
module VerilogMultiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] ,
         \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180;
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INV_X1 U2 ( .A(n110), .ZN(n25) );
  INV_X1 U3 ( .A(n107), .ZN(n23) );
  INV_X1 U4 ( .A(n131), .ZN(n21) );
  INV_X1 U5 ( .A(n111), .ZN(n14) );
  INV_X1 U6 ( .A(n88), .ZN(n12) );
  INV_X1 U7 ( .A(n80), .ZN(n10) );
  INV_X1 U8 ( .A(n72), .ZN(n8) );
  INV_X1 U9 ( .A(n64), .ZN(n6) );
  INV_X1 U10 ( .A(n56), .ZN(n4) );
  INV_X1 U11 ( .A(n145), .ZN(n29) );
  INV_X1 U12 ( .A(n48), .ZN(n2) );
  INV_X1 U13 ( .A(n106), .ZN(n24) );
  INV_X1 U14 ( .A(n144), .ZN(n27) );
  INV_X1 U15 ( .A(n142), .ZN(n26) );
  INV_X1 U16 ( .A(n149), .ZN(n31) );
  INV_X1 U17 ( .A(n127), .ZN(n20) );
  INV_X1 U18 ( .A(n122), .ZN(n18) );
  INV_X1 U19 ( .A(n102), .ZN(n17) );
  INV_X1 U20 ( .A(n97), .ZN(n15) );
  INV_X1 U21 ( .A(n90), .ZN(n13) );
  INV_X1 U22 ( .A(n82), .ZN(n11) );
  INV_X1 U23 ( .A(n74), .ZN(n9) );
  INV_X1 U24 ( .A(n66), .ZN(n7) );
  INV_X1 U25 ( .A(n58), .ZN(n5) );
  INV_X1 U26 ( .A(n50), .ZN(n3) );
  INV_X1 U27 ( .A(n42), .ZN(n1) );
  INV_X1 U28 ( .A(n158), .ZN(n34) );
  INV_X1 U29 ( .A(n165), .ZN(n36) );
  INV_X1 U30 ( .A(n130), .ZN(n19) );
  INV_X1 U31 ( .A(n148), .ZN(n28) );
  INV_X1 U32 ( .A(n170), .ZN(n33) );
  INV_X1 U33 ( .A(n160), .ZN(n32) );
  INV_X1 U34 ( .A(n117), .ZN(n16) );
  INV_X1 U35 ( .A(n172), .ZN(n35) );
  INV_X1 U36 ( .A(n147), .ZN(n30) );
  INV_X1 U37 ( .A(n128), .ZN(n22) );
  INV_X1 U38 ( .A(n175), .ZN(n37) );
  INV_X1 U39 ( .A(n176), .ZN(n38) );
  INV_X1 U40 ( .A(n180), .ZN(SUM[30]) );
  XOR2_X1 U41 ( .A(n40), .B(n41), .Z(SUM[61]) );
  XOR2_X1 U42 ( .A(B[61]), .B(A[61]), .Z(n41) );
  OAI21_X1 U43 ( .B1(n42), .B2(n43), .A(n44), .ZN(n40) );
  XOR2_X1 U44 ( .A(n45), .B(n43), .Z(SUM[60]) );
  AOI21_X1 U45 ( .B1(n2), .B2(n46), .A(n47), .ZN(n43) );
  NAND2_X1 U46 ( .A1(n1), .A2(n44), .ZN(n45) );
  NAND2_X1 U47 ( .A1(B[60]), .A2(A[60]), .ZN(n44) );
  NOR2_X1 U48 ( .A1(B[60]), .A2(A[60]), .ZN(n42) );
  XOR2_X1 U49 ( .A(n46), .B(n49), .Z(SUM[59]) );
  NOR2_X1 U50 ( .A1(n47), .A2(n48), .ZN(n49) );
  NOR2_X1 U51 ( .A1(B[59]), .A2(A[59]), .ZN(n48) );
  AND2_X1 U52 ( .A1(B[59]), .A2(A[59]), .ZN(n47) );
  OAI21_X1 U53 ( .B1(n50), .B2(n51), .A(n52), .ZN(n46) );
  XOR2_X1 U54 ( .A(n53), .B(n51), .Z(SUM[58]) );
  AOI21_X1 U55 ( .B1(n4), .B2(n54), .A(n55), .ZN(n51) );
  NAND2_X1 U56 ( .A1(n3), .A2(n52), .ZN(n53) );
  NAND2_X1 U57 ( .A1(B[58]), .A2(A[58]), .ZN(n52) );
  NOR2_X1 U58 ( .A1(B[58]), .A2(A[58]), .ZN(n50) );
  XOR2_X1 U59 ( .A(n54), .B(n57), .Z(SUM[57]) );
  NOR2_X1 U60 ( .A1(n55), .A2(n56), .ZN(n57) );
  NOR2_X1 U61 ( .A1(B[57]), .A2(A[57]), .ZN(n56) );
  AND2_X1 U62 ( .A1(B[57]), .A2(A[57]), .ZN(n55) );
  OAI21_X1 U63 ( .B1(n58), .B2(n59), .A(n60), .ZN(n54) );
  XOR2_X1 U64 ( .A(n61), .B(n59), .Z(SUM[56]) );
  AOI21_X1 U65 ( .B1(n6), .B2(n62), .A(n63), .ZN(n59) );
  NAND2_X1 U66 ( .A1(n5), .A2(n60), .ZN(n61) );
  NAND2_X1 U67 ( .A1(B[56]), .A2(A[56]), .ZN(n60) );
  NOR2_X1 U68 ( .A1(B[56]), .A2(A[56]), .ZN(n58) );
  XOR2_X1 U69 ( .A(n62), .B(n65), .Z(SUM[55]) );
  NOR2_X1 U70 ( .A1(n63), .A2(n64), .ZN(n65) );
  NOR2_X1 U71 ( .A1(B[55]), .A2(A[55]), .ZN(n64) );
  AND2_X1 U72 ( .A1(B[55]), .A2(A[55]), .ZN(n63) );
  OAI21_X1 U73 ( .B1(n66), .B2(n67), .A(n68), .ZN(n62) );
  XOR2_X1 U74 ( .A(n69), .B(n67), .Z(SUM[54]) );
  AOI21_X1 U75 ( .B1(n8), .B2(n70), .A(n71), .ZN(n67) );
  NAND2_X1 U76 ( .A1(n7), .A2(n68), .ZN(n69) );
  NAND2_X1 U77 ( .A1(B[54]), .A2(A[54]), .ZN(n68) );
  NOR2_X1 U78 ( .A1(B[54]), .A2(A[54]), .ZN(n66) );
  XOR2_X1 U79 ( .A(n70), .B(n73), .Z(SUM[53]) );
  NOR2_X1 U80 ( .A1(n71), .A2(n72), .ZN(n73) );
  NOR2_X1 U81 ( .A1(B[53]), .A2(A[53]), .ZN(n72) );
  AND2_X1 U82 ( .A1(B[53]), .A2(A[53]), .ZN(n71) );
  OAI21_X1 U83 ( .B1(n74), .B2(n75), .A(n76), .ZN(n70) );
  XOR2_X1 U84 ( .A(n77), .B(n75), .Z(SUM[52]) );
  AOI21_X1 U85 ( .B1(n10), .B2(n78), .A(n79), .ZN(n75) );
  NAND2_X1 U86 ( .A1(n9), .A2(n76), .ZN(n77) );
  NAND2_X1 U87 ( .A1(B[52]), .A2(A[52]), .ZN(n76) );
  NOR2_X1 U88 ( .A1(B[52]), .A2(A[52]), .ZN(n74) );
  XOR2_X1 U89 ( .A(n78), .B(n81), .Z(SUM[51]) );
  NOR2_X1 U90 ( .A1(n79), .A2(n80), .ZN(n81) );
  NOR2_X1 U91 ( .A1(B[51]), .A2(A[51]), .ZN(n80) );
  AND2_X1 U92 ( .A1(B[51]), .A2(A[51]), .ZN(n79) );
  OAI21_X1 U93 ( .B1(n82), .B2(n83), .A(n84), .ZN(n78) );
  XOR2_X1 U94 ( .A(n85), .B(n83), .Z(SUM[50]) );
  AOI21_X1 U95 ( .B1(n12), .B2(n86), .A(n87), .ZN(n83) );
  NAND2_X1 U96 ( .A1(n11), .A2(n84), .ZN(n85) );
  NAND2_X1 U97 ( .A1(B[50]), .A2(A[50]), .ZN(n84) );
  NOR2_X1 U98 ( .A1(B[50]), .A2(A[50]), .ZN(n82) );
  XOR2_X1 U99 ( .A(n86), .B(n89), .Z(SUM[49]) );
  NOR2_X1 U100 ( .A1(n87), .A2(n88), .ZN(n89) );
  NOR2_X1 U101 ( .A1(B[49]), .A2(A[49]), .ZN(n88) );
  AND2_X1 U102 ( .A1(B[49]), .A2(A[49]), .ZN(n87) );
  OAI21_X1 U103 ( .B1(n90), .B2(n91), .A(n92), .ZN(n86) );
  XOR2_X1 U104 ( .A(n93), .B(n91), .Z(SUM[48]) );
  AOI21_X1 U105 ( .B1(n14), .B2(n94), .A(n95), .ZN(n91) );
  OAI21_X1 U106 ( .B1(n96), .B2(n97), .A(n98), .ZN(n94) );
  AOI21_X1 U107 ( .B1(n16), .B2(n99), .A(n100), .ZN(n96) );
  OAI21_X1 U108 ( .B1(n101), .B2(n102), .A(n103), .ZN(n99) );
  AOI21_X1 U109 ( .B1(n24), .B2(n104), .A(n105), .ZN(n101) );
  AOI221_X1 U110 ( .B1(n107), .B2(n108), .C1(n109), .C2(n107), .A(n110), .ZN(
        n106) );
  NAND2_X1 U111 ( .A1(n13), .A2(n92), .ZN(n93) );
  NAND2_X1 U112 ( .A1(B[48]), .A2(A[48]), .ZN(n92) );
  NOR2_X1 U113 ( .A1(B[48]), .A2(A[48]), .ZN(n90) );
  XOR2_X1 U114 ( .A(n112), .B(n113), .Z(SUM[47]) );
  NOR2_X1 U115 ( .A1(n95), .A2(n111), .ZN(n113) );
  NOR2_X1 U116 ( .A1(B[47]), .A2(A[47]), .ZN(n111) );
  AND2_X1 U117 ( .A1(B[47]), .A2(A[47]), .ZN(n95) );
  OAI21_X1 U118 ( .B1(n97), .B2(n114), .A(n98), .ZN(n112) );
  XOR2_X1 U119 ( .A(n115), .B(n114), .Z(SUM[46]) );
  AOI21_X1 U120 ( .B1(n16), .B2(n116), .A(n100), .ZN(n114) );
  NAND2_X1 U121 ( .A1(n15), .A2(n98), .ZN(n115) );
  NAND2_X1 U122 ( .A1(B[46]), .A2(A[46]), .ZN(n98) );
  NOR2_X1 U123 ( .A1(B[46]), .A2(A[46]), .ZN(n97) );
  XOR2_X1 U124 ( .A(n116), .B(n118), .Z(SUM[45]) );
  NOR2_X1 U125 ( .A1(n100), .A2(n117), .ZN(n118) );
  NOR2_X1 U126 ( .A1(B[45]), .A2(A[45]), .ZN(n117) );
  AND2_X1 U127 ( .A1(B[45]), .A2(A[45]), .ZN(n100) );
  OAI21_X1 U128 ( .B1(n102), .B2(n119), .A(n103), .ZN(n116) );
  XOR2_X1 U129 ( .A(n120), .B(n119), .Z(SUM[44]) );
  AOI21_X1 U130 ( .B1(n121), .B2(n104), .A(n105), .ZN(n119) );
  OAI21_X1 U131 ( .B1(n122), .B2(n123), .A(n124), .ZN(n105) );
  AOI21_X1 U132 ( .B1(n125), .B2(n19), .A(n126), .ZN(n123) );
  OAI21_X1 U133 ( .B1(n127), .B2(n128), .A(n129), .ZN(n125) );
  NOR4_X1 U134 ( .A1(n122), .A2(n130), .A3(n127), .A4(n131), .ZN(n104) );
  NAND2_X1 U135 ( .A1(n17), .A2(n103), .ZN(n120) );
  NAND2_X1 U136 ( .A1(B[44]), .A2(A[44]), .ZN(n103) );
  NOR2_X1 U137 ( .A1(B[44]), .A2(A[44]), .ZN(n102) );
  XOR2_X1 U138 ( .A(n132), .B(n133), .Z(SUM[43]) );
  AOI21_X1 U139 ( .B1(n134), .B2(n19), .A(n126), .ZN(n133) );
  NAND2_X1 U140 ( .A1(n18), .A2(n124), .ZN(n132) );
  NAND2_X1 U141 ( .A1(B[43]), .A2(A[43]), .ZN(n124) );
  NOR2_X1 U142 ( .A1(B[43]), .A2(A[43]), .ZN(n122) );
  XOR2_X1 U143 ( .A(n134), .B(n135), .Z(SUM[42]) );
  NOR2_X1 U144 ( .A1(n126), .A2(n130), .ZN(n135) );
  NOR2_X1 U145 ( .A1(B[42]), .A2(A[42]), .ZN(n130) );
  AND2_X1 U146 ( .A1(B[42]), .A2(A[42]), .ZN(n126) );
  OAI21_X1 U147 ( .B1(n127), .B2(n136), .A(n129), .ZN(n134) );
  XOR2_X1 U148 ( .A(n137), .B(n136), .Z(SUM[41]) );
  AOI21_X1 U149 ( .B1(n21), .B2(n121), .A(n22), .ZN(n136) );
  NAND2_X1 U150 ( .A1(n20), .A2(n129), .ZN(n137) );
  NAND2_X1 U151 ( .A1(B[41]), .A2(A[41]), .ZN(n129) );
  NOR2_X1 U152 ( .A1(B[41]), .A2(A[41]), .ZN(n127) );
  XOR2_X1 U153 ( .A(n121), .B(n138), .Z(SUM[40]) );
  NOR2_X1 U154 ( .A1(n22), .A2(n131), .ZN(n138) );
  NOR2_X1 U155 ( .A1(B[40]), .A2(A[40]), .ZN(n131) );
  NAND2_X1 U156 ( .A1(B[40]), .A2(A[40]), .ZN(n128) );
  OAI21_X1 U157 ( .B1(n139), .B2(n23), .A(n25), .ZN(n121) );
  OAI21_X1 U158 ( .B1(n140), .B2(n141), .A(n142), .ZN(n110) );
  AOI21_X1 U159 ( .B1(n143), .B2(n28), .A(n27), .ZN(n141) );
  OAI21_X1 U160 ( .B1(n145), .B2(n146), .A(n147), .ZN(n143) );
  NOR4_X1 U161 ( .A1(n140), .A2(n148), .A3(n145), .A4(n149), .ZN(n107) );
  XOR2_X1 U162 ( .A(n150), .B(n151), .Z(SUM[39]) );
  NOR2_X1 U163 ( .A1(n26), .A2(n140), .ZN(n151) );
  NOR2_X1 U164 ( .A1(B[39]), .A2(A[39]), .ZN(n140) );
  NAND2_X1 U165 ( .A1(B[39]), .A2(A[39]), .ZN(n142) );
  OAI21_X1 U166 ( .B1(n148), .B2(n152), .A(n144), .ZN(n150) );
  XOR2_X1 U167 ( .A(n153), .B(n152), .Z(SUM[38]) );
  AOI21_X1 U168 ( .B1(n29), .B2(n154), .A(n30), .ZN(n152) );
  NAND2_X1 U169 ( .A1(n28), .A2(n144), .ZN(n153) );
  NAND2_X1 U170 ( .A1(B[38]), .A2(A[38]), .ZN(n144) );
  NOR2_X1 U171 ( .A1(B[38]), .A2(A[38]), .ZN(n148) );
  XOR2_X1 U172 ( .A(n154), .B(n155), .Z(SUM[37]) );
  NOR2_X1 U173 ( .A1(n30), .A2(n145), .ZN(n155) );
  NOR2_X1 U174 ( .A1(B[37]), .A2(A[37]), .ZN(n145) );
  NAND2_X1 U175 ( .A1(B[37]), .A2(A[37]), .ZN(n147) );
  OAI21_X1 U176 ( .B1(n149), .B2(n139), .A(n146), .ZN(n154) );
  XOR2_X1 U177 ( .A(n156), .B(n139), .Z(SUM[36]) );
  NOR2_X1 U178 ( .A1(n108), .A2(n109), .ZN(n139) );
  NOR4_X1 U179 ( .A1(n37), .A2(n157), .A3(n158), .A4(n159), .ZN(n109) );
  NAND2_X1 U180 ( .A1(n33), .A2(n32), .ZN(n159) );
  OAI21_X1 U181 ( .B1(n160), .B2(n161), .A(n162), .ZN(n108) );
  AOI21_X1 U182 ( .B1(n163), .B2(n33), .A(n164), .ZN(n161) );
  OAI21_X1 U183 ( .B1(n158), .B2(n165), .A(n166), .ZN(n163) );
  NAND2_X1 U184 ( .A1(n31), .A2(n146), .ZN(n156) );
  NAND2_X1 U185 ( .A1(B[36]), .A2(A[36]), .ZN(n146) );
  NOR2_X1 U186 ( .A1(B[36]), .A2(A[36]), .ZN(n149) );
  XOR2_X1 U187 ( .A(n167), .B(n168), .Z(SUM[35]) );
  AOI21_X1 U188 ( .B1(n169), .B2(n33), .A(n164), .ZN(n168) );
  NAND2_X1 U189 ( .A1(n32), .A2(n162), .ZN(n167) );
  NAND2_X1 U190 ( .A1(B[35]), .A2(A[35]), .ZN(n162) );
  NOR2_X1 U191 ( .A1(B[35]), .A2(A[35]), .ZN(n160) );
  XOR2_X1 U192 ( .A(n169), .B(n171), .Z(SUM[34]) );
  NOR2_X1 U193 ( .A1(n164), .A2(n170), .ZN(n171) );
  NOR2_X1 U194 ( .A1(B[34]), .A2(A[34]), .ZN(n170) );
  AND2_X1 U195 ( .A1(B[34]), .A2(A[34]), .ZN(n164) );
  OAI21_X1 U196 ( .B1(n158), .B2(n35), .A(n166), .ZN(n169) );
  XNOR2_X1 U197 ( .A(n173), .B(n172), .ZN(SUM[33]) );
  OAI21_X1 U198 ( .B1(n157), .B2(n37), .A(n165), .ZN(n172) );
  NAND2_X1 U199 ( .A1(n34), .A2(n166), .ZN(n173) );
  NAND2_X1 U200 ( .A1(B[33]), .A2(A[33]), .ZN(n166) );
  NOR2_X1 U201 ( .A1(B[33]), .A2(A[33]), .ZN(n158) );
  XNOR2_X1 U202 ( .A(n37), .B(n174), .ZN(SUM[32]) );
  NOR2_X1 U203 ( .A1(n36), .A2(n157), .ZN(n174) );
  NOR2_X1 U204 ( .A1(B[32]), .A2(A[32]), .ZN(n157) );
  NAND2_X1 U205 ( .A1(B[32]), .A2(A[32]), .ZN(n165) );
  OAI21_X1 U206 ( .B1(n176), .B2(n177), .A(n178), .ZN(n175) );
  XOR2_X1 U207 ( .A(n177), .B(n179), .Z(SUM[31]) );
  NAND2_X1 U208 ( .A1(n38), .A2(n178), .ZN(n179) );
  NAND2_X1 U209 ( .A1(B[31]), .A2(A[31]), .ZN(n178) );
  NOR2_X1 U210 ( .A1(B[31]), .A2(A[31]), .ZN(n176) );
  OAI21_X1 U211 ( .B1(B[30]), .B2(A[30]), .A(n177), .ZN(n180) );
  NAND2_X1 U212 ( .A1(B[30]), .A2(A[30]), .ZN(n177) );
endmodule


module VerilogMultiplier_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \ab[31][31] , \ab[31][30] , \ab[31][29] , \ab[31][28] , \ab[31][27] ,
         \ab[31][26] , \ab[31][25] , \ab[31][24] , \ab[31][23] , \ab[31][22] ,
         \ab[31][21] , \ab[31][20] , \ab[31][19] , \ab[31][18] , \ab[31][17] ,
         \ab[31][16] , \ab[31][15] , \ab[31][14] , \ab[31][13] , \ab[31][12] ,
         \ab[31][11] , \ab[31][10] , \ab[31][9] , \ab[31][8] , \ab[31][7] ,
         \ab[31][6] , \ab[31][5] , \ab[31][4] , \ab[31][3] , \ab[31][2] ,
         \ab[31][1] , \ab[31][0] , \ab[30][31] , \ab[30][30] , \ab[30][29] ,
         \ab[30][28] , \ab[30][27] , \ab[30][26] , \ab[30][25] , \ab[30][24] ,
         \ab[30][23] , \ab[30][22] , \ab[30][21] , \ab[30][20] , \ab[30][19] ,
         \ab[30][18] , \ab[30][17] , \ab[30][16] , \ab[30][15] , \ab[30][14] ,
         \ab[30][13] , \ab[30][12] , \ab[30][11] , \ab[30][10] , \ab[30][9] ,
         \ab[30][8] , \ab[30][7] , \ab[30][6] , \ab[30][5] , \ab[30][4] ,
         \ab[30][3] , \ab[30][2] , \ab[30][1] , \ab[30][0] , \ab[29][31] ,
         \ab[29][30] , \ab[29][29] , \ab[29][28] , \ab[29][27] , \ab[29][26] ,
         \ab[29][25] , \ab[29][24] , \ab[29][23] , \ab[29][22] , \ab[29][21] ,
         \ab[29][20] , \ab[29][19] , \ab[29][18] , \ab[29][17] , \ab[29][16] ,
         \ab[29][15] , \ab[29][14] , \ab[29][13] , \ab[29][12] , \ab[29][11] ,
         \ab[29][10] , \ab[29][9] , \ab[29][8] , \ab[29][7] , \ab[29][6] ,
         \ab[29][5] , \ab[29][4] , \ab[29][3] , \ab[29][2] , \ab[29][1] ,
         \ab[29][0] , \ab[28][31] , \ab[28][30] , \ab[28][29] , \ab[28][28] ,
         \ab[28][27] , \ab[28][26] , \ab[28][25] , \ab[28][24] , \ab[28][23] ,
         \ab[28][22] , \ab[28][21] , \ab[28][20] , \ab[28][19] , \ab[28][18] ,
         \ab[28][17] , \ab[28][16] , \ab[28][15] , \ab[28][14] , \ab[28][13] ,
         \ab[28][12] , \ab[28][11] , \ab[28][10] , \ab[28][9] , \ab[28][8] ,
         \ab[28][7] , \ab[28][6] , \ab[28][5] , \ab[28][4] , \ab[28][3] ,
         \ab[28][2] , \ab[28][1] , \ab[28][0] , \ab[27][31] , \ab[27][30] ,
         \ab[27][29] , \ab[27][28] , \ab[27][27] , \ab[27][26] , \ab[27][25] ,
         \ab[27][24] , \ab[27][23] , \ab[27][22] , \ab[27][21] , \ab[27][20] ,
         \ab[27][19] , \ab[27][18] , \ab[27][17] , \ab[27][16] , \ab[27][15] ,
         \ab[27][14] , \ab[27][13] , \ab[27][12] , \ab[27][11] , \ab[27][10] ,
         \ab[27][9] , \ab[27][8] , \ab[27][7] , \ab[27][6] , \ab[27][5] ,
         \ab[27][4] , \ab[27][3] , \ab[27][2] , \ab[27][1] , \ab[27][0] ,
         \ab[26][31] , \ab[26][30] , \ab[26][29] , \ab[26][28] , \ab[26][27] ,
         \ab[26][26] , \ab[26][25] , \ab[26][24] , \ab[26][23] , \ab[26][22] ,
         \ab[26][21] , \ab[26][20] , \ab[26][19] , \ab[26][18] , \ab[26][17] ,
         \ab[26][16] , \ab[26][15] , \ab[26][14] , \ab[26][13] , \ab[26][12] ,
         \ab[26][11] , \ab[26][10] , \ab[26][9] , \ab[26][8] , \ab[26][7] ,
         \ab[26][6] , \ab[26][5] , \ab[26][4] , \ab[26][3] , \ab[26][2] ,
         \ab[26][1] , \ab[26][0] , \ab[25][31] , \ab[25][30] , \ab[25][29] ,
         \ab[25][28] , \ab[25][27] , \ab[25][26] , \ab[25][25] , \ab[25][24] ,
         \ab[25][23] , \ab[25][22] , \ab[25][21] , \ab[25][20] , \ab[25][19] ,
         \ab[25][18] , \ab[25][17] , \ab[25][16] , \ab[25][15] , \ab[25][14] ,
         \ab[25][13] , \ab[25][12] , \ab[25][11] , \ab[25][10] , \ab[25][9] ,
         \ab[25][8] , \ab[25][7] , \ab[25][6] , \ab[25][5] , \ab[25][4] ,
         \ab[25][3] , \ab[25][2] , \ab[25][1] , \ab[25][0] , \ab[24][31] ,
         \ab[24][30] , \ab[24][29] , \ab[24][28] , \ab[24][27] , \ab[24][26] ,
         \ab[24][25] , \ab[24][24] , \ab[24][23] , \ab[24][22] , \ab[24][21] ,
         \ab[24][20] , \ab[24][19] , \ab[24][18] , \ab[24][17] , \ab[24][16] ,
         \ab[24][15] , \ab[24][14] , \ab[24][13] , \ab[24][12] , \ab[24][11] ,
         \ab[24][10] , \ab[24][9] , \ab[24][8] , \ab[24][7] , \ab[24][6] ,
         \ab[24][5] , \ab[24][4] , \ab[24][3] , \ab[24][2] , \ab[24][1] ,
         \ab[24][0] , \ab[23][31] , \ab[23][30] , \ab[23][29] , \ab[23][28] ,
         \ab[23][27] , \ab[23][26] , \ab[23][25] , \ab[23][24] , \ab[23][23] ,
         \ab[23][22] , \ab[23][21] , \ab[23][20] , \ab[23][19] , \ab[23][18] ,
         \ab[23][17] , \ab[23][16] , \ab[23][15] , \ab[23][14] , \ab[23][13] ,
         \ab[23][12] , \ab[23][11] , \ab[23][10] , \ab[23][9] , \ab[23][8] ,
         \ab[23][7] , \ab[23][6] , \ab[23][5] , \ab[23][4] , \ab[23][3] ,
         \ab[23][2] , \ab[23][1] , \ab[23][0] , \ab[22][31] , \ab[22][30] ,
         \ab[22][29] , \ab[22][28] , \ab[22][27] , \ab[22][26] , \ab[22][25] ,
         \ab[22][24] , \ab[22][23] , \ab[22][22] , \ab[22][21] , \ab[22][20] ,
         \ab[22][19] , \ab[22][18] , \ab[22][17] , \ab[22][16] , \ab[22][15] ,
         \ab[22][14] , \ab[22][13] , \ab[22][12] , \ab[22][11] , \ab[22][10] ,
         \ab[22][9] , \ab[22][8] , \ab[22][7] , \ab[22][6] , \ab[22][5] ,
         \ab[22][4] , \ab[22][3] , \ab[22][2] , \ab[22][1] , \ab[22][0] ,
         \ab[21][31] , \ab[21][30] , \ab[21][29] , \ab[21][28] , \ab[21][27] ,
         \ab[21][26] , \ab[21][25] , \ab[21][24] , \ab[21][23] , \ab[21][22] ,
         \ab[21][21] , \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] ,
         \ab[21][16] , \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] ,
         \ab[21][11] , \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] ,
         \ab[21][6] , \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] ,
         \ab[21][1] , \ab[21][0] , \ab[20][31] , \ab[20][30] , \ab[20][29] ,
         \ab[20][28] , \ab[20][27] , \ab[20][26] , \ab[20][25] , \ab[20][24] ,
         \ab[20][23] , \ab[20][22] , \ab[20][21] , \ab[20][20] , \ab[20][19] ,
         \ab[20][18] , \ab[20][17] , \ab[20][16] , \ab[20][15] , \ab[20][14] ,
         \ab[20][13] , \ab[20][12] , \ab[20][11] , \ab[20][10] , \ab[20][9] ,
         \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][5] , \ab[20][4] ,
         \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] , \ab[19][31] ,
         \ab[19][30] , \ab[19][29] , \ab[19][28] , \ab[19][27] , \ab[19][26] ,
         \ab[19][25] , \ab[19][24] , \ab[19][23] , \ab[19][22] , \ab[19][21] ,
         \ab[19][20] , \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] ,
         \ab[19][15] , \ab[19][14] , \ab[19][13] , \ab[19][12] , \ab[19][11] ,
         \ab[19][10] , \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] ,
         \ab[19][5] , \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] ,
         \ab[19][0] , \ab[18][31] , \ab[18][30] , \ab[18][29] , \ab[18][28] ,
         \ab[18][27] , \ab[18][26] , \ab[18][25] , \ab[18][24] , \ab[18][23] ,
         \ab[18][22] , \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] ,
         \ab[18][17] , \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] ,
         \ab[18][12] , \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] ,
         \ab[18][7] , \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] ,
         \ab[18][2] , \ab[18][1] , \ab[18][0] , \ab[17][31] , \ab[17][30] ,
         \ab[17][29] , \ab[17][28] , \ab[17][27] , \ab[17][26] , \ab[17][25] ,
         \ab[17][24] , \ab[17][23] , \ab[17][22] , \ab[17][21] , \ab[17][20] ,
         \ab[17][19] , \ab[17][18] , \ab[17][17] , \ab[17][16] , \ab[17][15] ,
         \ab[17][14] , \ab[17][13] , \ab[17][12] , \ab[17][11] , \ab[17][10] ,
         \ab[17][9] , \ab[17][8] , \ab[17][7] , \ab[17][6] , \ab[17][5] ,
         \ab[17][4] , \ab[17][3] , \ab[17][2] , \ab[17][1] , \ab[17][0] ,
         \ab[16][31] , \ab[16][30] , \ab[16][29] , \ab[16][28] , \ab[16][27] ,
         \ab[16][26] , \ab[16][25] , \ab[16][24] , \ab[16][23] , \ab[16][22] ,
         \ab[16][21] , \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] ,
         \ab[16][16] , \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] ,
         \ab[16][11] , \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] ,
         \ab[16][6] , \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] ,
         \ab[16][1] , \ab[16][0] , \ab[15][31] , \ab[15][30] , \ab[15][29] ,
         \ab[15][28] , \ab[15][27] , \ab[15][26] , \ab[15][25] , \ab[15][24] ,
         \ab[15][23] , \ab[15][22] , \ab[15][21] , \ab[15][20] , \ab[15][19] ,
         \ab[15][18] , \ab[15][17] , \ab[15][16] , \ab[15][15] , \ab[15][14] ,
         \ab[15][13] , \ab[15][12] , \ab[15][11] , \ab[15][10] , \ab[15][9] ,
         \ab[15][8] , \ab[15][7] , \ab[15][6] , \ab[15][5] , \ab[15][4] ,
         \ab[15][3] , \ab[15][2] , \ab[15][1] , \ab[15][0] , \ab[14][31] ,
         \ab[14][30] , \ab[14][29] , \ab[14][28] , \ab[14][27] , \ab[14][26] ,
         \ab[14][25] , \ab[14][24] , \ab[14][23] , \ab[14][22] , \ab[14][21] ,
         \ab[14][20] , \ab[14][19] , \ab[14][18] , \ab[14][17] , \ab[14][16] ,
         \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] ,
         \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] ,
         \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] ,
         \ab[14][0] , \ab[13][31] , \ab[13][30] , \ab[13][29] , \ab[13][28] ,
         \ab[13][27] , \ab[13][26] , \ab[13][25] , \ab[13][24] , \ab[13][23] ,
         \ab[13][22] , \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] ,
         \ab[13][17] , \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][31] , \ab[12][30] ,
         \ab[12][29] , \ab[12][28] , \ab[12][27] , \ab[12][26] , \ab[12][25] ,
         \ab[12][24] , \ab[12][23] , \ab[12][22] , \ab[12][21] , \ab[12][20] ,
         \ab[12][19] , \ab[12][18] , \ab[12][17] , \ab[12][16] , \ab[12][15] ,
         \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] ,
         \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] ,
         \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][31] , \ab[11][30] , \ab[11][29] , \ab[11][28] , \ab[11][27] ,
         \ab[11][26] , \ab[11][25] , \ab[11][24] , \ab[11][23] , \ab[11][22] ,
         \ab[11][21] , \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] ,
         \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] ,
         \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] ,
         \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] ,
         \ab[11][1] , \ab[11][0] , \ab[10][31] , \ab[10][30] , \ab[10][29] ,
         \ab[10][28] , \ab[10][27] , \ab[10][26] , \ab[10][25] , \ab[10][24] ,
         \ab[10][23] , \ab[10][22] , \ab[10][21] , \ab[10][20] , \ab[10][19] ,
         \ab[10][18] , \ab[10][17] , \ab[10][16] , \ab[10][15] , \ab[10][14] ,
         \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] ,
         \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] ,
         \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][31] ,
         \ab[9][30] , \ab[9][29] , \ab[9][28] , \ab[9][27] , \ab[9][26] ,
         \ab[9][25] , \ab[9][24] , \ab[9][23] , \ab[9][22] , \ab[9][21] ,
         \ab[9][20] , \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] ,
         \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] ,
         \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] ,
         \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] ,
         \ab[9][0] , \ab[8][31] , \ab[8][30] , \ab[8][29] , \ab[8][28] ,
         \ab[8][27] , \ab[8][26] , \ab[8][25] , \ab[8][24] , \ab[8][23] ,
         \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] ,
         \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][31] , \ab[7][30] ,
         \ab[7][29] , \ab[7][28] , \ab[7][27] , \ab[7][26] , \ab[7][25] ,
         \ab[7][24] , \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] ,
         \ab[7][19] , \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][31] , \ab[6][30] , \ab[6][29] , \ab[6][28] , \ab[6][27] ,
         \ab[6][26] , \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] ,
         \ab[6][21] , \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] ,
         \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] ,
         \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] ,
         \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] ,
         \ab[6][1] , \ab[6][0] , \ab[5][31] , \ab[5][30] , \ab[5][29] ,
         \ab[5][28] , \ab[5][27] , \ab[5][26] , \ab[5][25] , \ab[5][24] ,
         \ab[5][23] , \ab[5][22] , \ab[5][21] , \ab[5][20] , \ab[5][19] ,
         \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][15] , \ab[5][14] ,
         \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] ,
         \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] ,
         \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][31] ,
         \ab[4][30] , \ab[4][29] , \ab[4][28] , \ab[4][27] , \ab[4][26] ,
         \ab[4][25] , \ab[4][24] , \ab[4][23] , \ab[4][22] , \ab[4][21] ,
         \ab[4][20] , \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] ,
         \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] ,
         \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] ,
         \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] ,
         \ab[4][0] , \ab[3][31] , \ab[3][30] , \ab[3][29] , \ab[3][28] ,
         \ab[3][27] , \ab[3][26] , \ab[3][25] , \ab[3][24] , \ab[3][23] ,
         \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] ,
         \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][31] , \ab[2][30] ,
         \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] , \ab[2][25] ,
         \ab[2][24] , \ab[2][23] , \ab[2][22] , \ab[2][21] , \ab[2][20] ,
         \ab[2][19] , \ab[2][18] , \ab[2][17] , \ab[2][16] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][31] , \ab[1][30] , \ab[1][29] , \ab[1][28] , \ab[1][27] ,
         \ab[1][26] , \ab[1][25] , \ab[1][24] , \ab[1][23] , \ab[1][22] ,
         \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] ,
         \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] ,
         \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] ,
         \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] ,
         \ab[1][1] , \ab[1][0] , \ab[0][31] , \ab[0][30] , \ab[0][29] ,
         \ab[0][28] , \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] ,
         \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] ,
         \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[15][30] ,
         \CARRYB[15][29] , \CARRYB[15][28] , \CARRYB[15][27] ,
         \CARRYB[15][26] , \CARRYB[15][25] , \CARRYB[15][24] ,
         \CARRYB[15][23] , \CARRYB[15][22] , \CARRYB[15][21] ,
         \CARRYB[15][20] , \CARRYB[15][19] , \CARRYB[15][18] ,
         \CARRYB[15][17] , \CARRYB[15][16] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][30] , \CARRYB[13][29] , \CARRYB[13][28] ,
         \CARRYB[13][27] , \CARRYB[13][26] , \CARRYB[13][25] ,
         \CARRYB[13][24] , \CARRYB[13][23] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][30] , \CARRYB[11][29] , \CARRYB[11][28] ,
         \CARRYB[11][27] , \CARRYB[11][26] , \CARRYB[11][25] ,
         \CARRYB[11][24] , \CARRYB[11][23] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][30] , \CARRYB[10][29] , \CARRYB[10][28] ,
         \CARRYB[10][27] , \CARRYB[10][26] , \CARRYB[10][25] ,
         \CARRYB[10][24] , \CARRYB[10][23] , \CARRYB[10][22] ,
         \CARRYB[10][21] , \CARRYB[10][20] , \CARRYB[10][19] ,
         \CARRYB[10][18] , \CARRYB[10][17] , \CARRYB[10][16] ,
         \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][30] , \CARRYB[9][29] , \CARRYB[9][28] ,
         \CARRYB[9][27] , \CARRYB[9][26] , \CARRYB[9][25] , \CARRYB[9][24] ,
         \CARRYB[9][23] , \CARRYB[9][22] , \CARRYB[9][21] , \CARRYB[9][20] ,
         \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] , \CARRYB[9][16] ,
         \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] ,
         \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] ,
         \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] ,
         \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] ,
         \CARRYB[8][30] , \CARRYB[8][29] , \CARRYB[8][28] , \CARRYB[8][27] ,
         \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] , \CARRYB[8][23] ,
         \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] , \CARRYB[8][19] ,
         \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] , \CARRYB[8][15] ,
         \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] ,
         \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] ,
         \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] ,
         \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][30] ,
         \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] , \CARRYB[7][26] ,
         \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] ,
         \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] ,
         \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][30] , \CARRYB[6][29] ,
         \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][30] , \CARRYB[5][29] , \CARRYB[5][28] ,
         \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] , \CARRYB[5][24] ,
         \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] , \CARRYB[5][20] ,
         \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] , \CARRYB[5][16] ,
         \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] ,
         \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] ,
         \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] ,
         \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] ,
         \CARRYB[4][30] , \CARRYB[4][29] , \CARRYB[4][28] , \CARRYB[4][27] ,
         \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] , \CARRYB[4][23] ,
         \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] , \CARRYB[4][19] ,
         \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][15] ,
         \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] ,
         \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] ,
         \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] ,
         \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][30] ,
         \CARRYB[3][29] , \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] ,
         \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][30] , \CARRYB[2][29] ,
         \CARRYB[2][28] , \CARRYB[2][27] , \CARRYB[2][26] , \CARRYB[2][25] ,
         \CARRYB[2][24] , \CARRYB[2][23] , \CARRYB[2][22] , \CARRYB[2][21] ,
         \CARRYB[2][20] , \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] ,
         \CARRYB[2][16] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[15][30] , \SUMB[15][29] , \SUMB[15][28] ,
         \SUMB[15][27] , \SUMB[15][26] , \SUMB[15][25] , \SUMB[15][24] ,
         \SUMB[15][23] , \SUMB[15][22] , \SUMB[15][21] , \SUMB[15][20] ,
         \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] , \SUMB[15][16] ,
         \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] ,
         \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] ,
         \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] ,
         \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][30] ,
         \SUMB[14][29] , \SUMB[14][28] , \SUMB[14][27] , \SUMB[14][26] ,
         \SUMB[14][25] , \SUMB[14][24] , \SUMB[14][23] , \SUMB[14][22] ,
         \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] , \SUMB[14][18] ,
         \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][30] , \SUMB[13][29] , \SUMB[13][28] ,
         \SUMB[13][27] , \SUMB[13][26] , \SUMB[13][25] , \SUMB[13][24] ,
         \SUMB[13][23] , \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] ,
         \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] ,
         \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][30] ,
         \SUMB[12][29] , \SUMB[12][28] , \SUMB[12][27] , \SUMB[12][26] ,
         \SUMB[12][25] , \SUMB[12][24] , \SUMB[12][23] , \SUMB[12][22] ,
         \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] ,
         \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][30] , \SUMB[11][29] , \SUMB[11][28] ,
         \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] ,
         \SUMB[11][23] , \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] ,
         \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][30] ,
         \SUMB[10][29] , \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] ,
         \SUMB[10][25] , \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] ,
         \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] ,
         \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][30] , \SUMB[9][29] , \SUMB[9][28] ,
         \SUMB[9][27] , \SUMB[9][26] , \SUMB[9][25] , \SUMB[9][24] ,
         \SUMB[9][23] , \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] ,
         \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] ,
         \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][30] , \SUMB[8][29] ,
         \SUMB[8][28] , \SUMB[8][27] , \SUMB[8][26] , \SUMB[8][25] ,
         \SUMB[8][24] , \SUMB[8][23] , \SUMB[8][22] , \SUMB[8][21] ,
         \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] , \SUMB[8][17] ,
         \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][30] ,
         \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] , \SUMB[7][26] ,
         \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][30] ,
         \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] ,
         \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][30] ,
         \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] ,
         \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][30] ,
         \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] ,
         \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \CARRYB[31][31] , \CARRYB[31][30] , \CARRYB[31][29] ,
         \CARRYB[31][28] , \CARRYB[31][27] , \CARRYB[31][26] ,
         \CARRYB[31][25] , \CARRYB[31][24] , \CARRYB[31][23] ,
         \CARRYB[31][22] , \CARRYB[31][21] , \CARRYB[31][20] ,
         \CARRYB[31][19] , \CARRYB[31][18] , \CARRYB[31][17] ,
         \CARRYB[31][16] , \CARRYB[31][15] , \CARRYB[31][14] ,
         \CARRYB[31][13] , \CARRYB[31][12] , \CARRYB[31][11] ,
         \CARRYB[31][10] , \CARRYB[31][9] , \CARRYB[31][8] , \CARRYB[31][7] ,
         \CARRYB[31][6] , \CARRYB[31][5] , \CARRYB[31][4] , \CARRYB[31][3] ,
         \CARRYB[31][2] , \CARRYB[31][1] , \CARRYB[31][0] , \CARRYB[30][30] ,
         \CARRYB[30][29] , \CARRYB[30][28] , \CARRYB[30][27] ,
         \CARRYB[30][26] , \CARRYB[30][25] , \CARRYB[30][24] ,
         \CARRYB[30][23] , \CARRYB[30][22] , \CARRYB[30][21] ,
         \CARRYB[30][20] , \CARRYB[30][19] , \CARRYB[30][18] ,
         \CARRYB[30][17] , \CARRYB[30][16] , \CARRYB[30][15] ,
         \CARRYB[30][14] , \CARRYB[30][13] , \CARRYB[30][12] ,
         \CARRYB[30][11] , \CARRYB[30][10] , \CARRYB[30][9] , \CARRYB[30][8] ,
         \CARRYB[30][7] , \CARRYB[30][6] , \CARRYB[30][5] , \CARRYB[30][4] ,
         \CARRYB[30][3] , \CARRYB[30][2] , \CARRYB[30][1] , \CARRYB[30][0] ,
         \CARRYB[29][30] , \CARRYB[29][29] , \CARRYB[29][28] ,
         \CARRYB[29][27] , \CARRYB[29][26] , \CARRYB[29][25] ,
         \CARRYB[29][24] , \CARRYB[29][23] , \CARRYB[29][22] ,
         \CARRYB[29][21] , \CARRYB[29][20] , \CARRYB[29][19] ,
         \CARRYB[29][18] , \CARRYB[29][17] , \CARRYB[29][16] ,
         \CARRYB[29][15] , \CARRYB[29][14] , \CARRYB[29][13] ,
         \CARRYB[29][12] , \CARRYB[29][11] , \CARRYB[29][10] , \CARRYB[29][9] ,
         \CARRYB[29][8] , \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][5] ,
         \CARRYB[29][4] , \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][30] , \CARRYB[28][29] , \CARRYB[28][28] ,
         \CARRYB[28][27] , \CARRYB[28][26] , \CARRYB[28][25] ,
         \CARRYB[28][24] , \CARRYB[28][23] , \CARRYB[28][22] ,
         \CARRYB[28][21] , \CARRYB[28][20] , \CARRYB[28][19] ,
         \CARRYB[28][18] , \CARRYB[28][17] , \CARRYB[28][16] ,
         \CARRYB[28][15] , \CARRYB[28][14] , \CARRYB[28][13] ,
         \CARRYB[28][12] , \CARRYB[28][11] , \CARRYB[28][10] , \CARRYB[28][9] ,
         \CARRYB[28][8] , \CARRYB[28][7] , \CARRYB[28][6] , \CARRYB[28][5] ,
         \CARRYB[28][4] , \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][30] , \CARRYB[27][29] , \CARRYB[27][28] ,
         \CARRYB[27][27] , \CARRYB[27][26] , \CARRYB[27][25] ,
         \CARRYB[27][24] , \CARRYB[27][23] , \CARRYB[27][22] ,
         \CARRYB[27][21] , \CARRYB[27][20] , \CARRYB[27][19] ,
         \CARRYB[27][18] , \CARRYB[27][17] , \CARRYB[27][16] ,
         \CARRYB[27][15] , \CARRYB[27][14] , \CARRYB[27][13] ,
         \CARRYB[27][12] , \CARRYB[27][11] , \CARRYB[27][10] , \CARRYB[27][9] ,
         \CARRYB[27][8] , \CARRYB[27][7] , \CARRYB[27][6] , \CARRYB[27][5] ,
         \CARRYB[27][4] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][30] , \CARRYB[25][29] , \CARRYB[25][28] ,
         \CARRYB[25][27] , \CARRYB[25][26] , \CARRYB[25][25] ,
         \CARRYB[25][24] , \CARRYB[25][23] , \CARRYB[25][22] ,
         \CARRYB[25][21] , \CARRYB[25][20] , \CARRYB[25][19] ,
         \CARRYB[25][18] , \CARRYB[25][17] , \CARRYB[25][16] ,
         \CARRYB[25][15] , \CARRYB[25][14] , \CARRYB[25][13] ,
         \CARRYB[25][12] , \CARRYB[25][11] , \CARRYB[25][10] , \CARRYB[25][9] ,
         \CARRYB[25][8] , \CARRYB[25][7] , \CARRYB[25][6] , \CARRYB[25][5] ,
         \CARRYB[25][4] , \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] ,
         \CARRYB[25][0] , \CARRYB[24][30] , \CARRYB[24][29] , \CARRYB[24][28] ,
         \CARRYB[24][27] , \CARRYB[24][26] , \CARRYB[24][25] ,
         \CARRYB[24][24] , \CARRYB[24][23] , \CARRYB[24][22] ,
         \CARRYB[24][21] , \CARRYB[24][20] , \CARRYB[24][19] ,
         \CARRYB[24][18] , \CARRYB[24][17] , \CARRYB[24][16] ,
         \CARRYB[24][15] , \CARRYB[24][14] , \CARRYB[24][13] ,
         \CARRYB[24][12] , \CARRYB[24][11] , \CARRYB[24][10] , \CARRYB[24][9] ,
         \CARRYB[24][8] , \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] ,
         \CARRYB[24][4] , \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] ,
         \CARRYB[24][0] , \CARRYB[23][30] , \CARRYB[23][29] , \CARRYB[23][28] ,
         \CARRYB[23][27] , \CARRYB[23][26] , \CARRYB[23][25] ,
         \CARRYB[23][24] , \CARRYB[23][23] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][30] , \CARRYB[22][29] , \CARRYB[22][28] ,
         \CARRYB[22][27] , \CARRYB[22][26] , \CARRYB[22][25] ,
         \CARRYB[22][24] , \CARRYB[22][23] , \CARRYB[22][22] ,
         \CARRYB[22][21] , \CARRYB[22][20] , \CARRYB[22][19] ,
         \CARRYB[22][18] , \CARRYB[22][17] , \CARRYB[22][16] ,
         \CARRYB[22][15] , \CARRYB[22][14] , \CARRYB[22][13] ,
         \CARRYB[22][12] , \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] ,
         \CARRYB[22][8] , \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][30] , \CARRYB[21][29] , \CARRYB[21][28] ,
         \CARRYB[21][27] , \CARRYB[21][26] , \CARRYB[21][25] ,
         \CARRYB[21][24] , \CARRYB[21][23] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][30] , \CARRYB[19][29] , \CARRYB[19][28] ,
         \CARRYB[19][27] , \CARRYB[19][26] , \CARRYB[19][25] ,
         \CARRYB[19][24] , \CARRYB[19][23] , \CARRYB[19][22] ,
         \CARRYB[19][21] , \CARRYB[19][20] , \CARRYB[19][19] ,
         \CARRYB[19][18] , \CARRYB[19][17] , \CARRYB[19][16] ,
         \CARRYB[19][15] , \CARRYB[19][14] , \CARRYB[19][13] ,
         \CARRYB[19][12] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] ,
         \CARRYB[19][8] , \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] ,
         \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] ,
         \CARRYB[19][0] , \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][30] , \CARRYB[17][29] , \CARRYB[17][28] ,
         \CARRYB[17][27] , \CARRYB[17][26] , \CARRYB[17][25] ,
         \CARRYB[17][24] , \CARRYB[17][23] , \CARRYB[17][22] ,
         \CARRYB[17][21] , \CARRYB[17][20] , \CARRYB[17][19] ,
         \CARRYB[17][18] , \CARRYB[17][17] , \CARRYB[17][16] ,
         \CARRYB[17][15] , \CARRYB[17][14] , \CARRYB[17][13] ,
         \CARRYB[17][12] , \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] ,
         \CARRYB[17][8] , \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \SUMB[31][31] , \SUMB[31][30] , \SUMB[31][29] ,
         \SUMB[31][28] , \SUMB[31][27] , \SUMB[31][26] , \SUMB[31][25] ,
         \SUMB[31][24] , \SUMB[31][23] , \SUMB[31][22] , \SUMB[31][21] ,
         \SUMB[31][20] , \SUMB[31][19] , \SUMB[31][18] , \SUMB[31][17] ,
         \SUMB[31][16] , \SUMB[31][15] , \SUMB[31][14] , \SUMB[31][13] ,
         \SUMB[31][12] , \SUMB[31][11] , \SUMB[31][10] , \SUMB[31][9] ,
         \SUMB[31][8] , \SUMB[31][7] , \SUMB[31][6] , \SUMB[31][5] ,
         \SUMB[31][4] , \SUMB[31][3] , \SUMB[31][2] , \SUMB[31][1] ,
         \SUMB[31][0] , \SUMB[30][30] , \SUMB[30][29] , \SUMB[30][28] ,
         \SUMB[30][27] , \SUMB[30][26] , \SUMB[30][25] , \SUMB[30][24] ,
         \SUMB[30][23] , \SUMB[30][22] , \SUMB[30][21] , \SUMB[30][20] ,
         \SUMB[30][19] , \SUMB[30][18] , \SUMB[30][17] , \SUMB[30][16] ,
         \SUMB[30][15] , \SUMB[30][14] , \SUMB[30][13] , \SUMB[30][12] ,
         \SUMB[30][11] , \SUMB[30][10] , \SUMB[30][9] , \SUMB[30][8] ,
         \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][5] , \SUMB[30][4] ,
         \SUMB[30][3] , \SUMB[30][2] , \SUMB[30][1] , \SUMB[29][30] ,
         \SUMB[29][29] , \SUMB[29][28] , \SUMB[29][27] , \SUMB[29][26] ,
         \SUMB[29][25] , \SUMB[29][24] , \SUMB[29][23] , \SUMB[29][22] ,
         \SUMB[29][21] , \SUMB[29][20] , \SUMB[29][19] , \SUMB[29][18] ,
         \SUMB[29][17] , \SUMB[29][16] , \SUMB[29][15] , \SUMB[29][14] ,
         \SUMB[29][13] , \SUMB[29][12] , \SUMB[29][11] , \SUMB[29][10] ,
         \SUMB[29][9] , \SUMB[29][8] , \SUMB[29][7] , \SUMB[29][6] ,
         \SUMB[29][5] , \SUMB[29][4] , \SUMB[29][3] , \SUMB[29][2] ,
         \SUMB[29][1] , \SUMB[28][30] , \SUMB[28][29] , \SUMB[28][28] ,
         \SUMB[28][27] , \SUMB[28][26] , \SUMB[28][25] , \SUMB[28][24] ,
         \SUMB[28][23] , \SUMB[28][22] , \SUMB[28][21] , \SUMB[28][20] ,
         \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] , \SUMB[28][16] ,
         \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] , \SUMB[28][12] ,
         \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] , \SUMB[28][8] ,
         \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] , \SUMB[28][4] ,
         \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][30] ,
         \SUMB[27][29] , \SUMB[27][28] , \SUMB[27][27] , \SUMB[27][26] ,
         \SUMB[27][25] , \SUMB[27][24] , \SUMB[27][23] , \SUMB[27][22] ,
         \SUMB[27][21] , \SUMB[27][20] , \SUMB[27][19] , \SUMB[27][18] ,
         \SUMB[27][17] , \SUMB[27][16] , \SUMB[27][15] , \SUMB[27][14] ,
         \SUMB[27][13] , \SUMB[27][12] , \SUMB[27][11] , \SUMB[27][10] ,
         \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] , \SUMB[27][6] ,
         \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] , \SUMB[27][2] ,
         \SUMB[27][1] , \SUMB[26][30] , \SUMB[26][29] , \SUMB[26][28] ,
         \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] , \SUMB[26][24] ,
         \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] , \SUMB[26][20] ,
         \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] , \SUMB[26][16] ,
         \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] , \SUMB[26][12] ,
         \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] , \SUMB[26][8] ,
         \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][30] ,
         \SUMB[25][29] , \SUMB[25][28] , \SUMB[25][27] , \SUMB[25][26] ,
         \SUMB[25][25] , \SUMB[25][24] , \SUMB[25][23] , \SUMB[25][22] ,
         \SUMB[25][21] , \SUMB[25][20] , \SUMB[25][19] , \SUMB[25][18] ,
         \SUMB[25][17] , \SUMB[25][16] , \SUMB[25][15] , \SUMB[25][14] ,
         \SUMB[25][13] , \SUMB[25][12] , \SUMB[25][11] , \SUMB[25][10] ,
         \SUMB[25][9] , \SUMB[25][8] , \SUMB[25][7] , \SUMB[25][6] ,
         \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] ,
         \SUMB[25][1] , \SUMB[24][30] , \SUMB[24][29] , \SUMB[24][28] ,
         \SUMB[24][27] , \SUMB[24][26] , \SUMB[24][25] , \SUMB[24][24] ,
         \SUMB[24][23] , \SUMB[24][22] , \SUMB[24][21] , \SUMB[24][20] ,
         \SUMB[24][19] , \SUMB[24][18] , \SUMB[24][17] , \SUMB[24][16] ,
         \SUMB[24][15] , \SUMB[24][14] , \SUMB[24][13] , \SUMB[24][12] ,
         \SUMB[24][11] , \SUMB[24][10] , \SUMB[24][9] , \SUMB[24][8] ,
         \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][30] ,
         \SUMB[23][29] , \SUMB[23][28] , \SUMB[23][27] , \SUMB[23][26] ,
         \SUMB[23][25] , \SUMB[23][24] , \SUMB[23][23] , \SUMB[23][22] ,
         \SUMB[23][21] , \SUMB[23][20] , \SUMB[23][19] , \SUMB[23][18] ,
         \SUMB[23][17] , \SUMB[23][16] , \SUMB[23][15] , \SUMB[23][14] ,
         \SUMB[23][13] , \SUMB[23][12] , \SUMB[23][11] , \SUMB[23][10] ,
         \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] , \SUMB[23][6] ,
         \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] ,
         \SUMB[23][1] , \SUMB[22][30] , \SUMB[22][29] , \SUMB[22][28] ,
         \SUMB[22][27] , \SUMB[22][26] , \SUMB[22][25] , \SUMB[22][24] ,
         \SUMB[22][23] , \SUMB[22][22] , \SUMB[22][21] , \SUMB[22][20] ,
         \SUMB[22][19] , \SUMB[22][18] , \SUMB[22][17] , \SUMB[22][16] ,
         \SUMB[22][15] , \SUMB[22][14] , \SUMB[22][13] , \SUMB[22][12] ,
         \SUMB[22][11] , \SUMB[22][10] , \SUMB[22][9] , \SUMB[22][8] ,
         \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] ,
         \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][30] ,
         \SUMB[21][29] , \SUMB[21][28] , \SUMB[21][27] , \SUMB[21][26] ,
         \SUMB[21][25] , \SUMB[21][24] , \SUMB[21][23] , \SUMB[21][22] ,
         \SUMB[21][21] , \SUMB[21][20] , \SUMB[21][19] , \SUMB[21][18] ,
         \SUMB[21][17] , \SUMB[21][16] , \SUMB[21][15] , \SUMB[21][14] ,
         \SUMB[21][13] , \SUMB[21][12] , \SUMB[21][11] , \SUMB[21][10] ,
         \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] , \SUMB[21][6] ,
         \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] ,
         \SUMB[21][1] , \SUMB[20][30] , \SUMB[20][29] , \SUMB[20][28] ,
         \SUMB[20][27] , \SUMB[20][26] , \SUMB[20][25] , \SUMB[20][24] ,
         \SUMB[20][23] , \SUMB[20][22] , \SUMB[20][21] , \SUMB[20][20] ,
         \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] , \SUMB[20][16] ,
         \SUMB[20][15] , \SUMB[20][14] , \SUMB[20][13] , \SUMB[20][12] ,
         \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] ,
         \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][30] ,
         \SUMB[19][29] , \SUMB[19][28] , \SUMB[19][27] , \SUMB[19][26] ,
         \SUMB[19][25] , \SUMB[19][24] , \SUMB[19][23] , \SUMB[19][22] ,
         \SUMB[19][21] , \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] ,
         \SUMB[19][17] , \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] ,
         \SUMB[19][13] , \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] ,
         \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][30] , \SUMB[18][29] , \SUMB[18][28] ,
         \SUMB[18][27] , \SUMB[18][26] , \SUMB[18][25] , \SUMB[18][24] ,
         \SUMB[18][23] , \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] ,
         \SUMB[18][19] , \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] ,
         \SUMB[18][15] , \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] ,
         \SUMB[18][11] , \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] ,
         \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] ,
         \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][30] ,
         \SUMB[17][29] , \SUMB[17][28] , \SUMB[17][27] , \SUMB[17][26] ,
         \SUMB[17][25] , \SUMB[17][24] , \SUMB[17][23] , \SUMB[17][22] ,
         \SUMB[17][21] , \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] ,
         \SUMB[17][17] , \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] ,
         \SUMB[17][13] , \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] ,
         \SUMB[17][9] , \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] ,
         \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] ,
         \SUMB[17][1] , \SUMB[16][30] , \SUMB[16][29] , \SUMB[16][28] ,
         \SUMB[16][27] , \SUMB[16][26] , \SUMB[16][25] , \SUMB[16][24] ,
         \SUMB[16][23] , \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] ,
         \SUMB[16][19] , \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] ,
         \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] ,
         \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] ,
         \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , ZA, ZB, \A1[29] ,
         \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[30] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380;
  assign ZA = A[31];
  assign ZB = B[31];

  FA_X1 S14_31_0 ( .A(ZA), .B(ZB), .CI(\SUMB[31][0] ), .CO(\A2[30] ), .S(
        \A1[29] ) );
  FA_X1 S4_0 ( .A(\ab[31][0] ), .B(\CARRYB[30][0] ), .CI(\SUMB[30][1] ), .CO(
        \CARRYB[31][0] ), .S(\SUMB[31][0] ) );
  FA_X1 S4_1 ( .A(\ab[31][1] ), .B(\CARRYB[30][1] ), .CI(\SUMB[30][2] ), .CO(
        \CARRYB[31][1] ), .S(\SUMB[31][1] ) );
  FA_X1 S4_2 ( .A(\ab[31][2] ), .B(\CARRYB[30][2] ), .CI(\SUMB[30][3] ), .CO(
        \CARRYB[31][2] ), .S(\SUMB[31][2] ) );
  FA_X1 S4_3 ( .A(\ab[31][3] ), .B(\CARRYB[30][3] ), .CI(\SUMB[30][4] ), .CO(
        \CARRYB[31][3] ), .S(\SUMB[31][3] ) );
  FA_X1 S4_4 ( .A(\ab[31][4] ), .B(\CARRYB[30][4] ), .CI(\SUMB[30][5] ), .CO(
        \CARRYB[31][4] ), .S(\SUMB[31][4] ) );
  FA_X1 S4_5 ( .A(\ab[31][5] ), .B(\CARRYB[30][5] ), .CI(\SUMB[30][6] ), .CO(
        \CARRYB[31][5] ), .S(\SUMB[31][5] ) );
  FA_X1 S4_6 ( .A(\ab[31][6] ), .B(\CARRYB[30][6] ), .CI(\SUMB[30][7] ), .CO(
        \CARRYB[31][6] ), .S(\SUMB[31][6] ) );
  FA_X1 S4_7 ( .A(\ab[31][7] ), .B(\CARRYB[30][7] ), .CI(\SUMB[30][8] ), .CO(
        \CARRYB[31][7] ), .S(\SUMB[31][7] ) );
  FA_X1 S4_8 ( .A(\ab[31][8] ), .B(\CARRYB[30][8] ), .CI(\SUMB[30][9] ), .CO(
        \CARRYB[31][8] ), .S(\SUMB[31][8] ) );
  FA_X1 S4_9 ( .A(\ab[31][9] ), .B(\CARRYB[30][9] ), .CI(\SUMB[30][10] ), .CO(
        \CARRYB[31][9] ), .S(\SUMB[31][9] ) );
  FA_X1 S4_10 ( .A(\ab[31][10] ), .B(\CARRYB[30][10] ), .CI(\SUMB[30][11] ), 
        .CO(\CARRYB[31][10] ), .S(\SUMB[31][10] ) );
  FA_X1 S4_11 ( .A(\ab[31][11] ), .B(\CARRYB[30][11] ), .CI(\SUMB[30][12] ), 
        .CO(\CARRYB[31][11] ), .S(\SUMB[31][11] ) );
  FA_X1 S4_12 ( .A(\ab[31][12] ), .B(\CARRYB[30][12] ), .CI(\SUMB[30][13] ), 
        .CO(\CARRYB[31][12] ), .S(\SUMB[31][12] ) );
  FA_X1 S4_13 ( .A(\ab[31][13] ), .B(\CARRYB[30][13] ), .CI(\SUMB[30][14] ), 
        .CO(\CARRYB[31][13] ), .S(\SUMB[31][13] ) );
  FA_X1 S4_14 ( .A(\ab[31][14] ), .B(\CARRYB[30][14] ), .CI(\SUMB[30][15] ), 
        .CO(\CARRYB[31][14] ), .S(\SUMB[31][14] ) );
  FA_X1 S4_15 ( .A(\ab[31][15] ), .B(\CARRYB[30][15] ), .CI(\SUMB[30][16] ), 
        .CO(\CARRYB[31][15] ), .S(\SUMB[31][15] ) );
  FA_X1 S4_16 ( .A(\ab[31][16] ), .B(\CARRYB[30][16] ), .CI(\SUMB[30][17] ), 
        .CO(\CARRYB[31][16] ), .S(\SUMB[31][16] ) );
  FA_X1 S4_17 ( .A(\ab[31][17] ), .B(\CARRYB[30][17] ), .CI(\SUMB[30][18] ), 
        .CO(\CARRYB[31][17] ), .S(\SUMB[31][17] ) );
  FA_X1 S4_18 ( .A(\ab[31][18] ), .B(\CARRYB[30][18] ), .CI(\SUMB[30][19] ), 
        .CO(\CARRYB[31][18] ), .S(\SUMB[31][18] ) );
  FA_X1 S4_19 ( .A(\ab[31][19] ), .B(\CARRYB[30][19] ), .CI(\SUMB[30][20] ), 
        .CO(\CARRYB[31][19] ), .S(\SUMB[31][19] ) );
  FA_X1 S4_20 ( .A(\ab[31][20] ), .B(\CARRYB[30][20] ), .CI(\SUMB[30][21] ), 
        .CO(\CARRYB[31][20] ), .S(\SUMB[31][20] ) );
  FA_X1 S4_21 ( .A(\ab[31][21] ), .B(\CARRYB[30][21] ), .CI(\SUMB[30][22] ), 
        .CO(\CARRYB[31][21] ), .S(\SUMB[31][21] ) );
  FA_X1 S4_22 ( .A(\ab[31][22] ), .B(\CARRYB[30][22] ), .CI(\SUMB[30][23] ), 
        .CO(\CARRYB[31][22] ), .S(\SUMB[31][22] ) );
  FA_X1 S4_23 ( .A(\ab[31][23] ), .B(\CARRYB[30][23] ), .CI(\SUMB[30][24] ), 
        .CO(\CARRYB[31][23] ), .S(\SUMB[31][23] ) );
  FA_X1 S4_24 ( .A(\ab[31][24] ), .B(\CARRYB[30][24] ), .CI(\SUMB[30][25] ), 
        .CO(\CARRYB[31][24] ), .S(\SUMB[31][24] ) );
  FA_X1 S4_25 ( .A(\ab[31][25] ), .B(\CARRYB[30][25] ), .CI(\SUMB[30][26] ), 
        .CO(\CARRYB[31][25] ), .S(\SUMB[31][25] ) );
  FA_X1 S4_26 ( .A(\ab[31][26] ), .B(\CARRYB[30][26] ), .CI(\SUMB[30][27] ), 
        .CO(\CARRYB[31][26] ), .S(\SUMB[31][26] ) );
  FA_X1 S4_27 ( .A(\ab[31][27] ), .B(\CARRYB[30][27] ), .CI(\SUMB[30][28] ), 
        .CO(\CARRYB[31][27] ), .S(\SUMB[31][27] ) );
  FA_X1 S4_28 ( .A(\ab[31][28] ), .B(\CARRYB[30][28] ), .CI(\SUMB[30][29] ), 
        .CO(\CARRYB[31][28] ), .S(\SUMB[31][28] ) );
  FA_X1 S4_29 ( .A(\ab[31][29] ), .B(\CARRYB[30][29] ), .CI(\SUMB[30][30] ), 
        .CO(\CARRYB[31][29] ), .S(\SUMB[31][29] ) );
  FA_X1 S5_30 ( .A(\ab[31][30] ), .B(\CARRYB[30][30] ), .CI(\ab[30][31] ), 
        .CO(\CARRYB[31][30] ), .S(\SUMB[31][30] ) );
  FA_X1 S14_31 ( .A(n126), .B(n221), .CI(\ab[31][31] ), .CO(\CARRYB[31][31] ), 
        .S(\SUMB[31][31] ) );
  FA_X1 S1_30_0 ( .A(\ab[30][0] ), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), 
        .CO(\CARRYB[30][0] ), .S(\A1[28] ) );
  FA_X1 S2_30_1 ( .A(\ab[30][1] ), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), 
        .CO(\CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FA_X1 S2_30_2 ( .A(\ab[30][2] ), .B(\CARRYB[29][2] ), .CI(\SUMB[29][3] ), 
        .CO(\CARRYB[30][2] ), .S(\SUMB[30][2] ) );
  FA_X1 S2_30_3 ( .A(\ab[30][3] ), .B(\CARRYB[29][3] ), .CI(\SUMB[29][4] ), 
        .CO(\CARRYB[30][3] ), .S(\SUMB[30][3] ) );
  FA_X1 S2_30_4 ( .A(\ab[30][4] ), .B(\CARRYB[29][4] ), .CI(\SUMB[29][5] ), 
        .CO(\CARRYB[30][4] ), .S(\SUMB[30][4] ) );
  FA_X1 S2_30_5 ( .A(\ab[30][5] ), .B(\CARRYB[29][5] ), .CI(\SUMB[29][6] ), 
        .CO(\CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FA_X1 S2_30_6 ( .A(\ab[30][6] ), .B(\CARRYB[29][6] ), .CI(\SUMB[29][7] ), 
        .CO(\CARRYB[30][6] ), .S(\SUMB[30][6] ) );
  FA_X1 S2_30_7 ( .A(\ab[30][7] ), .B(\CARRYB[29][7] ), .CI(\SUMB[29][8] ), 
        .CO(\CARRYB[30][7] ), .S(\SUMB[30][7] ) );
  FA_X1 S2_30_8 ( .A(\ab[30][8] ), .B(\CARRYB[29][8] ), .CI(\SUMB[29][9] ), 
        .CO(\CARRYB[30][8] ), .S(\SUMB[30][8] ) );
  FA_X1 S2_30_9 ( .A(\ab[30][9] ), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), 
        .CO(\CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FA_X1 S2_30_10 ( .A(\ab[30][10] ), .B(\CARRYB[29][10] ), .CI(\SUMB[29][11] ), 
        .CO(\CARRYB[30][10] ), .S(\SUMB[30][10] ) );
  FA_X1 S2_30_11 ( .A(\ab[30][11] ), .B(\CARRYB[29][11] ), .CI(\SUMB[29][12] ), 
        .CO(\CARRYB[30][11] ), .S(\SUMB[30][11] ) );
  FA_X1 S2_30_12 ( .A(\ab[30][12] ), .B(\CARRYB[29][12] ), .CI(\SUMB[29][13] ), 
        .CO(\CARRYB[30][12] ), .S(\SUMB[30][12] ) );
  FA_X1 S2_30_13 ( .A(\ab[30][13] ), .B(\CARRYB[29][13] ), .CI(\SUMB[29][14] ), 
        .CO(\CARRYB[30][13] ), .S(\SUMB[30][13] ) );
  FA_X1 S2_30_14 ( .A(\ab[30][14] ), .B(\CARRYB[29][14] ), .CI(\SUMB[29][15] ), 
        .CO(\CARRYB[30][14] ), .S(\SUMB[30][14] ) );
  FA_X1 S2_30_15 ( .A(\ab[30][15] ), .B(\CARRYB[29][15] ), .CI(\SUMB[29][16] ), 
        .CO(\CARRYB[30][15] ), .S(\SUMB[30][15] ) );
  FA_X1 S2_30_16 ( .A(\ab[30][16] ), .B(\CARRYB[29][16] ), .CI(\SUMB[29][17] ), 
        .CO(\CARRYB[30][16] ), .S(\SUMB[30][16] ) );
  FA_X1 S2_30_17 ( .A(\ab[30][17] ), .B(\CARRYB[29][17] ), .CI(\SUMB[29][18] ), 
        .CO(\CARRYB[30][17] ), .S(\SUMB[30][17] ) );
  FA_X1 S2_30_18 ( .A(\ab[30][18] ), .B(\CARRYB[29][18] ), .CI(\SUMB[29][19] ), 
        .CO(\CARRYB[30][18] ), .S(\SUMB[30][18] ) );
  FA_X1 S2_30_19 ( .A(\ab[30][19] ), .B(\CARRYB[29][19] ), .CI(\SUMB[29][20] ), 
        .CO(\CARRYB[30][19] ), .S(\SUMB[30][19] ) );
  FA_X1 S2_30_20 ( .A(\ab[30][20] ), .B(\CARRYB[29][20] ), .CI(\SUMB[29][21] ), 
        .CO(\CARRYB[30][20] ), .S(\SUMB[30][20] ) );
  FA_X1 S2_30_21 ( .A(\ab[30][21] ), .B(\CARRYB[29][21] ), .CI(\SUMB[29][22] ), 
        .CO(\CARRYB[30][21] ), .S(\SUMB[30][21] ) );
  FA_X1 S2_30_22 ( .A(\ab[30][22] ), .B(\CARRYB[29][22] ), .CI(\SUMB[29][23] ), 
        .CO(\CARRYB[30][22] ), .S(\SUMB[30][22] ) );
  FA_X1 S2_30_23 ( .A(\ab[30][23] ), .B(\CARRYB[29][23] ), .CI(\SUMB[29][24] ), 
        .CO(\CARRYB[30][23] ), .S(\SUMB[30][23] ) );
  FA_X1 S2_30_24 ( .A(\ab[30][24] ), .B(\CARRYB[29][24] ), .CI(\SUMB[29][25] ), 
        .CO(\CARRYB[30][24] ), .S(\SUMB[30][24] ) );
  FA_X1 S2_30_25 ( .A(\ab[30][25] ), .B(\CARRYB[29][25] ), .CI(\SUMB[29][26] ), 
        .CO(\CARRYB[30][25] ), .S(\SUMB[30][25] ) );
  FA_X1 S2_30_26 ( .A(\ab[30][26] ), .B(\CARRYB[29][26] ), .CI(\SUMB[29][27] ), 
        .CO(\CARRYB[30][26] ), .S(\SUMB[30][26] ) );
  FA_X1 S2_30_27 ( .A(\ab[30][27] ), .B(\CARRYB[29][27] ), .CI(\SUMB[29][28] ), 
        .CO(\CARRYB[30][27] ), .S(\SUMB[30][27] ) );
  FA_X1 S2_30_28 ( .A(\ab[30][28] ), .B(\CARRYB[29][28] ), .CI(\SUMB[29][29] ), 
        .CO(\CARRYB[30][28] ), .S(\SUMB[30][28] ) );
  FA_X1 S2_30_29 ( .A(\ab[30][29] ), .B(\CARRYB[29][29] ), .CI(\SUMB[29][30] ), 
        .CO(\CARRYB[30][29] ), .S(\SUMB[30][29] ) );
  FA_X1 S3_30_30 ( .A(\ab[30][30] ), .B(\CARRYB[29][30] ), .CI(\ab[29][31] ), 
        .CO(\CARRYB[30][30] ), .S(\SUMB[30][30] ) );
  FA_X1 S1_29_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), 
        .CO(\CARRYB[29][0] ), .S(\A1[27] ) );
  FA_X1 S2_29_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), 
        .CO(\CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA_X1 S2_29_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), 
        .CO(\CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA_X1 S2_29_3 ( .A(\ab[29][3] ), .B(\CARRYB[28][3] ), .CI(\SUMB[28][4] ), 
        .CO(\CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA_X1 S2_29_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), 
        .CO(\CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA_X1 S2_29_5 ( .A(\ab[29][5] ), .B(\CARRYB[28][5] ), .CI(\SUMB[28][6] ), 
        .CO(\CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA_X1 S2_29_6 ( .A(\ab[29][6] ), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), 
        .CO(\CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA_X1 S2_29_7 ( .A(\ab[29][7] ), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), 
        .CO(\CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA_X1 S2_29_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), 
        .CO(\CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA_X1 S2_29_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), 
        .CO(\CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA_X1 S2_29_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), 
        .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA_X1 S2_29_11 ( .A(\ab[29][11] ), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), 
        .CO(\CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA_X1 S2_29_12 ( .A(\ab[29][12] ), .B(\CARRYB[28][12] ), .CI(\SUMB[28][13] ), 
        .CO(\CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA_X1 S2_29_13 ( .A(\ab[29][13] ), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), 
        .CO(\CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA_X1 S2_29_14 ( .A(\ab[29][14] ), .B(\CARRYB[28][14] ), .CI(\SUMB[28][15] ), 
        .CO(\CARRYB[29][14] ), .S(\SUMB[29][14] ) );
  FA_X1 S2_29_15 ( .A(\ab[29][15] ), .B(\CARRYB[28][15] ), .CI(\SUMB[28][16] ), 
        .CO(\CARRYB[29][15] ), .S(\SUMB[29][15] ) );
  FA_X1 S2_29_16 ( .A(\ab[29][16] ), .B(\CARRYB[28][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA_X1 S2_29_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA_X1 S2_29_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA_X1 S2_29_19 ( .A(\ab[29][19] ), .B(\CARRYB[28][19] ), .CI(\SUMB[28][20] ), 
        .CO(\CARRYB[29][19] ), .S(\SUMB[29][19] ) );
  FA_X1 S2_29_20 ( .A(\ab[29][20] ), .B(\CARRYB[28][20] ), .CI(\SUMB[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA_X1 S2_29_21 ( .A(\ab[29][21] ), .B(\CARRYB[28][21] ), .CI(\SUMB[28][22] ), 
        .CO(\CARRYB[29][21] ), .S(\SUMB[29][21] ) );
  FA_X1 S2_29_22 ( .A(\ab[29][22] ), .B(\CARRYB[28][22] ), .CI(\SUMB[28][23] ), 
        .CO(\CARRYB[29][22] ), .S(\SUMB[29][22] ) );
  FA_X1 S2_29_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), 
        .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FA_X1 S2_29_24 ( .A(\ab[29][24] ), .B(\CARRYB[28][24] ), .CI(\SUMB[28][25] ), 
        .CO(\CARRYB[29][24] ), .S(\SUMB[29][24] ) );
  FA_X1 S2_29_25 ( .A(\ab[29][25] ), .B(\CARRYB[28][25] ), .CI(\SUMB[28][26] ), 
        .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FA_X1 S2_29_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), 
        .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FA_X1 S2_29_27 ( .A(\ab[29][27] ), .B(\CARRYB[28][27] ), .CI(\SUMB[28][28] ), 
        .CO(\CARRYB[29][27] ), .S(\SUMB[29][27] ) );
  FA_X1 S2_29_28 ( .A(\ab[29][28] ), .B(\CARRYB[28][28] ), .CI(\SUMB[28][29] ), 
        .CO(\CARRYB[29][28] ), .S(\SUMB[29][28] ) );
  FA_X1 S2_29_29 ( .A(\ab[29][29] ), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), 
        .CO(\CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FA_X1 S3_29_30 ( .A(\ab[29][30] ), .B(\CARRYB[28][30] ), .CI(\ab[28][31] ), 
        .CO(\CARRYB[29][30] ), .S(\SUMB[29][30] ) );
  FA_X1 S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(\A1[26] ) );
  FA_X1 S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA_X1 S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA_X1 S2_28_3 ( .A(\ab[28][3] ), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), 
        .CO(\CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA_X1 S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA_X1 S2_28_5 ( .A(\ab[28][5] ), .B(\CARRYB[27][5] ), .CI(\SUMB[27][6] ), 
        .CO(\CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA_X1 S2_28_6 ( .A(\ab[28][6] ), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), 
        .CO(\CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA_X1 S2_28_7 ( .A(\ab[28][7] ), .B(\CARRYB[27][7] ), .CI(\SUMB[27][8] ), 
        .CO(\CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA_X1 S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA_X1 S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA_X1 S2_28_10 ( .A(\ab[28][10] ), .B(\CARRYB[27][10] ), .CI(\SUMB[27][11] ), 
        .CO(\CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA_X1 S2_28_11 ( .A(\ab[28][11] ), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), 
        .CO(\CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FA_X1 S2_28_12 ( .A(\ab[28][12] ), .B(\CARRYB[27][12] ), .CI(\SUMB[27][13] ), 
        .CO(\CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA_X1 S2_28_13 ( .A(\ab[28][13] ), .B(\CARRYB[27][13] ), .CI(\SUMB[27][14] ), 
        .CO(\CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA_X1 S2_28_14 ( .A(\ab[28][14] ), .B(\CARRYB[27][14] ), .CI(\SUMB[27][15] ), 
        .CO(\CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA_X1 S2_28_15 ( .A(\ab[28][15] ), .B(\CARRYB[27][15] ), .CI(\SUMB[27][16] ), 
        .CO(\CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA_X1 S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA_X1 S2_28_17 ( .A(\ab[28][17] ), .B(\CARRYB[27][17] ), .CI(\SUMB[27][18] ), 
        .CO(\CARRYB[28][17] ), .S(\SUMB[28][17] ) );
  FA_X1 S2_28_18 ( .A(\ab[28][18] ), .B(\CARRYB[27][18] ), .CI(\SUMB[27][19] ), 
        .CO(\CARRYB[28][18] ), .S(\SUMB[28][18] ) );
  FA_X1 S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA_X1 S2_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\SUMB[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA_X1 S2_28_21 ( .A(\ab[28][21] ), .B(\CARRYB[27][21] ), .CI(\SUMB[27][22] ), 
        .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FA_X1 S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), 
        .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FA_X1 S2_28_23 ( .A(\ab[28][23] ), .B(\CARRYB[27][23] ), .CI(\SUMB[27][24] ), 
        .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FA_X1 S2_28_24 ( .A(\ab[28][24] ), .B(\CARRYB[27][24] ), .CI(\SUMB[27][25] ), 
        .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FA_X1 S2_28_25 ( .A(\ab[28][25] ), .B(\CARRYB[27][25] ), .CI(\SUMB[27][26] ), 
        .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FA_X1 S2_28_26 ( .A(\ab[28][26] ), .B(\CARRYB[27][26] ), .CI(\SUMB[27][27] ), 
        .CO(\CARRYB[28][26] ), .S(\SUMB[28][26] ) );
  FA_X1 S2_28_27 ( .A(\ab[28][27] ), .B(\CARRYB[27][27] ), .CI(\SUMB[27][28] ), 
        .CO(\CARRYB[28][27] ), .S(\SUMB[28][27] ) );
  FA_X1 S2_28_28 ( .A(\ab[28][28] ), .B(\CARRYB[27][28] ), .CI(\SUMB[27][29] ), 
        .CO(\CARRYB[28][28] ), .S(\SUMB[28][28] ) );
  FA_X1 S2_28_29 ( .A(\ab[28][29] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), 
        .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FA_X1 S3_28_30 ( .A(\ab[28][30] ), .B(\CARRYB[27][30] ), .CI(\ab[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FA_X1 S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(\A1[25] ) );
  FA_X1 S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA_X1 S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA_X1 S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA_X1 S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA_X1 S2_27_5 ( .A(\ab[27][5] ), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), 
        .CO(\CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA_X1 S2_27_6 ( .A(\ab[27][6] ), .B(\CARRYB[26][6] ), .CI(\SUMB[26][7] ), 
        .CO(\CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA_X1 S2_27_7 ( .A(\ab[27][7] ), .B(\CARRYB[26][7] ), .CI(\SUMB[26][8] ), 
        .CO(\CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA_X1 S2_27_8 ( .A(\ab[27][8] ), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA_X1 S2_27_9 ( .A(\ab[27][9] ), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), 
        .CO(\CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA_X1 S2_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), 
        .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA_X1 S2_27_11 ( .A(\ab[27][11] ), .B(\CARRYB[26][11] ), .CI(\SUMB[26][12] ), 
        .CO(\CARRYB[27][11] ), .S(\SUMB[27][11] ) );
  FA_X1 S2_27_12 ( .A(\ab[27][12] ), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), 
        .CO(\CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA_X1 S2_27_13 ( .A(\ab[27][13] ), .B(\CARRYB[26][13] ), .CI(\SUMB[26][14] ), 
        .CO(\CARRYB[27][13] ), .S(\SUMB[27][13] ) );
  FA_X1 S2_27_14 ( .A(\ab[27][14] ), .B(\CARRYB[26][14] ), .CI(\SUMB[26][15] ), 
        .CO(\CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA_X1 S2_27_15 ( .A(\ab[27][15] ), .B(\CARRYB[26][15] ), .CI(\SUMB[26][16] ), 
        .CO(\CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA_X1 S2_27_16 ( .A(\ab[27][16] ), .B(\CARRYB[26][16] ), .CI(\SUMB[26][17] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA_X1 S2_27_17 ( .A(\ab[27][17] ), .B(\CARRYB[26][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA_X1 S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA_X1 S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA_X1 S2_27_20 ( .A(\ab[27][20] ), .B(\CARRYB[26][20] ), .CI(\SUMB[26][21] ), 
        .CO(\CARRYB[27][20] ), .S(\SUMB[27][20] ) );
  FA_X1 S2_27_21 ( .A(\ab[27][21] ), .B(\CARRYB[26][21] ), .CI(\SUMB[26][22] ), 
        .CO(\CARRYB[27][21] ), .S(\SUMB[27][21] ) );
  FA_X1 S2_27_22 ( .A(\ab[27][22] ), .B(\CARRYB[26][22] ), .CI(\SUMB[26][23] ), 
        .CO(\CARRYB[27][22] ), .S(\SUMB[27][22] ) );
  FA_X1 S2_27_23 ( .A(\ab[27][23] ), .B(\CARRYB[26][23] ), .CI(\SUMB[26][24] ), 
        .CO(\CARRYB[27][23] ), .S(\SUMB[27][23] ) );
  FA_X1 S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), 
        .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FA_X1 S2_27_25 ( .A(\ab[27][25] ), .B(\CARRYB[26][25] ), .CI(\SUMB[26][26] ), 
        .CO(\CARRYB[27][25] ), .S(\SUMB[27][25] ) );
  FA_X1 S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), 
        .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FA_X1 S2_27_27 ( .A(\ab[27][27] ), .B(\CARRYB[26][27] ), .CI(\SUMB[26][28] ), 
        .CO(\CARRYB[27][27] ), .S(\SUMB[27][27] ) );
  FA_X1 S2_27_28 ( .A(\ab[27][28] ), .B(\CARRYB[26][28] ), .CI(\SUMB[26][29] ), 
        .CO(\CARRYB[27][28] ), .S(\SUMB[27][28] ) );
  FA_X1 S2_27_29 ( .A(\ab[27][29] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), 
        .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FA_X1 S3_27_30 ( .A(\ab[27][30] ), .B(\CARRYB[26][30] ), .CI(\ab[26][31] ), 
        .CO(\CARRYB[27][30] ), .S(\SUMB[27][30] ) );
  FA_X1 S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(\A1[24] ) );
  FA_X1 S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA_X1 S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA_X1 S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA_X1 S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA_X1 S2_26_5 ( .A(\ab[26][5] ), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), 
        .CO(\CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA_X1 S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA_X1 S2_26_7 ( .A(\ab[26][7] ), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA_X1 S2_26_8 ( .A(\ab[26][8] ), .B(\CARRYB[25][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA_X1 S2_26_9 ( .A(\ab[26][9] ), .B(\CARRYB[25][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA_X1 S2_26_10 ( .A(\ab[26][10] ), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), 
        .CO(\CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA_X1 S2_26_11 ( .A(\ab[26][11] ), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), 
        .CO(\CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA_X1 S2_26_12 ( .A(\ab[26][12] ), .B(\CARRYB[25][12] ), .CI(\SUMB[25][13] ), 
        .CO(\CARRYB[26][12] ), .S(\SUMB[26][12] ) );
  FA_X1 S2_26_13 ( .A(\ab[26][13] ), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), 
        .CO(\CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA_X1 S2_26_14 ( .A(\ab[26][14] ), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), 
        .CO(\CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA_X1 S2_26_15 ( .A(\ab[26][15] ), .B(\CARRYB[25][15] ), .CI(\SUMB[25][16] ), 
        .CO(\CARRYB[26][15] ), .S(\SUMB[26][15] ) );
  FA_X1 S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA_X1 S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA_X1 S2_26_18 ( .A(\ab[26][18] ), .B(\CARRYB[25][18] ), .CI(\SUMB[25][19] ), 
        .CO(\CARRYB[26][18] ), .S(\SUMB[26][18] ) );
  FA_X1 S2_26_19 ( .A(\ab[26][19] ), .B(\CARRYB[25][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA_X1 S2_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\SUMB[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA_X1 S2_26_21 ( .A(\ab[26][21] ), .B(\CARRYB[25][21] ), .CI(\SUMB[25][22] ), 
        .CO(\CARRYB[26][21] ), .S(\SUMB[26][21] ) );
  FA_X1 S2_26_22 ( .A(\ab[26][22] ), .B(\CARRYB[25][22] ), .CI(\SUMB[25][23] ), 
        .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FA_X1 S2_26_23 ( .A(\ab[26][23] ), .B(\CARRYB[25][23] ), .CI(\SUMB[25][24] ), 
        .CO(\CARRYB[26][23] ), .S(\SUMB[26][23] ) );
  FA_X1 S2_26_24 ( .A(\ab[26][24] ), .B(\CARRYB[25][24] ), .CI(\SUMB[25][25] ), 
        .CO(\CARRYB[26][24] ), .S(\SUMB[26][24] ) );
  FA_X1 S2_26_25 ( .A(\ab[26][25] ), .B(\CARRYB[25][25] ), .CI(\SUMB[25][26] ), 
        .CO(\CARRYB[26][25] ), .S(\SUMB[26][25] ) );
  FA_X1 S2_26_26 ( .A(\ab[26][26] ), .B(\CARRYB[25][26] ), .CI(\SUMB[25][27] ), 
        .CO(\CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FA_X1 S2_26_27 ( .A(\ab[26][27] ), .B(\CARRYB[25][27] ), .CI(\SUMB[25][28] ), 
        .CO(\CARRYB[26][27] ), .S(\SUMB[26][27] ) );
  FA_X1 S2_26_28 ( .A(\ab[26][28] ), .B(\CARRYB[25][28] ), .CI(\SUMB[25][29] ), 
        .CO(\CARRYB[26][28] ), .S(\SUMB[26][28] ) );
  FA_X1 S2_26_29 ( .A(\ab[26][29] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), 
        .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FA_X1 S3_26_30 ( .A(\ab[26][30] ), .B(\CARRYB[25][30] ), .CI(\ab[25][31] ), 
        .CO(\CARRYB[26][30] ), .S(\SUMB[26][30] ) );
  FA_X1 S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(\A1[23] ) );
  FA_X1 S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA_X1 S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA_X1 S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA_X1 S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA_X1 S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA_X1 S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA_X1 S2_25_7 ( .A(\ab[25][7] ), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA_X1 S2_25_8 ( .A(\ab[25][8] ), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA_X1 S2_25_9 ( .A(\ab[25][9] ), .B(\CARRYB[24][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA_X1 S2_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), 
        .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA_X1 S2_25_11 ( .A(\ab[25][11] ), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), 
        .CO(\CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA_X1 S2_25_12 ( .A(\ab[25][12] ), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), 
        .CO(\CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA_X1 S2_25_13 ( .A(\ab[25][13] ), .B(\CARRYB[24][13] ), .CI(\SUMB[24][14] ), 
        .CO(\CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA_X1 S2_25_14 ( .A(\ab[25][14] ), .B(\CARRYB[24][14] ), .CI(\SUMB[24][15] ), 
        .CO(\CARRYB[25][14] ), .S(\SUMB[25][14] ) );
  FA_X1 S2_25_15 ( .A(\ab[25][15] ), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), 
        .CO(\CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA_X1 S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), 
        .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FA_X1 S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FA_X1 S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA_X1 S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA_X1 S2_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\SUMB[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA_X1 S2_25_21 ( .A(\ab[25][21] ), .B(\CARRYB[24][21] ), .CI(\SUMB[24][22] ), 
        .CO(\CARRYB[25][21] ), .S(\SUMB[25][21] ) );
  FA_X1 S2_25_22 ( .A(\ab[25][22] ), .B(\CARRYB[24][22] ), .CI(\SUMB[24][23] ), 
        .CO(\CARRYB[25][22] ), .S(\SUMB[25][22] ) );
  FA_X1 S2_25_23 ( .A(\ab[25][23] ), .B(\CARRYB[24][23] ), .CI(\SUMB[24][24] ), 
        .CO(\CARRYB[25][23] ), .S(\SUMB[25][23] ) );
  FA_X1 S2_25_24 ( .A(\ab[25][24] ), .B(\CARRYB[24][24] ), .CI(\SUMB[24][25] ), 
        .CO(\CARRYB[25][24] ), .S(\SUMB[25][24] ) );
  FA_X1 S2_25_25 ( .A(\ab[25][25] ), .B(\CARRYB[24][25] ), .CI(\SUMB[24][26] ), 
        .CO(\CARRYB[25][25] ), .S(\SUMB[25][25] ) );
  FA_X1 S2_25_26 ( .A(\ab[25][26] ), .B(\CARRYB[24][26] ), .CI(\SUMB[24][27] ), 
        .CO(\CARRYB[25][26] ), .S(\SUMB[25][26] ) );
  FA_X1 S2_25_27 ( .A(\ab[25][27] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), 
        .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FA_X1 S2_25_28 ( .A(\ab[25][28] ), .B(\CARRYB[24][28] ), .CI(\SUMB[24][29] ), 
        .CO(\CARRYB[25][28] ), .S(\SUMB[25][28] ) );
  FA_X1 S2_25_29 ( .A(\ab[25][29] ), .B(\CARRYB[24][29] ), .CI(\SUMB[24][30] ), 
        .CO(\CARRYB[25][29] ), .S(\SUMB[25][29] ) );
  FA_X1 S3_25_30 ( .A(\ab[25][30] ), .B(\CARRYB[24][30] ), .CI(\ab[24][31] ), 
        .CO(\CARRYB[25][30] ), .S(\SUMB[25][30] ) );
  FA_X1 S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(\A1[22] ) );
  FA_X1 S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA_X1 S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA_X1 S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA_X1 S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA_X1 S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA_X1 S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA_X1 S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA_X1 S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA_X1 S2_24_9 ( .A(\ab[24][9] ), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA_X1 S2_24_10 ( .A(\ab[24][10] ), .B(\CARRYB[23][10] ), .CI(\SUMB[23][11] ), 
        .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA_X1 S2_24_11 ( .A(\ab[24][11] ), .B(\CARRYB[23][11] ), .CI(\SUMB[23][12] ), 
        .CO(\CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FA_X1 S2_24_12 ( .A(\ab[24][12] ), .B(\CARRYB[23][12] ), .CI(\SUMB[23][13] ), 
        .CO(\CARRYB[24][12] ), .S(\SUMB[24][12] ) );
  FA_X1 S2_24_13 ( .A(\ab[24][13] ), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), 
        .CO(\CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA_X1 S2_24_14 ( .A(\ab[24][14] ), .B(\CARRYB[23][14] ), .CI(\SUMB[23][15] ), 
        .CO(\CARRYB[24][14] ), .S(\SUMB[24][14] ) );
  FA_X1 S2_24_15 ( .A(\ab[24][15] ), .B(\CARRYB[23][15] ), .CI(\SUMB[23][16] ), 
        .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA_X1 S2_24_16 ( .A(\ab[24][16] ), .B(\CARRYB[23][16] ), .CI(\SUMB[23][17] ), 
        .CO(\CARRYB[24][16] ), .S(\SUMB[24][16] ) );
  FA_X1 S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA_X1 S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA_X1 S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA_X1 S2_24_20 ( .A(\ab[24][20] ), .B(\CARRYB[23][20] ), .CI(\SUMB[23][21] ), 
        .CO(\CARRYB[24][20] ), .S(\SUMB[24][20] ) );
  FA_X1 S2_24_21 ( .A(\ab[24][21] ), .B(\CARRYB[23][21] ), .CI(\SUMB[23][22] ), 
        .CO(\CARRYB[24][21] ), .S(\SUMB[24][21] ) );
  FA_X1 S2_24_22 ( .A(\ab[24][22] ), .B(\CARRYB[23][22] ), .CI(\SUMB[23][23] ), 
        .CO(\CARRYB[24][22] ), .S(\SUMB[24][22] ) );
  FA_X1 S2_24_23 ( .A(\ab[24][23] ), .B(\CARRYB[23][23] ), .CI(\SUMB[23][24] ), 
        .CO(\CARRYB[24][23] ), .S(\SUMB[24][23] ) );
  FA_X1 S2_24_24 ( .A(\ab[24][24] ), .B(\CARRYB[23][24] ), .CI(\SUMB[23][25] ), 
        .CO(\CARRYB[24][24] ), .S(\SUMB[24][24] ) );
  FA_X1 S2_24_25 ( .A(\ab[24][25] ), .B(\CARRYB[23][25] ), .CI(\SUMB[23][26] ), 
        .CO(\CARRYB[24][25] ), .S(\SUMB[24][25] ) );
  FA_X1 S2_24_26 ( .A(\ab[24][26] ), .B(\CARRYB[23][26] ), .CI(\SUMB[23][27] ), 
        .CO(\CARRYB[24][26] ), .S(\SUMB[24][26] ) );
  FA_X1 S2_24_27 ( .A(\ab[24][27] ), .B(\CARRYB[23][27] ), .CI(\SUMB[23][28] ), 
        .CO(\CARRYB[24][27] ), .S(\SUMB[24][27] ) );
  FA_X1 S2_24_28 ( .A(\ab[24][28] ), .B(\CARRYB[23][28] ), .CI(\SUMB[23][29] ), 
        .CO(\CARRYB[24][28] ), .S(\SUMB[24][28] ) );
  FA_X1 S2_24_29 ( .A(\ab[24][29] ), .B(\CARRYB[23][29] ), .CI(\SUMB[23][30] ), 
        .CO(\CARRYB[24][29] ), .S(\SUMB[24][29] ) );
  FA_X1 S3_24_30 ( .A(\ab[24][30] ), .B(\CARRYB[23][30] ), .CI(\ab[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FA_X1 S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(\A1[21] ) );
  FA_X1 S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA_X1 S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA_X1 S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA_X1 S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA_X1 S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA_X1 S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA_X1 S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA_X1 S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA_X1 S2_23_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA_X1 S2_23_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA_X1 S2_23_11 ( .A(\ab[23][11] ), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA_X1 S2_23_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA_X1 S2_23_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA_X1 S2_23_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA_X1 S2_23_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA_X1 S2_23_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA_X1 S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA_X1 S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA_X1 S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA_X1 S2_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA_X1 S2_23_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA_X1 S2_23_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\SUMB[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA_X1 S2_23_23 ( .A(\ab[23][23] ), .B(\CARRYB[22][23] ), .CI(\SUMB[22][24] ), 
        .CO(\CARRYB[23][23] ), .S(\SUMB[23][23] ) );
  FA_X1 S2_23_24 ( .A(\ab[23][24] ), .B(\CARRYB[22][24] ), .CI(\SUMB[22][25] ), 
        .CO(\CARRYB[23][24] ), .S(\SUMB[23][24] ) );
  FA_X1 S2_23_25 ( .A(\ab[23][25] ), .B(\CARRYB[22][25] ), .CI(\SUMB[22][26] ), 
        .CO(\CARRYB[23][25] ), .S(\SUMB[23][25] ) );
  FA_X1 S2_23_26 ( .A(\ab[23][26] ), .B(\CARRYB[22][26] ), .CI(\SUMB[22][27] ), 
        .CO(\CARRYB[23][26] ), .S(\SUMB[23][26] ) );
  FA_X1 S2_23_27 ( .A(\ab[23][27] ), .B(\CARRYB[22][27] ), .CI(\SUMB[22][28] ), 
        .CO(\CARRYB[23][27] ), .S(\SUMB[23][27] ) );
  FA_X1 S2_23_28 ( .A(\ab[23][28] ), .B(\CARRYB[22][28] ), .CI(\SUMB[22][29] ), 
        .CO(\CARRYB[23][28] ), .S(\SUMB[23][28] ) );
  FA_X1 S2_23_29 ( .A(\ab[23][29] ), .B(\CARRYB[22][29] ), .CI(\SUMB[22][30] ), 
        .CO(\CARRYB[23][29] ), .S(\SUMB[23][29] ) );
  FA_X1 S3_23_30 ( .A(\ab[23][30] ), .B(\CARRYB[22][30] ), .CI(\ab[22][31] ), 
        .CO(\CARRYB[23][30] ), .S(\SUMB[23][30] ) );
  FA_X1 S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FA_X1 S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA_X1 S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA_X1 S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA_X1 S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA_X1 S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA_X1 S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA_X1 S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA_X1 S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA_X1 S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA_X1 S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA_X1 S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), 
        .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA_X1 S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), 
        .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA_X1 S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(\SUMB[21][14] ), 
        .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FA_X1 S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), 
        .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA_X1 S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA_X1 S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA_X1 S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA_X1 S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA_X1 S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA_X1 S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA_X1 S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA_X1 S2_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), 
        .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA_X1 S2_22_23 ( .A(\ab[22][23] ), .B(\CARRYB[21][23] ), .CI(\SUMB[21][24] ), 
        .CO(\CARRYB[22][23] ), .S(\SUMB[22][23] ) );
  FA_X1 S2_22_24 ( .A(\ab[22][24] ), .B(\CARRYB[21][24] ), .CI(\SUMB[21][25] ), 
        .CO(\CARRYB[22][24] ), .S(\SUMB[22][24] ) );
  FA_X1 S2_22_25 ( .A(\ab[22][25] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), 
        .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FA_X1 S2_22_26 ( .A(\ab[22][26] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), 
        .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FA_X1 S2_22_27 ( .A(\ab[22][27] ), .B(\CARRYB[21][27] ), .CI(\SUMB[21][28] ), 
        .CO(\CARRYB[22][27] ), .S(\SUMB[22][27] ) );
  FA_X1 S2_22_28 ( .A(\ab[22][28] ), .B(\CARRYB[21][28] ), .CI(\SUMB[21][29] ), 
        .CO(\CARRYB[22][28] ), .S(\SUMB[22][28] ) );
  FA_X1 S2_22_29 ( .A(\ab[22][29] ), .B(\CARRYB[21][29] ), .CI(\SUMB[21][30] ), 
        .CO(\CARRYB[22][29] ), .S(\SUMB[22][29] ) );
  FA_X1 S3_22_30 ( .A(\ab[22][30] ), .B(\CARRYB[21][30] ), .CI(\ab[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FA_X1 S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FA_X1 S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA_X1 S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA_X1 S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA_X1 S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA_X1 S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA_X1 S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA_X1 S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA_X1 S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA_X1 S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA_X1 S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA_X1 S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA_X1 S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA_X1 S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA_X1 S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA_X1 S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA_X1 S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA_X1 S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA_X1 S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA_X1 S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA_X1 S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA_X1 S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA_X1 S2_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA_X1 S2_21_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA_X1 S2_21_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA_X1 S2_21_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA_X1 S2_21_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA_X1 S2_21_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA_X1 S2_21_28 ( .A(\ab[21][28] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA_X1 S2_21_29 ( .A(\ab[21][29] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA_X1 S3_21_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\ab[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA_X1 S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA_X1 S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA_X1 S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA_X1 S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA_X1 S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA_X1 S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA_X1 S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA_X1 S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA_X1 S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA_X1 S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA_X1 S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA_X1 S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA_X1 S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA_X1 S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA_X1 S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA_X1 S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA_X1 S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA_X1 S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA_X1 S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA_X1 S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA_X1 S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA_X1 S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA_X1 S2_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA_X1 S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA_X1 S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA_X1 S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA_X1 S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA_X1 S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA_X1 S2_20_28 ( .A(\ab[20][28] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA_X1 S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA_X1 S3_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\ab[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA_X1 S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA_X1 S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA_X1 S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA_X1 S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA_X1 S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA_X1 S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA_X1 S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA_X1 S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA_X1 S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA_X1 S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA_X1 S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA_X1 S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA_X1 S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA_X1 S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA_X1 S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA_X1 S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA_X1 S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA_X1 S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA_X1 S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA_X1 S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA_X1 S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA_X1 S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA_X1 S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA_X1 S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA_X1 S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA_X1 S2_19_25 ( .A(\ab[19][25] ), .B(\CARRYB[18][25] ), .CI(\SUMB[18][26] ), 
        .CO(\CARRYB[19][25] ), .S(\SUMB[19][25] ) );
  FA_X1 S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA_X1 S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA_X1 S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA_X1 S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA_X1 S3_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\ab[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA_X1 S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA_X1 S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA_X1 S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA_X1 S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA_X1 S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA_X1 S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA_X1 S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA_X1 S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA_X1 S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA_X1 S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA_X1 S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA_X1 S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA_X1 S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA_X1 S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA_X1 S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA_X1 S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA_X1 S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA_X1 S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA_X1 S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA_X1 S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA_X1 S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA_X1 S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA_X1 S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA_X1 S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA_X1 S2_18_24 ( .A(\ab[18][24] ), .B(\CARRYB[17][24] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA_X1 S2_18_25 ( .A(\ab[18][25] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA_X1 S2_18_26 ( .A(\ab[18][26] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA_X1 S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA_X1 S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA_X1 S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA_X1 S3_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\ab[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA_X1 S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA_X1 S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA_X1 S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA_X1 S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA_X1 S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA_X1 S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA_X1 S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA_X1 S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA_X1 S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA_X1 S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA_X1 S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA_X1 S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA_X1 S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA_X1 S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA_X1 S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA_X1 S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA_X1 S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA_X1 S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA_X1 S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA_X1 S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA_X1 S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA_X1 S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA_X1 S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA_X1 S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA_X1 S2_17_24 ( .A(\ab[17][24] ), .B(\CARRYB[16][24] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA_X1 S2_17_25 ( .A(\ab[17][25] ), .B(\CARRYB[16][25] ), .CI(\SUMB[16][26] ), 
        .CO(\CARRYB[17][25] ), .S(\SUMB[17][25] ) );
  FA_X1 S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA_X1 S2_17_27 ( .A(\ab[17][27] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA_X1 S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA_X1 S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA_X1 S3_17_30 ( .A(\ab[17][30] ), .B(\CARRYB[16][30] ), .CI(\ab[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA_X1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA_X1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA_X1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA_X1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA_X1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA_X1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA_X1 S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA_X1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA_X1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA_X1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA_X1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA_X1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA_X1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA_X1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA_X1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA_X1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA_X1 S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA_X1 S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA_X1 S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA_X1 S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA_X1 S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA_X1 S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA_X1 S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA_X1 S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA_X1 S2_16_24 ( .A(\ab[16][24] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA_X1 S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA_X1 S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA_X1 S2_16_27 ( .A(\ab[16][27] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA_X1 S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA_X1 S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA_X1 S3_16_30 ( .A(\ab[16][30] ), .B(\CARRYB[15][30] ), .CI(\ab[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA_X1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA_X1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA_X1 S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA_X1 S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA_X1 S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA_X1 S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA_X1 S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA_X1 S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA_X1 S2_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA_X1 S2_15_23 ( .A(\ab[15][23] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA_X1 S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA_X1 S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA_X1 S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), 
        .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FA_X1 S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA_X1 S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA_X1 S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA_X1 S3_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\ab[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA_X1 S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA_X1 S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA_X1 S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA_X1 S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA_X1 S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA_X1 S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA_X1 S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA_X1 S2_14_23 ( .A(\ab[14][23] ), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), 
        .CO(\CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA_X1 S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), 
        .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA_X1 S2_14_25 ( .A(\ab[14][25] ), .B(\CARRYB[13][25] ), .CI(\SUMB[13][26] ), 
        .CO(\CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA_X1 S2_14_26 ( .A(\ab[14][26] ), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), 
        .CO(\CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA_X1 S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), 
        .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA_X1 S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA_X1 S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA_X1 S3_14_30 ( .A(\ab[14][30] ), .B(\CARRYB[13][30] ), .CI(\ab[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA_X1 S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA_X1 S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA_X1 S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA_X1 S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA_X1 S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA_X1 S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA_X1 S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA_X1 S2_13_23 ( .A(\ab[13][23] ), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), 
        .CO(\CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA_X1 S2_13_24 ( .A(\ab[13][24] ), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), 
        .CO(\CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA_X1 S2_13_25 ( .A(\ab[13][25] ), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), 
        .CO(\CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA_X1 S2_13_26 ( .A(\ab[13][26] ), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), 
        .CO(\CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA_X1 S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), 
        .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA_X1 S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), 
        .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA_X1 S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), 
        .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA_X1 S3_13_30 ( .A(\ab[13][30] ), .B(\CARRYB[12][30] ), .CI(\ab[12][31] ), 
        .CO(\CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA_X1 S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA_X1 S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA_X1 S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA_X1 S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA_X1 S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA_X1 S2_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\SUMB[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA_X1 S2_12_23 ( .A(\ab[12][23] ), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), 
        .CO(\CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA_X1 S2_12_24 ( .A(\ab[12][24] ), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), 
        .CO(\CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA_X1 S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), 
        .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA_X1 S2_12_26 ( .A(\ab[12][26] ), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), 
        .CO(\CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA_X1 S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), 
        .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA_X1 S2_12_28 ( .A(\ab[12][28] ), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), 
        .CO(\CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA_X1 S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), 
        .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA_X1 S3_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\ab[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA_X1 S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA_X1 S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA_X1 S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA_X1 S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA_X1 S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA_X1 S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA_X1 S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA_X1 S2_11_23 ( .A(\ab[11][23] ), .B(\CARRYB[10][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA_X1 S2_11_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA_X1 S2_11_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA_X1 S2_11_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA_X1 S2_11_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA_X1 S2_11_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA_X1 S2_11_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), 
        .CO(\CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA_X1 S3_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\ab[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA_X1 S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA_X1 S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA_X1 S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA_X1 S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA_X1 S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA_X1 S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA_X1 S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA_X1 S2_10_23 ( .A(\ab[10][23] ), .B(\CARRYB[9][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA_X1 S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA_X1 S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA_X1 S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA_X1 S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA_X1 S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA_X1 S2_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA_X1 S3_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\ab[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA_X1 S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA_X1 S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA_X1 S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA_X1 S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA_X1 S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA_X1 S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA_X1 S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA_X1 S2_9_23 ( .A(\ab[9][23] ), .B(\CARRYB[8][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA_X1 S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA_X1 S2_9_25 ( .A(\ab[9][25] ), .B(\CARRYB[8][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA_X1 S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA_X1 S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA_X1 S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA_X1 S2_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), 
        .CO(\CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA_X1 S3_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\ab[8][31] ), .CO(
        \CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA_X1 S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA_X1 S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA_X1 S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA_X1 S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA_X1 S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA_X1 S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA_X1 S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA_X1 S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA_X1 S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA_X1 S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA_X1 S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA_X1 S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA_X1 S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA_X1 S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA_X1 S3_8_30 ( .A(\ab[8][30] ), .B(\CARRYB[7][30] ), .CI(\ab[7][31] ), .CO(
        \CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA_X1 S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA_X1 S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA_X1 S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA_X1 S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA_X1 S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA_X1 S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA_X1 S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA_X1 S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA_X1 S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA_X1 S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA_X1 S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA_X1 S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA_X1 S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA_X1 S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA_X1 S3_7_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .CI(\ab[6][31] ), .CO(
        \CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA_X1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA_X1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA_X1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA_X1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA_X1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA_X1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA_X1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA_X1 S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA_X1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA_X1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA_X1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA_X1 S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA_X1 S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA_X1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA_X1 S3_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .CI(\ab[5][31] ), .CO(
        \CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA_X1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA_X1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA_X1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA_X1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA_X1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA_X1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA_X1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA_X1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA_X1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA_X1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA_X1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA_X1 S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA_X1 S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA_X1 S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\SUMB[4][30] ), 
        .CO(\CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA_X1 S3_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .CI(\ab[4][31] ), .CO(
        \CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA_X1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA_X1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA_X1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA_X1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA_X1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA_X1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA_X1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA_X1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA_X1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA_X1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA_X1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA_X1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA_X1 S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA_X1 S2_4_29 ( .A(\ab[4][29] ), .B(\CARRYB[3][29] ), .CI(\SUMB[3][30] ), 
        .CO(\CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA_X1 S3_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .CI(\ab[3][31] ), .CO(
        \CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA_X1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA_X1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA_X1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA_X1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA_X1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA_X1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA_X1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA_X1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA_X1 S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA_X1 S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA_X1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA_X1 S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA_X1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA_X1 S2_3_29 ( .A(\ab[3][29] ), .B(\CARRYB[2][29] ), .CI(\SUMB[2][30] ), 
        .CO(\CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA_X1 S3_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .CI(\ab[2][31] ), .CO(
        \CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n31), .CI(n62), .CO(\CARRYB[2][0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n30), .CI(n61), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n29), .CI(n60), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n28), .CI(n59), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n27), .CI(n58), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n26), .CI(n57), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n25), .CI(n56), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n24), .CI(n55), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n23), .CI(n54), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n22), .CI(n53), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n21), .CI(n52), .CO(\CARRYB[2][10] ), 
        .S(\SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n20), .CI(n51), .CO(\CARRYB[2][11] ), 
        .S(\SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n19), .CI(n50), .CO(\CARRYB[2][12] ), 
        .S(\SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n18), .CI(n49), .CO(\CARRYB[2][13] ), 
        .S(\SUMB[2][13] ) );
  FA_X1 S2_2_14 ( .A(\ab[2][14] ), .B(n17), .CI(n48), .CO(\CARRYB[2][14] ), 
        .S(\SUMB[2][14] ) );
  FA_X1 S2_2_15 ( .A(\ab[2][15] ), .B(n16), .CI(n47), .CO(\CARRYB[2][15] ), 
        .S(\SUMB[2][15] ) );
  FA_X1 S2_2_16 ( .A(\ab[2][16] ), .B(n15), .CI(n46), .CO(\CARRYB[2][16] ), 
        .S(\SUMB[2][16] ) );
  FA_X1 S2_2_17 ( .A(\ab[2][17] ), .B(n14), .CI(n45), .CO(\CARRYB[2][17] ), 
        .S(\SUMB[2][17] ) );
  FA_X1 S2_2_18 ( .A(\ab[2][18] ), .B(n13), .CI(n44), .CO(\CARRYB[2][18] ), 
        .S(\SUMB[2][18] ) );
  FA_X1 S2_2_19 ( .A(\ab[2][19] ), .B(n12), .CI(n43), .CO(\CARRYB[2][19] ), 
        .S(\SUMB[2][19] ) );
  FA_X1 S2_2_20 ( .A(\ab[2][20] ), .B(n11), .CI(n42), .CO(\CARRYB[2][20] ), 
        .S(\SUMB[2][20] ) );
  FA_X1 S2_2_21 ( .A(\ab[2][21] ), .B(n10), .CI(n41), .CO(\CARRYB[2][21] ), 
        .S(\SUMB[2][21] ) );
  FA_X1 S2_2_22 ( .A(\ab[2][22] ), .B(n9), .CI(n40), .CO(\CARRYB[2][22] ), .S(
        \SUMB[2][22] ) );
  FA_X1 S2_2_23 ( .A(\ab[2][23] ), .B(n8), .CI(n39), .CO(\CARRYB[2][23] ), .S(
        \SUMB[2][23] ) );
  FA_X1 S2_2_24 ( .A(\ab[2][24] ), .B(n7), .CI(n38), .CO(\CARRYB[2][24] ), .S(
        \SUMB[2][24] ) );
  FA_X1 S2_2_25 ( .A(\ab[2][25] ), .B(n6), .CI(n37), .CO(\CARRYB[2][25] ), .S(
        \SUMB[2][25] ) );
  FA_X1 S2_2_26 ( .A(\ab[2][26] ), .B(n5), .CI(n36), .CO(\CARRYB[2][26] ), .S(
        \SUMB[2][26] ) );
  FA_X1 S2_2_27 ( .A(\ab[2][27] ), .B(n4), .CI(n35), .CO(\CARRYB[2][27] ), .S(
        \SUMB[2][27] ) );
  FA_X1 S2_2_28 ( .A(\ab[2][28] ), .B(n3), .CI(n34), .CO(\CARRYB[2][28] ), .S(
        \SUMB[2][28] ) );
  FA_X1 S2_2_29 ( .A(\ab[2][29] ), .B(n2), .CI(n33), .CO(\CARRYB[2][29] ), .S(
        \SUMB[2][29] ) );
  FA_X1 S3_2_30 ( .A(\ab[2][30] ), .B(n32), .CI(\ab[1][31] ), .CO(
        \CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  VerilogMultiplier_DW01_add_0 FS_1 ( .A({n316, n112, n120, n110, n119, n109, 
        n118, n111, n117, n74, n101, n66, n100, n73, n99, n69, n98, n68, n67, 
        n102, n79, n72, n78, n70, n65, n77, n71, n97, n76, n75, n64, n80, 
        \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , 
        \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , 
        \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , 
        \A1[0] }), .B({n125, n116, n124, n115, n123, n114, n122, n113, n121, 
        n87, n107, n86, n106, n85, n105, n95, n104, n94, n93, n108, n92, n84, 
        n91, n96, n83, n90, n82, n103, n89, n88, n81, \A2[30] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[63:2]) );
  AND2_X1 U2 ( .A1(\ab[0][30] ), .A2(\ab[1][29] ), .ZN(n2) );
  AND2_X1 U3 ( .A1(\ab[0][29] ), .A2(\ab[1][28] ), .ZN(n3) );
  AND2_X1 U4 ( .A1(\ab[0][28] ), .A2(\ab[1][27] ), .ZN(n4) );
  AND2_X1 U5 ( .A1(\ab[0][27] ), .A2(\ab[1][26] ), .ZN(n5) );
  AND2_X1 U6 ( .A1(\ab[0][26] ), .A2(\ab[1][25] ), .ZN(n6) );
  AND2_X1 U7 ( .A1(\ab[0][25] ), .A2(\ab[1][24] ), .ZN(n7) );
  AND2_X1 U8 ( .A1(\ab[0][24] ), .A2(\ab[1][23] ), .ZN(n8) );
  AND2_X1 U9 ( .A1(\ab[0][23] ), .A2(\ab[1][22] ), .ZN(n9) );
  AND2_X1 U10 ( .A1(\ab[0][22] ), .A2(\ab[1][21] ), .ZN(n10) );
  AND2_X1 U11 ( .A1(\ab[0][21] ), .A2(\ab[1][20] ), .ZN(n11) );
  AND2_X1 U12 ( .A1(\ab[0][20] ), .A2(\ab[1][19] ), .ZN(n12) );
  AND2_X1 U13 ( .A1(\ab[0][19] ), .A2(\ab[1][18] ), .ZN(n13) );
  AND2_X1 U14 ( .A1(\ab[0][18] ), .A2(\ab[1][17] ), .ZN(n14) );
  AND2_X1 U15 ( .A1(\ab[0][17] ), .A2(\ab[1][16] ), .ZN(n15) );
  AND2_X1 U16 ( .A1(\ab[0][16] ), .A2(\ab[1][15] ), .ZN(n16) );
  AND2_X1 U17 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n17) );
  AND2_X1 U18 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n18) );
  AND2_X1 U19 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n19) );
  AND2_X1 U20 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n20) );
  AND2_X1 U21 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n21) );
  AND2_X1 U22 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n22) );
  AND2_X1 U23 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n23) );
  AND2_X1 U24 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n24) );
  AND2_X1 U25 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n25) );
  AND2_X1 U26 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n26) );
  AND2_X1 U27 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n27) );
  AND2_X1 U28 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n28) );
  AND2_X1 U29 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n29) );
  AND2_X1 U30 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n30) );
  AND2_X1 U31 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n31) );
  AND2_X1 U32 ( .A1(\ab[0][31] ), .A2(\ab[1][30] ), .ZN(n32) );
  XOR2_X1 U33 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Z(n33) );
  XOR2_X1 U34 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(n34) );
  XOR2_X1 U35 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(n35) );
  XOR2_X1 U36 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(n36) );
  XOR2_X1 U37 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(n37) );
  XOR2_X1 U38 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(n38) );
  XOR2_X1 U39 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(n39) );
  XOR2_X1 U40 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(n40) );
  XOR2_X1 U41 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(n41) );
  XOR2_X1 U42 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(n42) );
  XOR2_X1 U43 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(n43) );
  XOR2_X1 U44 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(n44) );
  XOR2_X1 U45 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(n45) );
  XOR2_X1 U46 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(n46) );
  XOR2_X1 U47 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(n47) );
  XOR2_X1 U48 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(n48) );
  XOR2_X1 U49 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n49) );
  XOR2_X1 U50 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n50) );
  XOR2_X1 U51 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n51) );
  XOR2_X1 U52 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n52) );
  XOR2_X1 U53 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n53) );
  XOR2_X1 U54 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n54) );
  XOR2_X1 U55 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n55) );
  XOR2_X1 U56 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n56) );
  XOR2_X1 U57 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n57) );
  XOR2_X1 U58 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n58) );
  XOR2_X1 U59 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n59) );
  XOR2_X1 U60 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n60) );
  XOR2_X1 U61 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n61) );
  XOR2_X1 U62 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n62) );
  XOR2_X1 U63 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  INV_X1 U64 ( .A(\CARRYB[31][31] ), .ZN(n316) );
  BUF_X1 U65 ( .A(n378), .Z(n307) );
  BUF_X1 U66 ( .A(n379), .Z(n310) );
  BUF_X1 U67 ( .A(n377), .Z(n304) );
  BUF_X1 U68 ( .A(n376), .Z(n301) );
  BUF_X1 U69 ( .A(n375), .Z(n298) );
  BUF_X1 U70 ( .A(n374), .Z(n295) );
  BUF_X1 U71 ( .A(n373), .Z(n292) );
  BUF_X1 U72 ( .A(n372), .Z(n289) );
  BUF_X1 U73 ( .A(n371), .Z(n286) );
  BUF_X1 U74 ( .A(n370), .Z(n283) );
  BUF_X1 U75 ( .A(n369), .Z(n280) );
  BUF_X1 U76 ( .A(n368), .Z(n277) );
  BUF_X1 U77 ( .A(n367), .Z(n274) );
  BUF_X1 U78 ( .A(n366), .Z(n271) );
  BUF_X1 U79 ( .A(n365), .Z(n268) );
  BUF_X1 U80 ( .A(n364), .Z(n265) );
  BUF_X1 U81 ( .A(n363), .Z(n262) );
  BUF_X1 U82 ( .A(n362), .Z(n259) );
  BUF_X1 U83 ( .A(n361), .Z(n256) );
  BUF_X1 U84 ( .A(n360), .Z(n253) );
  BUF_X1 U85 ( .A(n359), .Z(n250) );
  BUF_X1 U86 ( .A(n358), .Z(n247) );
  BUF_X1 U87 ( .A(n357), .Z(n244) );
  BUF_X1 U88 ( .A(n356), .Z(n241) );
  BUF_X1 U89 ( .A(n355), .Z(n238) );
  BUF_X1 U90 ( .A(n354), .Z(n235) );
  BUF_X1 U91 ( .A(n353), .Z(n232) );
  BUF_X1 U92 ( .A(n352), .Z(n229) );
  BUF_X1 U93 ( .A(n351), .Z(n226) );
  BUF_X1 U94 ( .A(n350), .Z(n223) );
  BUF_X1 U95 ( .A(n339), .Z(n192) );
  BUF_X1 U96 ( .A(n378), .Z(n308) );
  BUF_X1 U97 ( .A(n379), .Z(n311) );
  BUF_X1 U98 ( .A(n377), .Z(n305) );
  BUF_X1 U99 ( .A(n376), .Z(n302) );
  BUF_X1 U100 ( .A(n375), .Z(n299) );
  BUF_X1 U101 ( .A(n372), .Z(n290) );
  BUF_X1 U102 ( .A(n373), .Z(n293) );
  BUF_X1 U103 ( .A(n374), .Z(n296) );
  BUF_X1 U104 ( .A(n371), .Z(n287) );
  BUF_X1 U105 ( .A(n369), .Z(n281) );
  BUF_X1 U106 ( .A(n370), .Z(n284) );
  BUF_X1 U107 ( .A(n366), .Z(n272) );
  BUF_X1 U108 ( .A(n365), .Z(n269) );
  BUF_X1 U109 ( .A(n364), .Z(n266) );
  BUF_X1 U110 ( .A(n361), .Z(n257) );
  BUF_X1 U111 ( .A(n363), .Z(n263) );
  BUF_X1 U112 ( .A(n362), .Z(n260) );
  BUF_X1 U113 ( .A(n359), .Z(n251) );
  BUF_X1 U114 ( .A(n360), .Z(n254) );
  BUF_X1 U115 ( .A(n357), .Z(n245) );
  BUF_X1 U116 ( .A(n358), .Z(n248) );
  BUF_X1 U117 ( .A(n355), .Z(n239) );
  BUF_X1 U118 ( .A(n356), .Z(n242) );
  BUF_X1 U119 ( .A(n353), .Z(n233) );
  BUF_X1 U120 ( .A(n354), .Z(n236) );
  BUF_X1 U121 ( .A(n351), .Z(n227) );
  BUF_X1 U122 ( .A(n352), .Z(n230) );
  BUF_X1 U123 ( .A(n368), .Z(n278) );
  BUF_X1 U124 ( .A(n367), .Z(n275) );
  BUF_X1 U125 ( .A(n350), .Z(n224) );
  BUF_X1 U126 ( .A(n380), .Z(n313) );
  BUF_X1 U127 ( .A(n380), .Z(n314) );
  BUF_X1 U128 ( .A(n348), .Z(n218) );
  BUF_X1 U129 ( .A(n347), .Z(n215) );
  BUF_X1 U130 ( .A(n348), .Z(n219) );
  BUF_X1 U131 ( .A(n347), .Z(n216) );
  BUF_X1 U132 ( .A(n346), .Z(n213) );
  BUF_X1 U133 ( .A(n345), .Z(n209) );
  BUF_X1 U134 ( .A(n345), .Z(n210) );
  BUF_X1 U135 ( .A(n344), .Z(n206) );
  BUF_X1 U136 ( .A(n344), .Z(n207) );
  BUF_X1 U137 ( .A(n343), .Z(n203) );
  BUF_X1 U138 ( .A(n343), .Z(n204) );
  BUF_X1 U139 ( .A(n342), .Z(n200) );
  BUF_X1 U140 ( .A(n342), .Z(n201) );
  BUF_X1 U141 ( .A(n341), .Z(n197) );
  BUF_X1 U142 ( .A(n341), .Z(n198) );
  BUF_X1 U143 ( .A(n340), .Z(n194) );
  BUF_X1 U144 ( .A(n340), .Z(n195) );
  BUF_X1 U145 ( .A(n346), .Z(n212) );
  BUF_X1 U146 ( .A(n349), .Z(n221) );
  BUF_X1 U147 ( .A(n379), .Z(n312) );
  BUF_X1 U148 ( .A(n377), .Z(n306) );
  BUF_X1 U149 ( .A(n376), .Z(n303) );
  BUF_X1 U150 ( .A(n375), .Z(n300) );
  BUF_X1 U151 ( .A(n351), .Z(n228) );
  BUF_X1 U152 ( .A(n374), .Z(n297) );
  BUF_X1 U153 ( .A(n373), .Z(n294) );
  BUF_X1 U154 ( .A(n372), .Z(n291) );
  BUF_X1 U155 ( .A(n371), .Z(n288) );
  BUF_X1 U156 ( .A(n370), .Z(n285) );
  BUF_X1 U157 ( .A(n369), .Z(n282) );
  BUF_X1 U158 ( .A(n368), .Z(n279) );
  BUF_X1 U159 ( .A(n367), .Z(n276) );
  BUF_X1 U160 ( .A(n366), .Z(n273) );
  BUF_X1 U161 ( .A(n365), .Z(n270) );
  BUF_X1 U162 ( .A(n364), .Z(n267) );
  BUF_X1 U163 ( .A(n363), .Z(n264) );
  BUF_X1 U164 ( .A(n362), .Z(n261) );
  BUF_X1 U165 ( .A(n361), .Z(n258) );
  BUF_X1 U166 ( .A(n360), .Z(n255) );
  BUF_X1 U167 ( .A(n359), .Z(n252) );
  BUF_X1 U168 ( .A(n358), .Z(n249) );
  BUF_X1 U169 ( .A(n357), .Z(n246) );
  BUF_X1 U170 ( .A(n356), .Z(n243) );
  BUF_X1 U171 ( .A(n355), .Z(n240) );
  BUF_X1 U172 ( .A(n354), .Z(n237) );
  BUF_X1 U173 ( .A(n378), .Z(n309) );
  BUF_X1 U174 ( .A(n352), .Z(n231) );
  BUF_X1 U175 ( .A(n353), .Z(n234) );
  BUF_X1 U176 ( .A(n350), .Z(n225) );
  BUF_X1 U177 ( .A(n380), .Z(n315) );
  BUF_X1 U178 ( .A(n348), .Z(n220) );
  BUF_X1 U179 ( .A(n347), .Z(n217) );
  BUF_X1 U180 ( .A(n346), .Z(n214) );
  BUF_X1 U181 ( .A(n345), .Z(n211) );
  BUF_X1 U182 ( .A(n344), .Z(n208) );
  BUF_X1 U183 ( .A(n343), .Z(n205) );
  BUF_X1 U184 ( .A(n342), .Z(n202) );
  BUF_X1 U185 ( .A(n341), .Z(n199) );
  BUF_X1 U186 ( .A(n349), .Z(n222) );
  XOR2_X1 U187 ( .A(\CARRYB[31][1] ), .B(\SUMB[31][2] ), .Z(n64) );
  XOR2_X1 U188 ( .A(\CARRYB[31][7] ), .B(\SUMB[31][8] ), .Z(n65) );
  XOR2_X1 U189 ( .A(\CARRYB[31][20] ), .B(\SUMB[31][21] ), .Z(n66) );
  XOR2_X1 U190 ( .A(\CARRYB[31][13] ), .B(\SUMB[31][14] ), .Z(n67) );
  XOR2_X1 U191 ( .A(\CARRYB[31][14] ), .B(\SUMB[31][15] ), .Z(n68) );
  XOR2_X1 U192 ( .A(\CARRYB[31][16] ), .B(\SUMB[31][17] ), .Z(n69) );
  XOR2_X1 U193 ( .A(\CARRYB[31][8] ), .B(\SUMB[31][9] ), .Z(n70) );
  XOR2_X1 U194 ( .A(\CARRYB[31][5] ), .B(\SUMB[31][6] ), .Z(n71) );
  XOR2_X1 U195 ( .A(\CARRYB[31][10] ), .B(\SUMB[31][11] ), .Z(n72) );
  XOR2_X1 U196 ( .A(\CARRYB[31][18] ), .B(\SUMB[31][19] ), .Z(n73) );
  XOR2_X1 U197 ( .A(\CARRYB[31][22] ), .B(\SUMB[31][23] ), .Z(n74) );
  XOR2_X1 U198 ( .A(\CARRYB[31][2] ), .B(\SUMB[31][3] ), .Z(n75) );
  XOR2_X1 U199 ( .A(\CARRYB[31][3] ), .B(\SUMB[31][4] ), .Z(n76) );
  XOR2_X1 U200 ( .A(\CARRYB[31][6] ), .B(\SUMB[31][7] ), .Z(n77) );
  XOR2_X1 U201 ( .A(\CARRYB[31][9] ), .B(\SUMB[31][10] ), .Z(n78) );
  XOR2_X1 U202 ( .A(\CARRYB[31][11] ), .B(\SUMB[31][12] ), .Z(n79) );
  XOR2_X1 U203 ( .A(\CARRYB[31][0] ), .B(\SUMB[31][1] ), .Z(n80) );
  AND2_X1 U204 ( .A1(\CARRYB[31][0] ), .A2(\SUMB[31][1] ), .ZN(n81) );
  AND2_X1 U205 ( .A1(\CARRYB[31][4] ), .A2(\SUMB[31][5] ), .ZN(n82) );
  AND2_X1 U206 ( .A1(\CARRYB[31][6] ), .A2(\SUMB[31][7] ), .ZN(n83) );
  AND2_X1 U207 ( .A1(\CARRYB[31][9] ), .A2(\SUMB[31][10] ), .ZN(n84) );
  AND2_X1 U208 ( .A1(\CARRYB[31][17] ), .A2(\SUMB[31][18] ), .ZN(n85) );
  AND2_X1 U209 ( .A1(\CARRYB[31][19] ), .A2(\SUMB[31][20] ), .ZN(n86) );
  AND2_X1 U210 ( .A1(\CARRYB[31][21] ), .A2(\SUMB[31][22] ), .ZN(n87) );
  AND2_X1 U211 ( .A1(\CARRYB[31][1] ), .A2(\SUMB[31][2] ), .ZN(n88) );
  AND2_X1 U212 ( .A1(\CARRYB[31][2] ), .A2(\SUMB[31][3] ), .ZN(n89) );
  AND2_X1 U213 ( .A1(\CARRYB[31][5] ), .A2(\SUMB[31][6] ), .ZN(n90) );
  AND2_X1 U214 ( .A1(\CARRYB[31][8] ), .A2(\SUMB[31][9] ), .ZN(n91) );
  AND2_X1 U215 ( .A1(\CARRYB[31][10] ), .A2(\SUMB[31][11] ), .ZN(n92) );
  AND2_X1 U216 ( .A1(\CARRYB[31][12] ), .A2(\SUMB[31][13] ), .ZN(n93) );
  AND2_X1 U217 ( .A1(\CARRYB[31][13] ), .A2(\SUMB[31][14] ), .ZN(n94) );
  AND2_X1 U218 ( .A1(\CARRYB[31][15] ), .A2(\SUMB[31][16] ), .ZN(n95) );
  AND2_X1 U219 ( .A1(\CARRYB[31][7] ), .A2(\SUMB[31][8] ), .ZN(n96) );
  XOR2_X1 U220 ( .A(\CARRYB[31][4] ), .B(\SUMB[31][5] ), .Z(n97) );
  XOR2_X1 U221 ( .A(\CARRYB[31][15] ), .B(\SUMB[31][16] ), .Z(n98) );
  XOR2_X1 U222 ( .A(\CARRYB[31][17] ), .B(\SUMB[31][18] ), .Z(n99) );
  XOR2_X1 U223 ( .A(\CARRYB[31][19] ), .B(\SUMB[31][20] ), .Z(n100) );
  XOR2_X1 U224 ( .A(\CARRYB[31][21] ), .B(\SUMB[31][22] ), .Z(n101) );
  XOR2_X1 U225 ( .A(\CARRYB[31][12] ), .B(\SUMB[31][13] ), .Z(n102) );
  AND2_X1 U226 ( .A1(\CARRYB[31][3] ), .A2(\SUMB[31][4] ), .ZN(n103) );
  AND2_X1 U227 ( .A1(\CARRYB[31][14] ), .A2(\SUMB[31][15] ), .ZN(n104) );
  AND2_X1 U228 ( .A1(\CARRYB[31][16] ), .A2(\SUMB[31][17] ), .ZN(n105) );
  AND2_X1 U229 ( .A1(\CARRYB[31][18] ), .A2(\SUMB[31][19] ), .ZN(n106) );
  AND2_X1 U230 ( .A1(\CARRYB[31][20] ), .A2(\SUMB[31][21] ), .ZN(n107) );
  AND2_X1 U231 ( .A1(\CARRYB[31][11] ), .A2(\SUMB[31][12] ), .ZN(n108) );
  BUF_X1 U232 ( .A(n339), .Z(n191) );
  BUF_X1 U233 ( .A(n338), .Z(n188) );
  BUF_X1 U234 ( .A(n337), .Z(n185) );
  BUF_X1 U235 ( .A(n336), .Z(n182) );
  BUF_X1 U236 ( .A(n338), .Z(n189) );
  BUF_X1 U237 ( .A(n335), .Z(n179) );
  BUF_X1 U238 ( .A(n337), .Z(n186) );
  BUF_X1 U239 ( .A(n334), .Z(n176) );
  BUF_X1 U240 ( .A(n333), .Z(n173) );
  BUF_X1 U241 ( .A(n332), .Z(n170) );
  BUF_X1 U242 ( .A(n331), .Z(n167) );
  BUF_X1 U243 ( .A(n330), .Z(n164) );
  BUF_X1 U244 ( .A(n336), .Z(n183) );
  BUF_X1 U245 ( .A(n335), .Z(n180) );
  BUF_X1 U246 ( .A(n334), .Z(n177) );
  BUF_X1 U247 ( .A(n333), .Z(n174) );
  BUF_X1 U248 ( .A(n332), .Z(n171) );
  BUF_X1 U249 ( .A(n331), .Z(n168) );
  BUF_X1 U250 ( .A(n330), .Z(n165) );
  BUF_X1 U251 ( .A(n339), .Z(n193) );
  BUF_X1 U252 ( .A(n340), .Z(n196) );
  BUF_X1 U253 ( .A(n338), .Z(n190) );
  BUF_X1 U254 ( .A(n337), .Z(n187) );
  BUF_X1 U255 ( .A(n336), .Z(n184) );
  BUF_X1 U256 ( .A(n335), .Z(n181) );
  BUF_X1 U257 ( .A(n334), .Z(n178) );
  BUF_X1 U258 ( .A(n333), .Z(n175) );
  BUF_X1 U259 ( .A(n332), .Z(n172) );
  BUF_X1 U260 ( .A(n331), .Z(n169) );
  XOR2_X1 U261 ( .A(\CARRYB[31][26] ), .B(\SUMB[31][27] ), .Z(n109) );
  XOR2_X1 U262 ( .A(\CARRYB[31][28] ), .B(\SUMB[31][29] ), .Z(n110) );
  XOR2_X1 U263 ( .A(\CARRYB[31][24] ), .B(\SUMB[31][25] ), .Z(n111) );
  XOR2_X1 U264 ( .A(\CARRYB[31][30] ), .B(\SUMB[31][31] ), .Z(n112) );
  AND2_X1 U265 ( .A1(\CARRYB[31][23] ), .A2(\SUMB[31][24] ), .ZN(n113) );
  AND2_X1 U266 ( .A1(\CARRYB[31][25] ), .A2(\SUMB[31][26] ), .ZN(n114) );
  AND2_X1 U267 ( .A1(\CARRYB[31][27] ), .A2(\SUMB[31][28] ), .ZN(n115) );
  AND2_X1 U268 ( .A1(\CARRYB[31][29] ), .A2(\SUMB[31][30] ), .ZN(n116) );
  XOR2_X1 U269 ( .A(\CARRYB[31][23] ), .B(\SUMB[31][24] ), .Z(n117) );
  XOR2_X1 U270 ( .A(\CARRYB[31][25] ), .B(\SUMB[31][26] ), .Z(n118) );
  XOR2_X1 U271 ( .A(\CARRYB[31][27] ), .B(\SUMB[31][28] ), .Z(n119) );
  XOR2_X1 U272 ( .A(\CARRYB[31][29] ), .B(\SUMB[31][30] ), .Z(n120) );
  AND2_X1 U273 ( .A1(\CARRYB[31][22] ), .A2(\SUMB[31][23] ), .ZN(n121) );
  AND2_X1 U274 ( .A1(\CARRYB[31][24] ), .A2(\SUMB[31][25] ), .ZN(n122) );
  AND2_X1 U275 ( .A1(\CARRYB[31][26] ), .A2(\SUMB[31][27] ), .ZN(n123) );
  AND2_X1 U276 ( .A1(\CARRYB[31][28] ), .A2(\SUMB[31][29] ), .ZN(n124) );
  AND2_X1 U277 ( .A1(\CARRYB[31][30] ), .A2(\SUMB[31][31] ), .ZN(n125) );
  BUF_X1 U278 ( .A(n329), .Z(n161) );
  BUF_X1 U279 ( .A(n328), .Z(n158) );
  BUF_X1 U280 ( .A(n327), .Z(n155) );
  BUF_X1 U281 ( .A(n326), .Z(n152) );
  BUF_X1 U282 ( .A(n325), .Z(n149) );
  BUF_X1 U283 ( .A(n324), .Z(n146) );
  BUF_X1 U284 ( .A(n323), .Z(n143) );
  BUF_X1 U285 ( .A(n322), .Z(n140) );
  BUF_X1 U286 ( .A(n321), .Z(n137) );
  BUF_X1 U287 ( .A(n329), .Z(n162) );
  BUF_X1 U288 ( .A(n328), .Z(n159) );
  BUF_X1 U289 ( .A(n327), .Z(n156) );
  BUF_X1 U290 ( .A(n326), .Z(n153) );
  BUF_X1 U291 ( .A(n325), .Z(n150) );
  BUF_X1 U292 ( .A(n324), .Z(n147) );
  BUF_X1 U293 ( .A(n323), .Z(n144) );
  BUF_X1 U294 ( .A(n322), .Z(n141) );
  BUF_X1 U295 ( .A(n330), .Z(n166) );
  BUF_X1 U296 ( .A(n329), .Z(n163) );
  BUF_X1 U297 ( .A(n328), .Z(n160) );
  BUF_X1 U298 ( .A(n327), .Z(n157) );
  BUF_X1 U299 ( .A(n326), .Z(n154) );
  BUF_X1 U300 ( .A(n325), .Z(n151) );
  BUF_X1 U301 ( .A(n324), .Z(n148) );
  BUF_X1 U302 ( .A(n323), .Z(n145) );
  BUF_X1 U303 ( .A(n322), .Z(n142) );
  BUF_X1 U304 ( .A(n321), .Z(n139) );
  BUF_X1 U305 ( .A(n320), .Z(n134) );
  BUF_X1 U306 ( .A(n319), .Z(n131) );
  BUF_X1 U307 ( .A(n318), .Z(n128) );
  BUF_X1 U308 ( .A(n317), .Z(n127) );
  BUF_X1 U309 ( .A(n321), .Z(n138) );
  BUF_X1 U310 ( .A(n320), .Z(n135) );
  BUF_X1 U311 ( .A(n319), .Z(n132) );
  BUF_X1 U312 ( .A(n318), .Z(n129) );
  BUF_X1 U313 ( .A(n317), .Z(n126) );
  BUF_X1 U314 ( .A(n320), .Z(n136) );
  BUF_X1 U315 ( .A(n319), .Z(n133) );
  BUF_X1 U316 ( .A(n318), .Z(n130) );
  INV_X1 U317 ( .A(ZB), .ZN(n349) );
  INV_X1 U318 ( .A(B[2]), .ZN(n378) );
  INV_X1 U319 ( .A(B[1]), .ZN(n379) );
  INV_X1 U320 ( .A(B[3]), .ZN(n377) );
  INV_X1 U321 ( .A(B[4]), .ZN(n376) );
  INV_X1 U322 ( .A(B[5]), .ZN(n375) );
  INV_X1 U323 ( .A(B[6]), .ZN(n374) );
  INV_X1 U324 ( .A(B[7]), .ZN(n373) );
  INV_X1 U325 ( .A(B[8]), .ZN(n372) );
  INV_X1 U326 ( .A(B[9]), .ZN(n371) );
  INV_X1 U327 ( .A(B[10]), .ZN(n370) );
  INV_X1 U328 ( .A(B[11]), .ZN(n369) );
  INV_X1 U329 ( .A(B[12]), .ZN(n368) );
  INV_X1 U330 ( .A(B[13]), .ZN(n367) );
  INV_X1 U331 ( .A(B[14]), .ZN(n366) );
  INV_X1 U332 ( .A(B[15]), .ZN(n365) );
  INV_X1 U333 ( .A(B[16]), .ZN(n364) );
  INV_X1 U334 ( .A(B[17]), .ZN(n363) );
  INV_X1 U335 ( .A(B[18]), .ZN(n362) );
  INV_X1 U336 ( .A(B[19]), .ZN(n361) );
  INV_X1 U337 ( .A(B[20]), .ZN(n360) );
  INV_X1 U338 ( .A(B[21]), .ZN(n359) );
  INV_X1 U339 ( .A(B[22]), .ZN(n358) );
  INV_X1 U340 ( .A(B[23]), .ZN(n357) );
  INV_X1 U341 ( .A(B[24]), .ZN(n356) );
  INV_X1 U342 ( .A(B[25]), .ZN(n355) );
  INV_X1 U343 ( .A(B[26]), .ZN(n354) );
  INV_X1 U344 ( .A(B[27]), .ZN(n353) );
  INV_X1 U345 ( .A(B[28]), .ZN(n352) );
  INV_X1 U346 ( .A(A[0]), .ZN(n348) );
  INV_X1 U347 ( .A(B[29]), .ZN(n351) );
  INV_X1 U348 ( .A(B[30]), .ZN(n350) );
  INV_X1 U349 ( .A(A[1]), .ZN(n347) );
  INV_X1 U350 ( .A(A[2]), .ZN(n346) );
  INV_X1 U351 ( .A(A[3]), .ZN(n345) );
  INV_X1 U352 ( .A(A[4]), .ZN(n344) );
  INV_X1 U353 ( .A(A[5]), .ZN(n343) );
  INV_X1 U354 ( .A(A[6]), .ZN(n342) );
  INV_X1 U355 ( .A(A[7]), .ZN(n341) );
  INV_X1 U356 ( .A(A[8]), .ZN(n340) );
  INV_X1 U357 ( .A(A[9]), .ZN(n339) );
  INV_X1 U358 ( .A(B[0]), .ZN(n380) );
  INV_X1 U359 ( .A(A[10]), .ZN(n338) );
  INV_X1 U360 ( .A(A[11]), .ZN(n337) );
  INV_X1 U361 ( .A(A[12]), .ZN(n336) );
  INV_X1 U362 ( .A(A[13]), .ZN(n335) );
  INV_X1 U363 ( .A(A[14]), .ZN(n334) );
  INV_X1 U364 ( .A(A[15]), .ZN(n333) );
  INV_X1 U365 ( .A(A[16]), .ZN(n332) );
  INV_X1 U366 ( .A(A[17]), .ZN(n331) );
  INV_X1 U367 ( .A(A[18]), .ZN(n330) );
  INV_X1 U368 ( .A(A[19]), .ZN(n329) );
  INV_X1 U369 ( .A(A[20]), .ZN(n328) );
  INV_X1 U370 ( .A(A[21]), .ZN(n327) );
  INV_X1 U371 ( .A(A[22]), .ZN(n326) );
  INV_X1 U372 ( .A(A[23]), .ZN(n325) );
  INV_X1 U373 ( .A(A[24]), .ZN(n324) );
  INV_X1 U374 ( .A(A[25]), .ZN(n323) );
  INV_X1 U375 ( .A(A[26]), .ZN(n322) );
  INV_X1 U376 ( .A(A[27]), .ZN(n321) );
  INV_X1 U377 ( .A(A[28]), .ZN(n320) );
  INV_X1 U378 ( .A(A[29]), .ZN(n319) );
  INV_X1 U379 ( .A(A[30]), .ZN(n318) );
  INV_X1 U380 ( .A(ZA), .ZN(n317) );
  NOR2_X1 U381 ( .A1(n193), .A2(n288), .ZN(\ab[9][9] ) );
  NOR2_X1 U382 ( .A1(n193), .A2(n291), .ZN(\ab[9][8] ) );
  NOR2_X1 U383 ( .A1(n193), .A2(n294), .ZN(\ab[9][7] ) );
  NOR2_X1 U384 ( .A1(n193), .A2(n297), .ZN(\ab[9][6] ) );
  NOR2_X1 U385 ( .A1(n193), .A2(n300), .ZN(\ab[9][5] ) );
  NOR2_X1 U386 ( .A1(n193), .A2(n303), .ZN(\ab[9][4] ) );
  NOR2_X1 U387 ( .A1(n193), .A2(n306), .ZN(\ab[9][3] ) );
  NOR2_X1 U388 ( .A1(A[9]), .A2(n221), .ZN(\ab[9][31] ) );
  NOR2_X1 U389 ( .A1(n192), .A2(n225), .ZN(\ab[9][30] ) );
  NOR2_X1 U390 ( .A1(n192), .A2(n309), .ZN(\ab[9][2] ) );
  NOR2_X1 U391 ( .A1(n192), .A2(n228), .ZN(\ab[9][29] ) );
  NOR2_X1 U392 ( .A1(n192), .A2(n231), .ZN(\ab[9][28] ) );
  NOR2_X1 U393 ( .A1(n192), .A2(n234), .ZN(\ab[9][27] ) );
  NOR2_X1 U394 ( .A1(n192), .A2(n237), .ZN(\ab[9][26] ) );
  NOR2_X1 U395 ( .A1(n192), .A2(n240), .ZN(\ab[9][25] ) );
  NOR2_X1 U396 ( .A1(n192), .A2(n243), .ZN(\ab[9][24] ) );
  NOR2_X1 U397 ( .A1(n192), .A2(n246), .ZN(\ab[9][23] ) );
  NOR2_X1 U398 ( .A1(n192), .A2(n249), .ZN(\ab[9][22] ) );
  NOR2_X1 U399 ( .A1(n192), .A2(n252), .ZN(\ab[9][21] ) );
  NOR2_X1 U400 ( .A1(n192), .A2(n255), .ZN(\ab[9][20] ) );
  NOR2_X1 U401 ( .A1(n191), .A2(n312), .ZN(\ab[9][1] ) );
  NOR2_X1 U402 ( .A1(n191), .A2(n258), .ZN(\ab[9][19] ) );
  NOR2_X1 U403 ( .A1(n191), .A2(n261), .ZN(\ab[9][18] ) );
  NOR2_X1 U404 ( .A1(n191), .A2(n264), .ZN(\ab[9][17] ) );
  NOR2_X1 U405 ( .A1(n191), .A2(n267), .ZN(\ab[9][16] ) );
  NOR2_X1 U406 ( .A1(n191), .A2(n270), .ZN(\ab[9][15] ) );
  NOR2_X1 U407 ( .A1(n191), .A2(n273), .ZN(\ab[9][14] ) );
  NOR2_X1 U408 ( .A1(n191), .A2(n276), .ZN(\ab[9][13] ) );
  NOR2_X1 U409 ( .A1(n191), .A2(n279), .ZN(\ab[9][12] ) );
  NOR2_X1 U410 ( .A1(n191), .A2(n282), .ZN(\ab[9][11] ) );
  NOR2_X1 U411 ( .A1(n191), .A2(n285), .ZN(\ab[9][10] ) );
  NOR2_X1 U412 ( .A1(n191), .A2(n315), .ZN(\ab[9][0] ) );
  NOR2_X1 U413 ( .A1(n288), .A2(n196), .ZN(\ab[8][9] ) );
  NOR2_X1 U414 ( .A1(n291), .A2(n196), .ZN(\ab[8][8] ) );
  NOR2_X1 U415 ( .A1(n294), .A2(n196), .ZN(\ab[8][7] ) );
  NOR2_X1 U416 ( .A1(n297), .A2(n196), .ZN(\ab[8][6] ) );
  NOR2_X1 U417 ( .A1(n300), .A2(n196), .ZN(\ab[8][5] ) );
  NOR2_X1 U418 ( .A1(n303), .A2(n196), .ZN(\ab[8][4] ) );
  NOR2_X1 U419 ( .A1(n306), .A2(n196), .ZN(\ab[8][3] ) );
  NOR2_X1 U420 ( .A1(A[8]), .A2(n222), .ZN(\ab[8][31] ) );
  NOR2_X1 U421 ( .A1(n225), .A2(n195), .ZN(\ab[8][30] ) );
  NOR2_X1 U422 ( .A1(n309), .A2(n195), .ZN(\ab[8][2] ) );
  NOR2_X1 U423 ( .A1(n228), .A2(n195), .ZN(\ab[8][29] ) );
  NOR2_X1 U424 ( .A1(n231), .A2(n195), .ZN(\ab[8][28] ) );
  NOR2_X1 U425 ( .A1(n234), .A2(n195), .ZN(\ab[8][27] ) );
  NOR2_X1 U426 ( .A1(n237), .A2(n195), .ZN(\ab[8][26] ) );
  NOR2_X1 U427 ( .A1(n240), .A2(n195), .ZN(\ab[8][25] ) );
  NOR2_X1 U428 ( .A1(n243), .A2(n195), .ZN(\ab[8][24] ) );
  NOR2_X1 U429 ( .A1(n246), .A2(n195), .ZN(\ab[8][23] ) );
  NOR2_X1 U430 ( .A1(n249), .A2(n195), .ZN(\ab[8][22] ) );
  NOR2_X1 U431 ( .A1(n252), .A2(n195), .ZN(\ab[8][21] ) );
  NOR2_X1 U432 ( .A1(n255), .A2(n195), .ZN(\ab[8][20] ) );
  NOR2_X1 U433 ( .A1(n312), .A2(n194), .ZN(\ab[8][1] ) );
  NOR2_X1 U434 ( .A1(n258), .A2(n194), .ZN(\ab[8][19] ) );
  NOR2_X1 U435 ( .A1(n261), .A2(n194), .ZN(\ab[8][18] ) );
  NOR2_X1 U436 ( .A1(n264), .A2(n194), .ZN(\ab[8][17] ) );
  NOR2_X1 U437 ( .A1(n267), .A2(n194), .ZN(\ab[8][16] ) );
  NOR2_X1 U438 ( .A1(n270), .A2(n194), .ZN(\ab[8][15] ) );
  NOR2_X1 U439 ( .A1(n273), .A2(n194), .ZN(\ab[8][14] ) );
  NOR2_X1 U440 ( .A1(n276), .A2(n194), .ZN(\ab[8][13] ) );
  NOR2_X1 U441 ( .A1(n279), .A2(n194), .ZN(\ab[8][12] ) );
  NOR2_X1 U442 ( .A1(n282), .A2(n194), .ZN(\ab[8][11] ) );
  NOR2_X1 U443 ( .A1(n285), .A2(n194), .ZN(\ab[8][10] ) );
  NOR2_X1 U444 ( .A1(n315), .A2(n194), .ZN(\ab[8][0] ) );
  NOR2_X1 U445 ( .A1(n288), .A2(n199), .ZN(\ab[7][9] ) );
  NOR2_X1 U446 ( .A1(n291), .A2(n199), .ZN(\ab[7][8] ) );
  NOR2_X1 U447 ( .A1(n294), .A2(n199), .ZN(\ab[7][7] ) );
  NOR2_X1 U448 ( .A1(n297), .A2(n199), .ZN(\ab[7][6] ) );
  NOR2_X1 U449 ( .A1(n300), .A2(n199), .ZN(\ab[7][5] ) );
  NOR2_X1 U450 ( .A1(n303), .A2(n199), .ZN(\ab[7][4] ) );
  NOR2_X1 U451 ( .A1(n306), .A2(n199), .ZN(\ab[7][3] ) );
  NOR2_X1 U452 ( .A1(A[7]), .A2(n222), .ZN(\ab[7][31] ) );
  NOR2_X1 U453 ( .A1(n225), .A2(n198), .ZN(\ab[7][30] ) );
  NOR2_X1 U454 ( .A1(n309), .A2(n198), .ZN(\ab[7][2] ) );
  NOR2_X1 U455 ( .A1(n228), .A2(n198), .ZN(\ab[7][29] ) );
  NOR2_X1 U456 ( .A1(n231), .A2(n198), .ZN(\ab[7][28] ) );
  NOR2_X1 U457 ( .A1(n234), .A2(n198), .ZN(\ab[7][27] ) );
  NOR2_X1 U458 ( .A1(n237), .A2(n198), .ZN(\ab[7][26] ) );
  NOR2_X1 U459 ( .A1(n240), .A2(n198), .ZN(\ab[7][25] ) );
  NOR2_X1 U460 ( .A1(n243), .A2(n198), .ZN(\ab[7][24] ) );
  NOR2_X1 U461 ( .A1(n246), .A2(n198), .ZN(\ab[7][23] ) );
  NOR2_X1 U462 ( .A1(n249), .A2(n198), .ZN(\ab[7][22] ) );
  NOR2_X1 U463 ( .A1(n252), .A2(n198), .ZN(\ab[7][21] ) );
  NOR2_X1 U464 ( .A1(n255), .A2(n198), .ZN(\ab[7][20] ) );
  NOR2_X1 U465 ( .A1(n312), .A2(n197), .ZN(\ab[7][1] ) );
  NOR2_X1 U466 ( .A1(n258), .A2(n197), .ZN(\ab[7][19] ) );
  NOR2_X1 U467 ( .A1(n261), .A2(n197), .ZN(\ab[7][18] ) );
  NOR2_X1 U468 ( .A1(n264), .A2(n197), .ZN(\ab[7][17] ) );
  NOR2_X1 U469 ( .A1(n267), .A2(n197), .ZN(\ab[7][16] ) );
  NOR2_X1 U470 ( .A1(n270), .A2(n197), .ZN(\ab[7][15] ) );
  NOR2_X1 U471 ( .A1(n273), .A2(n197), .ZN(\ab[7][14] ) );
  NOR2_X1 U472 ( .A1(n276), .A2(n197), .ZN(\ab[7][13] ) );
  NOR2_X1 U473 ( .A1(n279), .A2(n197), .ZN(\ab[7][12] ) );
  NOR2_X1 U474 ( .A1(n282), .A2(n197), .ZN(\ab[7][11] ) );
  NOR2_X1 U475 ( .A1(n285), .A2(n197), .ZN(\ab[7][10] ) );
  NOR2_X1 U476 ( .A1(n315), .A2(n197), .ZN(\ab[7][0] ) );
  NOR2_X1 U477 ( .A1(n288), .A2(n202), .ZN(\ab[6][9] ) );
  NOR2_X1 U478 ( .A1(n291), .A2(n202), .ZN(\ab[6][8] ) );
  NOR2_X1 U479 ( .A1(n294), .A2(n202), .ZN(\ab[6][7] ) );
  NOR2_X1 U480 ( .A1(n297), .A2(n202), .ZN(\ab[6][6] ) );
  NOR2_X1 U481 ( .A1(n300), .A2(n202), .ZN(\ab[6][5] ) );
  NOR2_X1 U482 ( .A1(n303), .A2(n202), .ZN(\ab[6][4] ) );
  NOR2_X1 U483 ( .A1(n306), .A2(n202), .ZN(\ab[6][3] ) );
  NOR2_X1 U484 ( .A1(A[6]), .A2(n222), .ZN(\ab[6][31] ) );
  NOR2_X1 U485 ( .A1(n225), .A2(n201), .ZN(\ab[6][30] ) );
  NOR2_X1 U486 ( .A1(n309), .A2(n201), .ZN(\ab[6][2] ) );
  NOR2_X1 U487 ( .A1(n228), .A2(n201), .ZN(\ab[6][29] ) );
  NOR2_X1 U488 ( .A1(n231), .A2(n201), .ZN(\ab[6][28] ) );
  NOR2_X1 U489 ( .A1(n234), .A2(n201), .ZN(\ab[6][27] ) );
  NOR2_X1 U490 ( .A1(n237), .A2(n201), .ZN(\ab[6][26] ) );
  NOR2_X1 U491 ( .A1(n240), .A2(n201), .ZN(\ab[6][25] ) );
  NOR2_X1 U492 ( .A1(n243), .A2(n201), .ZN(\ab[6][24] ) );
  NOR2_X1 U493 ( .A1(n246), .A2(n201), .ZN(\ab[6][23] ) );
  NOR2_X1 U494 ( .A1(n249), .A2(n201), .ZN(\ab[6][22] ) );
  NOR2_X1 U495 ( .A1(n252), .A2(n201), .ZN(\ab[6][21] ) );
  NOR2_X1 U496 ( .A1(n255), .A2(n201), .ZN(\ab[6][20] ) );
  NOR2_X1 U497 ( .A1(n312), .A2(n200), .ZN(\ab[6][1] ) );
  NOR2_X1 U498 ( .A1(n258), .A2(n200), .ZN(\ab[6][19] ) );
  NOR2_X1 U499 ( .A1(n261), .A2(n200), .ZN(\ab[6][18] ) );
  NOR2_X1 U500 ( .A1(n264), .A2(n200), .ZN(\ab[6][17] ) );
  NOR2_X1 U501 ( .A1(n267), .A2(n200), .ZN(\ab[6][16] ) );
  NOR2_X1 U502 ( .A1(n270), .A2(n200), .ZN(\ab[6][15] ) );
  NOR2_X1 U503 ( .A1(n273), .A2(n200), .ZN(\ab[6][14] ) );
  NOR2_X1 U504 ( .A1(n276), .A2(n200), .ZN(\ab[6][13] ) );
  NOR2_X1 U505 ( .A1(n279), .A2(n200), .ZN(\ab[6][12] ) );
  NOR2_X1 U506 ( .A1(n282), .A2(n200), .ZN(\ab[6][11] ) );
  NOR2_X1 U507 ( .A1(n285), .A2(n200), .ZN(\ab[6][10] ) );
  NOR2_X1 U508 ( .A1(n315), .A2(n200), .ZN(\ab[6][0] ) );
  NOR2_X1 U509 ( .A1(n288), .A2(n205), .ZN(\ab[5][9] ) );
  NOR2_X1 U510 ( .A1(n291), .A2(n205), .ZN(\ab[5][8] ) );
  NOR2_X1 U511 ( .A1(n294), .A2(n205), .ZN(\ab[5][7] ) );
  NOR2_X1 U512 ( .A1(n297), .A2(n205), .ZN(\ab[5][6] ) );
  NOR2_X1 U513 ( .A1(n300), .A2(n205), .ZN(\ab[5][5] ) );
  NOR2_X1 U514 ( .A1(n303), .A2(n205), .ZN(\ab[5][4] ) );
  NOR2_X1 U515 ( .A1(n306), .A2(n205), .ZN(\ab[5][3] ) );
  NOR2_X1 U516 ( .A1(A[5]), .A2(n222), .ZN(\ab[5][31] ) );
  NOR2_X1 U517 ( .A1(n225), .A2(n204), .ZN(\ab[5][30] ) );
  NOR2_X1 U518 ( .A1(n309), .A2(n204), .ZN(\ab[5][2] ) );
  NOR2_X1 U519 ( .A1(n228), .A2(n204), .ZN(\ab[5][29] ) );
  NOR2_X1 U520 ( .A1(n231), .A2(n204), .ZN(\ab[5][28] ) );
  NOR2_X1 U521 ( .A1(n234), .A2(n204), .ZN(\ab[5][27] ) );
  NOR2_X1 U522 ( .A1(n237), .A2(n204), .ZN(\ab[5][26] ) );
  NOR2_X1 U523 ( .A1(n240), .A2(n204), .ZN(\ab[5][25] ) );
  NOR2_X1 U524 ( .A1(n243), .A2(n204), .ZN(\ab[5][24] ) );
  NOR2_X1 U525 ( .A1(n246), .A2(n204), .ZN(\ab[5][23] ) );
  NOR2_X1 U526 ( .A1(n249), .A2(n204), .ZN(\ab[5][22] ) );
  NOR2_X1 U527 ( .A1(n252), .A2(n204), .ZN(\ab[5][21] ) );
  NOR2_X1 U528 ( .A1(n255), .A2(n204), .ZN(\ab[5][20] ) );
  NOR2_X1 U529 ( .A1(n312), .A2(n203), .ZN(\ab[5][1] ) );
  NOR2_X1 U530 ( .A1(n258), .A2(n203), .ZN(\ab[5][19] ) );
  NOR2_X1 U531 ( .A1(n261), .A2(n203), .ZN(\ab[5][18] ) );
  NOR2_X1 U532 ( .A1(n264), .A2(n203), .ZN(\ab[5][17] ) );
  NOR2_X1 U533 ( .A1(n267), .A2(n203), .ZN(\ab[5][16] ) );
  NOR2_X1 U534 ( .A1(n270), .A2(n203), .ZN(\ab[5][15] ) );
  NOR2_X1 U535 ( .A1(n273), .A2(n203), .ZN(\ab[5][14] ) );
  NOR2_X1 U536 ( .A1(n276), .A2(n203), .ZN(\ab[5][13] ) );
  NOR2_X1 U537 ( .A1(n279), .A2(n203), .ZN(\ab[5][12] ) );
  NOR2_X1 U538 ( .A1(n282), .A2(n203), .ZN(\ab[5][11] ) );
  NOR2_X1 U539 ( .A1(n285), .A2(n203), .ZN(\ab[5][10] ) );
  NOR2_X1 U540 ( .A1(n315), .A2(n203), .ZN(\ab[5][0] ) );
  NOR2_X1 U541 ( .A1(n288), .A2(n208), .ZN(\ab[4][9] ) );
  NOR2_X1 U542 ( .A1(n291), .A2(n208), .ZN(\ab[4][8] ) );
  NOR2_X1 U543 ( .A1(n294), .A2(n208), .ZN(\ab[4][7] ) );
  NOR2_X1 U544 ( .A1(n297), .A2(n208), .ZN(\ab[4][6] ) );
  NOR2_X1 U545 ( .A1(n300), .A2(n208), .ZN(\ab[4][5] ) );
  NOR2_X1 U546 ( .A1(n303), .A2(n208), .ZN(\ab[4][4] ) );
  NOR2_X1 U547 ( .A1(n306), .A2(n208), .ZN(\ab[4][3] ) );
  NOR2_X1 U548 ( .A1(A[4]), .A2(n222), .ZN(\ab[4][31] ) );
  NOR2_X1 U549 ( .A1(n225), .A2(n207), .ZN(\ab[4][30] ) );
  NOR2_X1 U550 ( .A1(n309), .A2(n207), .ZN(\ab[4][2] ) );
  NOR2_X1 U551 ( .A1(n228), .A2(n207), .ZN(\ab[4][29] ) );
  NOR2_X1 U552 ( .A1(n231), .A2(n207), .ZN(\ab[4][28] ) );
  NOR2_X1 U553 ( .A1(n234), .A2(n207), .ZN(\ab[4][27] ) );
  NOR2_X1 U554 ( .A1(n237), .A2(n207), .ZN(\ab[4][26] ) );
  NOR2_X1 U555 ( .A1(n240), .A2(n207), .ZN(\ab[4][25] ) );
  NOR2_X1 U556 ( .A1(n243), .A2(n207), .ZN(\ab[4][24] ) );
  NOR2_X1 U557 ( .A1(n246), .A2(n207), .ZN(\ab[4][23] ) );
  NOR2_X1 U558 ( .A1(n249), .A2(n207), .ZN(\ab[4][22] ) );
  NOR2_X1 U559 ( .A1(n252), .A2(n207), .ZN(\ab[4][21] ) );
  NOR2_X1 U560 ( .A1(n255), .A2(n207), .ZN(\ab[4][20] ) );
  NOR2_X1 U561 ( .A1(n312), .A2(n206), .ZN(\ab[4][1] ) );
  NOR2_X1 U562 ( .A1(n258), .A2(n206), .ZN(\ab[4][19] ) );
  NOR2_X1 U563 ( .A1(n261), .A2(n206), .ZN(\ab[4][18] ) );
  NOR2_X1 U564 ( .A1(n264), .A2(n206), .ZN(\ab[4][17] ) );
  NOR2_X1 U565 ( .A1(n267), .A2(n206), .ZN(\ab[4][16] ) );
  NOR2_X1 U566 ( .A1(n270), .A2(n206), .ZN(\ab[4][15] ) );
  NOR2_X1 U567 ( .A1(n273), .A2(n206), .ZN(\ab[4][14] ) );
  NOR2_X1 U568 ( .A1(n276), .A2(n206), .ZN(\ab[4][13] ) );
  NOR2_X1 U569 ( .A1(n279), .A2(n206), .ZN(\ab[4][12] ) );
  NOR2_X1 U570 ( .A1(n282), .A2(n206), .ZN(\ab[4][11] ) );
  NOR2_X1 U571 ( .A1(n285), .A2(n206), .ZN(\ab[4][10] ) );
  NOR2_X1 U572 ( .A1(n315), .A2(n206), .ZN(\ab[4][0] ) );
  NOR2_X1 U573 ( .A1(n288), .A2(n211), .ZN(\ab[3][9] ) );
  NOR2_X1 U574 ( .A1(n291), .A2(n211), .ZN(\ab[3][8] ) );
  NOR2_X1 U575 ( .A1(n294), .A2(n211), .ZN(\ab[3][7] ) );
  NOR2_X1 U576 ( .A1(n297), .A2(n211), .ZN(\ab[3][6] ) );
  NOR2_X1 U577 ( .A1(n300), .A2(n211), .ZN(\ab[3][5] ) );
  NOR2_X1 U578 ( .A1(n303), .A2(n211), .ZN(\ab[3][4] ) );
  NOR2_X1 U579 ( .A1(n306), .A2(n211), .ZN(\ab[3][3] ) );
  NOR2_X1 U580 ( .A1(A[3]), .A2(n222), .ZN(\ab[3][31] ) );
  NOR2_X1 U581 ( .A1(n225), .A2(n210), .ZN(\ab[3][30] ) );
  NOR2_X1 U582 ( .A1(n309), .A2(n210), .ZN(\ab[3][2] ) );
  NOR2_X1 U583 ( .A1(n228), .A2(n210), .ZN(\ab[3][29] ) );
  NOR2_X1 U584 ( .A1(n231), .A2(n210), .ZN(\ab[3][28] ) );
  NOR2_X1 U585 ( .A1(n234), .A2(n210), .ZN(\ab[3][27] ) );
  NOR2_X1 U586 ( .A1(n237), .A2(n210), .ZN(\ab[3][26] ) );
  NOR2_X1 U587 ( .A1(n240), .A2(n210), .ZN(\ab[3][25] ) );
  NOR2_X1 U588 ( .A1(n243), .A2(n210), .ZN(\ab[3][24] ) );
  NOR2_X1 U589 ( .A1(n246), .A2(n210), .ZN(\ab[3][23] ) );
  NOR2_X1 U590 ( .A1(n249), .A2(n210), .ZN(\ab[3][22] ) );
  NOR2_X1 U591 ( .A1(n252), .A2(n210), .ZN(\ab[3][21] ) );
  NOR2_X1 U592 ( .A1(n255), .A2(n210), .ZN(\ab[3][20] ) );
  NOR2_X1 U593 ( .A1(n312), .A2(n209), .ZN(\ab[3][1] ) );
  NOR2_X1 U594 ( .A1(n258), .A2(n209), .ZN(\ab[3][19] ) );
  NOR2_X1 U595 ( .A1(n261), .A2(n209), .ZN(\ab[3][18] ) );
  NOR2_X1 U596 ( .A1(n264), .A2(n209), .ZN(\ab[3][17] ) );
  NOR2_X1 U597 ( .A1(n267), .A2(n209), .ZN(\ab[3][16] ) );
  NOR2_X1 U598 ( .A1(n270), .A2(n209), .ZN(\ab[3][15] ) );
  NOR2_X1 U599 ( .A1(n273), .A2(n209), .ZN(\ab[3][14] ) );
  NOR2_X1 U600 ( .A1(n276), .A2(n209), .ZN(\ab[3][13] ) );
  NOR2_X1 U601 ( .A1(n279), .A2(n209), .ZN(\ab[3][12] ) );
  NOR2_X1 U602 ( .A1(n282), .A2(n209), .ZN(\ab[3][11] ) );
  NOR2_X1 U603 ( .A1(n285), .A2(n209), .ZN(\ab[3][10] ) );
  NOR2_X1 U604 ( .A1(n315), .A2(n209), .ZN(\ab[3][0] ) );
  NOR2_X1 U605 ( .A1(B[9]), .A2(n127), .ZN(\ab[31][9] ) );
  NOR2_X1 U606 ( .A1(B[8]), .A2(n127), .ZN(\ab[31][8] ) );
  NOR2_X1 U607 ( .A1(B[7]), .A2(n127), .ZN(\ab[31][7] ) );
  NOR2_X1 U608 ( .A1(B[6]), .A2(n127), .ZN(\ab[31][6] ) );
  NOR2_X1 U609 ( .A1(B[5]), .A2(n127), .ZN(\ab[31][5] ) );
  NOR2_X1 U610 ( .A1(B[4]), .A2(n127), .ZN(\ab[31][4] ) );
  NOR2_X1 U611 ( .A1(B[3]), .A2(n127), .ZN(\ab[31][3] ) );
  NOR2_X1 U612 ( .A1(n221), .A2(n127), .ZN(\ab[31][31] ) );
  NOR2_X1 U613 ( .A1(B[30]), .A2(n127), .ZN(\ab[31][30] ) );
  NOR2_X1 U614 ( .A1(B[2]), .A2(n127), .ZN(\ab[31][2] ) );
  NOR2_X1 U615 ( .A1(B[29]), .A2(n127), .ZN(\ab[31][29] ) );
  NOR2_X1 U616 ( .A1(B[28]), .A2(n127), .ZN(\ab[31][28] ) );
  NOR2_X1 U617 ( .A1(B[27]), .A2(n126), .ZN(\ab[31][27] ) );
  NOR2_X1 U618 ( .A1(B[26]), .A2(n126), .ZN(\ab[31][26] ) );
  NOR2_X1 U619 ( .A1(B[25]), .A2(n126), .ZN(\ab[31][25] ) );
  NOR2_X1 U620 ( .A1(B[24]), .A2(n126), .ZN(\ab[31][24] ) );
  NOR2_X1 U621 ( .A1(B[23]), .A2(n126), .ZN(\ab[31][23] ) );
  NOR2_X1 U622 ( .A1(B[22]), .A2(n126), .ZN(\ab[31][22] ) );
  NOR2_X1 U623 ( .A1(B[21]), .A2(n126), .ZN(\ab[31][21] ) );
  NOR2_X1 U624 ( .A1(B[20]), .A2(n126), .ZN(\ab[31][20] ) );
  NOR2_X1 U625 ( .A1(B[1]), .A2(n126), .ZN(\ab[31][1] ) );
  NOR2_X1 U626 ( .A1(B[19]), .A2(n126), .ZN(\ab[31][19] ) );
  NOR2_X1 U627 ( .A1(B[18]), .A2(n126), .ZN(\ab[31][18] ) );
  NOR2_X1 U628 ( .A1(B[17]), .A2(n126), .ZN(\ab[31][17] ) );
  NOR2_X1 U629 ( .A1(B[16]), .A2(n126), .ZN(\ab[31][16] ) );
  NOR2_X1 U630 ( .A1(B[15]), .A2(n126), .ZN(\ab[31][15] ) );
  NOR2_X1 U631 ( .A1(B[14]), .A2(n126), .ZN(\ab[31][14] ) );
  NOR2_X1 U632 ( .A1(B[13]), .A2(n126), .ZN(\ab[31][13] ) );
  NOR2_X1 U633 ( .A1(B[12]), .A2(n126), .ZN(\ab[31][12] ) );
  NOR2_X1 U634 ( .A1(B[11]), .A2(n126), .ZN(\ab[31][11] ) );
  NOR2_X1 U635 ( .A1(B[10]), .A2(n126), .ZN(\ab[31][10] ) );
  NOR2_X1 U636 ( .A1(B[0]), .A2(n126), .ZN(\ab[31][0] ) );
  NOR2_X1 U637 ( .A1(n287), .A2(n130), .ZN(\ab[30][9] ) );
  NOR2_X1 U638 ( .A1(n290), .A2(n130), .ZN(\ab[30][8] ) );
  NOR2_X1 U639 ( .A1(n293), .A2(n130), .ZN(\ab[30][7] ) );
  NOR2_X1 U640 ( .A1(n296), .A2(n130), .ZN(\ab[30][6] ) );
  NOR2_X1 U641 ( .A1(n299), .A2(n130), .ZN(\ab[30][5] ) );
  NOR2_X1 U642 ( .A1(n302), .A2(n130), .ZN(\ab[30][4] ) );
  NOR2_X1 U643 ( .A1(n305), .A2(n130), .ZN(\ab[30][3] ) );
  NOR2_X1 U644 ( .A1(A[30]), .A2(n222), .ZN(\ab[30][31] ) );
  NOR2_X1 U645 ( .A1(n224), .A2(n129), .ZN(\ab[30][30] ) );
  NOR2_X1 U646 ( .A1(n308), .A2(n129), .ZN(\ab[30][2] ) );
  NOR2_X1 U647 ( .A1(n227), .A2(n129), .ZN(\ab[30][29] ) );
  NOR2_X1 U648 ( .A1(n230), .A2(n129), .ZN(\ab[30][28] ) );
  NOR2_X1 U649 ( .A1(n233), .A2(n129), .ZN(\ab[30][27] ) );
  NOR2_X1 U650 ( .A1(n236), .A2(n129), .ZN(\ab[30][26] ) );
  NOR2_X1 U651 ( .A1(n239), .A2(n129), .ZN(\ab[30][25] ) );
  NOR2_X1 U652 ( .A1(n242), .A2(n129), .ZN(\ab[30][24] ) );
  NOR2_X1 U653 ( .A1(n245), .A2(n129), .ZN(\ab[30][23] ) );
  NOR2_X1 U654 ( .A1(n248), .A2(n129), .ZN(\ab[30][22] ) );
  NOR2_X1 U655 ( .A1(n251), .A2(n129), .ZN(\ab[30][21] ) );
  NOR2_X1 U656 ( .A1(n254), .A2(n129), .ZN(\ab[30][20] ) );
  NOR2_X1 U657 ( .A1(n311), .A2(n128), .ZN(\ab[30][1] ) );
  NOR2_X1 U658 ( .A1(n257), .A2(n128), .ZN(\ab[30][19] ) );
  NOR2_X1 U659 ( .A1(n260), .A2(n128), .ZN(\ab[30][18] ) );
  NOR2_X1 U660 ( .A1(n263), .A2(n128), .ZN(\ab[30][17] ) );
  NOR2_X1 U661 ( .A1(n266), .A2(n128), .ZN(\ab[30][16] ) );
  NOR2_X1 U662 ( .A1(n269), .A2(n128), .ZN(\ab[30][15] ) );
  NOR2_X1 U663 ( .A1(n272), .A2(n128), .ZN(\ab[30][14] ) );
  NOR2_X1 U664 ( .A1(n275), .A2(n128), .ZN(\ab[30][13] ) );
  NOR2_X1 U665 ( .A1(n278), .A2(n128), .ZN(\ab[30][12] ) );
  NOR2_X1 U666 ( .A1(n281), .A2(n128), .ZN(\ab[30][11] ) );
  NOR2_X1 U667 ( .A1(n284), .A2(n128), .ZN(\ab[30][10] ) );
  NOR2_X1 U668 ( .A1(n314), .A2(n128), .ZN(\ab[30][0] ) );
  NOR2_X1 U669 ( .A1(n287), .A2(n214), .ZN(\ab[2][9] ) );
  NOR2_X1 U670 ( .A1(n290), .A2(n214), .ZN(\ab[2][8] ) );
  NOR2_X1 U671 ( .A1(n293), .A2(n214), .ZN(\ab[2][7] ) );
  NOR2_X1 U672 ( .A1(n296), .A2(n214), .ZN(\ab[2][6] ) );
  NOR2_X1 U673 ( .A1(n299), .A2(n214), .ZN(\ab[2][5] ) );
  NOR2_X1 U674 ( .A1(n302), .A2(n214), .ZN(\ab[2][4] ) );
  NOR2_X1 U675 ( .A1(n305), .A2(n214), .ZN(\ab[2][3] ) );
  NOR2_X1 U676 ( .A1(A[2]), .A2(n222), .ZN(\ab[2][31] ) );
  NOR2_X1 U677 ( .A1(n224), .A2(n213), .ZN(\ab[2][30] ) );
  NOR2_X1 U678 ( .A1(n308), .A2(n213), .ZN(\ab[2][2] ) );
  NOR2_X1 U679 ( .A1(n227), .A2(n213), .ZN(\ab[2][29] ) );
  NOR2_X1 U680 ( .A1(n230), .A2(n213), .ZN(\ab[2][28] ) );
  NOR2_X1 U681 ( .A1(n233), .A2(n213), .ZN(\ab[2][27] ) );
  NOR2_X1 U682 ( .A1(n236), .A2(n213), .ZN(\ab[2][26] ) );
  NOR2_X1 U683 ( .A1(n239), .A2(n213), .ZN(\ab[2][25] ) );
  NOR2_X1 U684 ( .A1(n242), .A2(n213), .ZN(\ab[2][24] ) );
  NOR2_X1 U685 ( .A1(n245), .A2(n213), .ZN(\ab[2][23] ) );
  NOR2_X1 U686 ( .A1(n248), .A2(n213), .ZN(\ab[2][22] ) );
  NOR2_X1 U687 ( .A1(n251), .A2(n213), .ZN(\ab[2][21] ) );
  NOR2_X1 U688 ( .A1(n254), .A2(n213), .ZN(\ab[2][20] ) );
  NOR2_X1 U689 ( .A1(n311), .A2(n212), .ZN(\ab[2][1] ) );
  NOR2_X1 U690 ( .A1(n257), .A2(n212), .ZN(\ab[2][19] ) );
  NOR2_X1 U691 ( .A1(n260), .A2(n212), .ZN(\ab[2][18] ) );
  NOR2_X1 U692 ( .A1(n263), .A2(n212), .ZN(\ab[2][17] ) );
  NOR2_X1 U693 ( .A1(n266), .A2(n212), .ZN(\ab[2][16] ) );
  NOR2_X1 U694 ( .A1(n269), .A2(n212), .ZN(\ab[2][15] ) );
  NOR2_X1 U695 ( .A1(n272), .A2(n212), .ZN(\ab[2][14] ) );
  NOR2_X1 U696 ( .A1(n275), .A2(n212), .ZN(\ab[2][13] ) );
  NOR2_X1 U697 ( .A1(n278), .A2(n212), .ZN(\ab[2][12] ) );
  NOR2_X1 U698 ( .A1(n281), .A2(n212), .ZN(\ab[2][11] ) );
  NOR2_X1 U699 ( .A1(n284), .A2(n212), .ZN(\ab[2][10] ) );
  NOR2_X1 U700 ( .A1(n314), .A2(n212), .ZN(\ab[2][0] ) );
  NOR2_X1 U701 ( .A1(n287), .A2(n133), .ZN(\ab[29][9] ) );
  NOR2_X1 U702 ( .A1(n290), .A2(n133), .ZN(\ab[29][8] ) );
  NOR2_X1 U703 ( .A1(n293), .A2(n133), .ZN(\ab[29][7] ) );
  NOR2_X1 U704 ( .A1(n296), .A2(n133), .ZN(\ab[29][6] ) );
  NOR2_X1 U705 ( .A1(n299), .A2(n133), .ZN(\ab[29][5] ) );
  NOR2_X1 U706 ( .A1(n302), .A2(n133), .ZN(\ab[29][4] ) );
  NOR2_X1 U707 ( .A1(n305), .A2(n133), .ZN(\ab[29][3] ) );
  NOR2_X1 U708 ( .A1(A[29]), .A2(n222), .ZN(\ab[29][31] ) );
  NOR2_X1 U709 ( .A1(n224), .A2(n132), .ZN(\ab[29][30] ) );
  NOR2_X1 U710 ( .A1(n308), .A2(n132), .ZN(\ab[29][2] ) );
  NOR2_X1 U711 ( .A1(n227), .A2(n132), .ZN(\ab[29][29] ) );
  NOR2_X1 U712 ( .A1(n230), .A2(n132), .ZN(\ab[29][28] ) );
  NOR2_X1 U713 ( .A1(n233), .A2(n132), .ZN(\ab[29][27] ) );
  NOR2_X1 U714 ( .A1(n236), .A2(n132), .ZN(\ab[29][26] ) );
  NOR2_X1 U715 ( .A1(n239), .A2(n132), .ZN(\ab[29][25] ) );
  NOR2_X1 U716 ( .A1(n242), .A2(n132), .ZN(\ab[29][24] ) );
  NOR2_X1 U717 ( .A1(n245), .A2(n132), .ZN(\ab[29][23] ) );
  NOR2_X1 U718 ( .A1(n248), .A2(n132), .ZN(\ab[29][22] ) );
  NOR2_X1 U719 ( .A1(n251), .A2(n132), .ZN(\ab[29][21] ) );
  NOR2_X1 U720 ( .A1(n254), .A2(n132), .ZN(\ab[29][20] ) );
  NOR2_X1 U721 ( .A1(n311), .A2(n131), .ZN(\ab[29][1] ) );
  NOR2_X1 U722 ( .A1(n257), .A2(n131), .ZN(\ab[29][19] ) );
  NOR2_X1 U723 ( .A1(n260), .A2(n131), .ZN(\ab[29][18] ) );
  NOR2_X1 U724 ( .A1(n263), .A2(n131), .ZN(\ab[29][17] ) );
  NOR2_X1 U725 ( .A1(n266), .A2(n131), .ZN(\ab[29][16] ) );
  NOR2_X1 U726 ( .A1(n269), .A2(n131), .ZN(\ab[29][15] ) );
  NOR2_X1 U727 ( .A1(n272), .A2(n131), .ZN(\ab[29][14] ) );
  NOR2_X1 U728 ( .A1(n275), .A2(n131), .ZN(\ab[29][13] ) );
  NOR2_X1 U729 ( .A1(n278), .A2(n131), .ZN(\ab[29][12] ) );
  NOR2_X1 U730 ( .A1(n281), .A2(n131), .ZN(\ab[29][11] ) );
  NOR2_X1 U731 ( .A1(n284), .A2(n131), .ZN(\ab[29][10] ) );
  NOR2_X1 U732 ( .A1(n314), .A2(n131), .ZN(\ab[29][0] ) );
  NOR2_X1 U733 ( .A1(n287), .A2(n136), .ZN(\ab[28][9] ) );
  NOR2_X1 U734 ( .A1(n290), .A2(n136), .ZN(\ab[28][8] ) );
  NOR2_X1 U735 ( .A1(n293), .A2(n136), .ZN(\ab[28][7] ) );
  NOR2_X1 U736 ( .A1(n296), .A2(n136), .ZN(\ab[28][6] ) );
  NOR2_X1 U737 ( .A1(n299), .A2(n136), .ZN(\ab[28][5] ) );
  NOR2_X1 U738 ( .A1(n302), .A2(n136), .ZN(\ab[28][4] ) );
  NOR2_X1 U739 ( .A1(n305), .A2(n136), .ZN(\ab[28][3] ) );
  NOR2_X1 U740 ( .A1(A[28]), .A2(n222), .ZN(\ab[28][31] ) );
  NOR2_X1 U741 ( .A1(n224), .A2(n135), .ZN(\ab[28][30] ) );
  NOR2_X1 U742 ( .A1(n308), .A2(n135), .ZN(\ab[28][2] ) );
  NOR2_X1 U743 ( .A1(n227), .A2(n135), .ZN(\ab[28][29] ) );
  NOR2_X1 U744 ( .A1(n230), .A2(n135), .ZN(\ab[28][28] ) );
  NOR2_X1 U745 ( .A1(n233), .A2(n135), .ZN(\ab[28][27] ) );
  NOR2_X1 U746 ( .A1(n236), .A2(n135), .ZN(\ab[28][26] ) );
  NOR2_X1 U747 ( .A1(n239), .A2(n135), .ZN(\ab[28][25] ) );
  NOR2_X1 U748 ( .A1(n242), .A2(n135), .ZN(\ab[28][24] ) );
  NOR2_X1 U749 ( .A1(n245), .A2(n135), .ZN(\ab[28][23] ) );
  NOR2_X1 U750 ( .A1(n248), .A2(n135), .ZN(\ab[28][22] ) );
  NOR2_X1 U751 ( .A1(n251), .A2(n135), .ZN(\ab[28][21] ) );
  NOR2_X1 U752 ( .A1(n254), .A2(n135), .ZN(\ab[28][20] ) );
  NOR2_X1 U753 ( .A1(n311), .A2(n134), .ZN(\ab[28][1] ) );
  NOR2_X1 U754 ( .A1(n257), .A2(n134), .ZN(\ab[28][19] ) );
  NOR2_X1 U755 ( .A1(n260), .A2(n134), .ZN(\ab[28][18] ) );
  NOR2_X1 U756 ( .A1(n263), .A2(n134), .ZN(\ab[28][17] ) );
  NOR2_X1 U757 ( .A1(n266), .A2(n134), .ZN(\ab[28][16] ) );
  NOR2_X1 U758 ( .A1(n269), .A2(n134), .ZN(\ab[28][15] ) );
  NOR2_X1 U759 ( .A1(n272), .A2(n134), .ZN(\ab[28][14] ) );
  NOR2_X1 U760 ( .A1(n275), .A2(n134), .ZN(\ab[28][13] ) );
  NOR2_X1 U761 ( .A1(n278), .A2(n134), .ZN(\ab[28][12] ) );
  NOR2_X1 U762 ( .A1(n281), .A2(n134), .ZN(\ab[28][11] ) );
  NOR2_X1 U763 ( .A1(n284), .A2(n134), .ZN(\ab[28][10] ) );
  NOR2_X1 U764 ( .A1(n314), .A2(n134), .ZN(\ab[28][0] ) );
  NOR2_X1 U765 ( .A1(n287), .A2(n139), .ZN(\ab[27][9] ) );
  NOR2_X1 U766 ( .A1(n290), .A2(n139), .ZN(\ab[27][8] ) );
  NOR2_X1 U767 ( .A1(n293), .A2(n139), .ZN(\ab[27][7] ) );
  NOR2_X1 U768 ( .A1(n296), .A2(n139), .ZN(\ab[27][6] ) );
  NOR2_X1 U769 ( .A1(n299), .A2(n139), .ZN(\ab[27][5] ) );
  NOR2_X1 U770 ( .A1(n302), .A2(n139), .ZN(\ab[27][4] ) );
  NOR2_X1 U771 ( .A1(n305), .A2(n139), .ZN(\ab[27][3] ) );
  NOR2_X1 U772 ( .A1(A[27]), .A2(n222), .ZN(\ab[27][31] ) );
  NOR2_X1 U773 ( .A1(n224), .A2(n138), .ZN(\ab[27][30] ) );
  NOR2_X1 U774 ( .A1(n308), .A2(n138), .ZN(\ab[27][2] ) );
  NOR2_X1 U775 ( .A1(n227), .A2(n138), .ZN(\ab[27][29] ) );
  NOR2_X1 U776 ( .A1(n230), .A2(n138), .ZN(\ab[27][28] ) );
  NOR2_X1 U777 ( .A1(n233), .A2(n138), .ZN(\ab[27][27] ) );
  NOR2_X1 U778 ( .A1(n236), .A2(n138), .ZN(\ab[27][26] ) );
  NOR2_X1 U779 ( .A1(n239), .A2(n138), .ZN(\ab[27][25] ) );
  NOR2_X1 U780 ( .A1(n242), .A2(n138), .ZN(\ab[27][24] ) );
  NOR2_X1 U781 ( .A1(n245), .A2(n138), .ZN(\ab[27][23] ) );
  NOR2_X1 U782 ( .A1(n248), .A2(n138), .ZN(\ab[27][22] ) );
  NOR2_X1 U783 ( .A1(n251), .A2(n138), .ZN(\ab[27][21] ) );
  NOR2_X1 U784 ( .A1(n254), .A2(n138), .ZN(\ab[27][20] ) );
  NOR2_X1 U785 ( .A1(n311), .A2(n137), .ZN(\ab[27][1] ) );
  NOR2_X1 U786 ( .A1(n257), .A2(n137), .ZN(\ab[27][19] ) );
  NOR2_X1 U787 ( .A1(n260), .A2(n137), .ZN(\ab[27][18] ) );
  NOR2_X1 U788 ( .A1(n263), .A2(n137), .ZN(\ab[27][17] ) );
  NOR2_X1 U789 ( .A1(n266), .A2(n137), .ZN(\ab[27][16] ) );
  NOR2_X1 U790 ( .A1(n269), .A2(n137), .ZN(\ab[27][15] ) );
  NOR2_X1 U791 ( .A1(n272), .A2(n137), .ZN(\ab[27][14] ) );
  NOR2_X1 U792 ( .A1(n275), .A2(n137), .ZN(\ab[27][13] ) );
  NOR2_X1 U793 ( .A1(n278), .A2(n137), .ZN(\ab[27][12] ) );
  NOR2_X1 U794 ( .A1(n281), .A2(n137), .ZN(\ab[27][11] ) );
  NOR2_X1 U795 ( .A1(n284), .A2(n137), .ZN(\ab[27][10] ) );
  NOR2_X1 U796 ( .A1(n314), .A2(n137), .ZN(\ab[27][0] ) );
  NOR2_X1 U797 ( .A1(n287), .A2(n142), .ZN(\ab[26][9] ) );
  NOR2_X1 U798 ( .A1(n290), .A2(n142), .ZN(\ab[26][8] ) );
  NOR2_X1 U799 ( .A1(n293), .A2(n142), .ZN(\ab[26][7] ) );
  NOR2_X1 U800 ( .A1(n296), .A2(n142), .ZN(\ab[26][6] ) );
  NOR2_X1 U801 ( .A1(n299), .A2(n142), .ZN(\ab[26][5] ) );
  NOR2_X1 U802 ( .A1(n302), .A2(n142), .ZN(\ab[26][4] ) );
  NOR2_X1 U803 ( .A1(n305), .A2(n142), .ZN(\ab[26][3] ) );
  NOR2_X1 U804 ( .A1(A[26]), .A2(n222), .ZN(\ab[26][31] ) );
  NOR2_X1 U805 ( .A1(n224), .A2(n141), .ZN(\ab[26][30] ) );
  NOR2_X1 U806 ( .A1(n308), .A2(n141), .ZN(\ab[26][2] ) );
  NOR2_X1 U807 ( .A1(n227), .A2(n141), .ZN(\ab[26][29] ) );
  NOR2_X1 U808 ( .A1(n230), .A2(n141), .ZN(\ab[26][28] ) );
  NOR2_X1 U809 ( .A1(n233), .A2(n141), .ZN(\ab[26][27] ) );
  NOR2_X1 U810 ( .A1(n236), .A2(n141), .ZN(\ab[26][26] ) );
  NOR2_X1 U811 ( .A1(n239), .A2(n141), .ZN(\ab[26][25] ) );
  NOR2_X1 U812 ( .A1(n242), .A2(n141), .ZN(\ab[26][24] ) );
  NOR2_X1 U813 ( .A1(n245), .A2(n141), .ZN(\ab[26][23] ) );
  NOR2_X1 U814 ( .A1(n248), .A2(n141), .ZN(\ab[26][22] ) );
  NOR2_X1 U815 ( .A1(n251), .A2(n141), .ZN(\ab[26][21] ) );
  NOR2_X1 U816 ( .A1(n254), .A2(n141), .ZN(\ab[26][20] ) );
  NOR2_X1 U817 ( .A1(n311), .A2(n140), .ZN(\ab[26][1] ) );
  NOR2_X1 U818 ( .A1(n257), .A2(n140), .ZN(\ab[26][19] ) );
  NOR2_X1 U819 ( .A1(n260), .A2(n140), .ZN(\ab[26][18] ) );
  NOR2_X1 U820 ( .A1(n263), .A2(n140), .ZN(\ab[26][17] ) );
  NOR2_X1 U821 ( .A1(n266), .A2(n140), .ZN(\ab[26][16] ) );
  NOR2_X1 U822 ( .A1(n269), .A2(n140), .ZN(\ab[26][15] ) );
  NOR2_X1 U823 ( .A1(n272), .A2(n140), .ZN(\ab[26][14] ) );
  NOR2_X1 U824 ( .A1(n275), .A2(n140), .ZN(\ab[26][13] ) );
  NOR2_X1 U825 ( .A1(n278), .A2(n140), .ZN(\ab[26][12] ) );
  NOR2_X1 U826 ( .A1(n281), .A2(n140), .ZN(\ab[26][11] ) );
  NOR2_X1 U827 ( .A1(n284), .A2(n140), .ZN(\ab[26][10] ) );
  NOR2_X1 U828 ( .A1(n314), .A2(n140), .ZN(\ab[26][0] ) );
  NOR2_X1 U829 ( .A1(n287), .A2(n145), .ZN(\ab[25][9] ) );
  NOR2_X1 U830 ( .A1(n290), .A2(n145), .ZN(\ab[25][8] ) );
  NOR2_X1 U831 ( .A1(n293), .A2(n145), .ZN(\ab[25][7] ) );
  NOR2_X1 U832 ( .A1(n296), .A2(n145), .ZN(\ab[25][6] ) );
  NOR2_X1 U833 ( .A1(n299), .A2(n145), .ZN(\ab[25][5] ) );
  NOR2_X1 U834 ( .A1(n302), .A2(n145), .ZN(\ab[25][4] ) );
  NOR2_X1 U835 ( .A1(n305), .A2(n145), .ZN(\ab[25][3] ) );
  NOR2_X1 U836 ( .A1(A[25]), .A2(n222), .ZN(\ab[25][31] ) );
  NOR2_X1 U837 ( .A1(n224), .A2(n144), .ZN(\ab[25][30] ) );
  NOR2_X1 U838 ( .A1(n308), .A2(n144), .ZN(\ab[25][2] ) );
  NOR2_X1 U839 ( .A1(n227), .A2(n144), .ZN(\ab[25][29] ) );
  NOR2_X1 U840 ( .A1(n230), .A2(n144), .ZN(\ab[25][28] ) );
  NOR2_X1 U841 ( .A1(n233), .A2(n144), .ZN(\ab[25][27] ) );
  NOR2_X1 U842 ( .A1(n236), .A2(n144), .ZN(\ab[25][26] ) );
  NOR2_X1 U843 ( .A1(n239), .A2(n144), .ZN(\ab[25][25] ) );
  NOR2_X1 U844 ( .A1(n242), .A2(n144), .ZN(\ab[25][24] ) );
  NOR2_X1 U845 ( .A1(n245), .A2(n144), .ZN(\ab[25][23] ) );
  NOR2_X1 U846 ( .A1(n248), .A2(n144), .ZN(\ab[25][22] ) );
  NOR2_X1 U847 ( .A1(n251), .A2(n144), .ZN(\ab[25][21] ) );
  NOR2_X1 U848 ( .A1(n254), .A2(n144), .ZN(\ab[25][20] ) );
  NOR2_X1 U849 ( .A1(n311), .A2(n143), .ZN(\ab[25][1] ) );
  NOR2_X1 U850 ( .A1(n257), .A2(n143), .ZN(\ab[25][19] ) );
  NOR2_X1 U851 ( .A1(n260), .A2(n143), .ZN(\ab[25][18] ) );
  NOR2_X1 U852 ( .A1(n263), .A2(n143), .ZN(\ab[25][17] ) );
  NOR2_X1 U853 ( .A1(n266), .A2(n143), .ZN(\ab[25][16] ) );
  NOR2_X1 U854 ( .A1(n269), .A2(n143), .ZN(\ab[25][15] ) );
  NOR2_X1 U855 ( .A1(n272), .A2(n143), .ZN(\ab[25][14] ) );
  NOR2_X1 U856 ( .A1(n275), .A2(n143), .ZN(\ab[25][13] ) );
  NOR2_X1 U857 ( .A1(n278), .A2(n143), .ZN(\ab[25][12] ) );
  NOR2_X1 U858 ( .A1(n281), .A2(n143), .ZN(\ab[25][11] ) );
  NOR2_X1 U859 ( .A1(n284), .A2(n143), .ZN(\ab[25][10] ) );
  NOR2_X1 U860 ( .A1(n314), .A2(n143), .ZN(\ab[25][0] ) );
  NOR2_X1 U861 ( .A1(n287), .A2(n148), .ZN(\ab[24][9] ) );
  NOR2_X1 U862 ( .A1(n290), .A2(n148), .ZN(\ab[24][8] ) );
  NOR2_X1 U863 ( .A1(n293), .A2(n148), .ZN(\ab[24][7] ) );
  NOR2_X1 U864 ( .A1(n296), .A2(n148), .ZN(\ab[24][6] ) );
  NOR2_X1 U865 ( .A1(n299), .A2(n148), .ZN(\ab[24][5] ) );
  NOR2_X1 U866 ( .A1(n302), .A2(n148), .ZN(\ab[24][4] ) );
  NOR2_X1 U867 ( .A1(n305), .A2(n148), .ZN(\ab[24][3] ) );
  NOR2_X1 U868 ( .A1(A[24]), .A2(n221), .ZN(\ab[24][31] ) );
  NOR2_X1 U869 ( .A1(n224), .A2(n147), .ZN(\ab[24][30] ) );
  NOR2_X1 U870 ( .A1(n308), .A2(n147), .ZN(\ab[24][2] ) );
  NOR2_X1 U871 ( .A1(n227), .A2(n147), .ZN(\ab[24][29] ) );
  NOR2_X1 U872 ( .A1(n230), .A2(n147), .ZN(\ab[24][28] ) );
  NOR2_X1 U873 ( .A1(n233), .A2(n147), .ZN(\ab[24][27] ) );
  NOR2_X1 U874 ( .A1(n236), .A2(n147), .ZN(\ab[24][26] ) );
  NOR2_X1 U875 ( .A1(n239), .A2(n147), .ZN(\ab[24][25] ) );
  NOR2_X1 U876 ( .A1(n242), .A2(n147), .ZN(\ab[24][24] ) );
  NOR2_X1 U877 ( .A1(n245), .A2(n147), .ZN(\ab[24][23] ) );
  NOR2_X1 U878 ( .A1(n248), .A2(n147), .ZN(\ab[24][22] ) );
  NOR2_X1 U879 ( .A1(n251), .A2(n147), .ZN(\ab[24][21] ) );
  NOR2_X1 U880 ( .A1(n254), .A2(n147), .ZN(\ab[24][20] ) );
  NOR2_X1 U881 ( .A1(n311), .A2(n146), .ZN(\ab[24][1] ) );
  NOR2_X1 U882 ( .A1(n257), .A2(n146), .ZN(\ab[24][19] ) );
  NOR2_X1 U883 ( .A1(n260), .A2(n146), .ZN(\ab[24][18] ) );
  NOR2_X1 U884 ( .A1(n263), .A2(n146), .ZN(\ab[24][17] ) );
  NOR2_X1 U885 ( .A1(n266), .A2(n146), .ZN(\ab[24][16] ) );
  NOR2_X1 U886 ( .A1(n269), .A2(n146), .ZN(\ab[24][15] ) );
  NOR2_X1 U887 ( .A1(n272), .A2(n146), .ZN(\ab[24][14] ) );
  NOR2_X1 U888 ( .A1(n275), .A2(n146), .ZN(\ab[24][13] ) );
  NOR2_X1 U889 ( .A1(n278), .A2(n146), .ZN(\ab[24][12] ) );
  NOR2_X1 U890 ( .A1(n281), .A2(n146), .ZN(\ab[24][11] ) );
  NOR2_X1 U891 ( .A1(n284), .A2(n146), .ZN(\ab[24][10] ) );
  NOR2_X1 U892 ( .A1(n314), .A2(n146), .ZN(\ab[24][0] ) );
  NOR2_X1 U893 ( .A1(n287), .A2(n151), .ZN(\ab[23][9] ) );
  NOR2_X1 U894 ( .A1(n290), .A2(n151), .ZN(\ab[23][8] ) );
  NOR2_X1 U895 ( .A1(n293), .A2(n151), .ZN(\ab[23][7] ) );
  NOR2_X1 U896 ( .A1(n296), .A2(n151), .ZN(\ab[23][6] ) );
  NOR2_X1 U897 ( .A1(n299), .A2(n151), .ZN(\ab[23][5] ) );
  NOR2_X1 U898 ( .A1(n302), .A2(n151), .ZN(\ab[23][4] ) );
  NOR2_X1 U899 ( .A1(n305), .A2(n151), .ZN(\ab[23][3] ) );
  NOR2_X1 U900 ( .A1(A[23]), .A2(n221), .ZN(\ab[23][31] ) );
  NOR2_X1 U901 ( .A1(n224), .A2(n150), .ZN(\ab[23][30] ) );
  NOR2_X1 U902 ( .A1(n308), .A2(n150), .ZN(\ab[23][2] ) );
  NOR2_X1 U903 ( .A1(n227), .A2(n150), .ZN(\ab[23][29] ) );
  NOR2_X1 U904 ( .A1(n230), .A2(n150), .ZN(\ab[23][28] ) );
  NOR2_X1 U905 ( .A1(n233), .A2(n150), .ZN(\ab[23][27] ) );
  NOR2_X1 U906 ( .A1(n236), .A2(n150), .ZN(\ab[23][26] ) );
  NOR2_X1 U907 ( .A1(n239), .A2(n150), .ZN(\ab[23][25] ) );
  NOR2_X1 U908 ( .A1(n242), .A2(n150), .ZN(\ab[23][24] ) );
  NOR2_X1 U909 ( .A1(n245), .A2(n150), .ZN(\ab[23][23] ) );
  NOR2_X1 U910 ( .A1(n248), .A2(n150), .ZN(\ab[23][22] ) );
  NOR2_X1 U911 ( .A1(n251), .A2(n150), .ZN(\ab[23][21] ) );
  NOR2_X1 U912 ( .A1(n254), .A2(n150), .ZN(\ab[23][20] ) );
  NOR2_X1 U913 ( .A1(n311), .A2(n149), .ZN(\ab[23][1] ) );
  NOR2_X1 U914 ( .A1(n257), .A2(n149), .ZN(\ab[23][19] ) );
  NOR2_X1 U915 ( .A1(n260), .A2(n149), .ZN(\ab[23][18] ) );
  NOR2_X1 U916 ( .A1(n263), .A2(n149), .ZN(\ab[23][17] ) );
  NOR2_X1 U917 ( .A1(n266), .A2(n149), .ZN(\ab[23][16] ) );
  NOR2_X1 U918 ( .A1(n269), .A2(n149), .ZN(\ab[23][15] ) );
  NOR2_X1 U919 ( .A1(n272), .A2(n149), .ZN(\ab[23][14] ) );
  NOR2_X1 U920 ( .A1(n275), .A2(n149), .ZN(\ab[23][13] ) );
  NOR2_X1 U921 ( .A1(n278), .A2(n149), .ZN(\ab[23][12] ) );
  NOR2_X1 U922 ( .A1(n281), .A2(n149), .ZN(\ab[23][11] ) );
  NOR2_X1 U923 ( .A1(n284), .A2(n149), .ZN(\ab[23][10] ) );
  NOR2_X1 U924 ( .A1(n314), .A2(n149), .ZN(\ab[23][0] ) );
  NOR2_X1 U925 ( .A1(n287), .A2(n154), .ZN(\ab[22][9] ) );
  NOR2_X1 U926 ( .A1(n290), .A2(n154), .ZN(\ab[22][8] ) );
  NOR2_X1 U927 ( .A1(n293), .A2(n154), .ZN(\ab[22][7] ) );
  NOR2_X1 U928 ( .A1(n296), .A2(n154), .ZN(\ab[22][6] ) );
  NOR2_X1 U929 ( .A1(n299), .A2(n154), .ZN(\ab[22][5] ) );
  NOR2_X1 U930 ( .A1(n302), .A2(n154), .ZN(\ab[22][4] ) );
  NOR2_X1 U931 ( .A1(n305), .A2(n154), .ZN(\ab[22][3] ) );
  NOR2_X1 U932 ( .A1(A[22]), .A2(n221), .ZN(\ab[22][31] ) );
  NOR2_X1 U933 ( .A1(n224), .A2(n153), .ZN(\ab[22][30] ) );
  NOR2_X1 U934 ( .A1(n308), .A2(n153), .ZN(\ab[22][2] ) );
  NOR2_X1 U935 ( .A1(n227), .A2(n153), .ZN(\ab[22][29] ) );
  NOR2_X1 U936 ( .A1(n230), .A2(n153), .ZN(\ab[22][28] ) );
  NOR2_X1 U937 ( .A1(n233), .A2(n153), .ZN(\ab[22][27] ) );
  NOR2_X1 U938 ( .A1(n236), .A2(n153), .ZN(\ab[22][26] ) );
  NOR2_X1 U939 ( .A1(n239), .A2(n153), .ZN(\ab[22][25] ) );
  NOR2_X1 U940 ( .A1(n242), .A2(n153), .ZN(\ab[22][24] ) );
  NOR2_X1 U941 ( .A1(n245), .A2(n153), .ZN(\ab[22][23] ) );
  NOR2_X1 U942 ( .A1(n248), .A2(n153), .ZN(\ab[22][22] ) );
  NOR2_X1 U943 ( .A1(n251), .A2(n153), .ZN(\ab[22][21] ) );
  NOR2_X1 U944 ( .A1(n254), .A2(n153), .ZN(\ab[22][20] ) );
  NOR2_X1 U945 ( .A1(n311), .A2(n152), .ZN(\ab[22][1] ) );
  NOR2_X1 U946 ( .A1(n257), .A2(n152), .ZN(\ab[22][19] ) );
  NOR2_X1 U947 ( .A1(n260), .A2(n152), .ZN(\ab[22][18] ) );
  NOR2_X1 U948 ( .A1(n263), .A2(n152), .ZN(\ab[22][17] ) );
  NOR2_X1 U949 ( .A1(n266), .A2(n152), .ZN(\ab[22][16] ) );
  NOR2_X1 U950 ( .A1(n269), .A2(n152), .ZN(\ab[22][15] ) );
  NOR2_X1 U951 ( .A1(n272), .A2(n152), .ZN(\ab[22][14] ) );
  NOR2_X1 U952 ( .A1(n275), .A2(n152), .ZN(\ab[22][13] ) );
  NOR2_X1 U953 ( .A1(n278), .A2(n152), .ZN(\ab[22][12] ) );
  NOR2_X1 U954 ( .A1(n281), .A2(n152), .ZN(\ab[22][11] ) );
  NOR2_X1 U955 ( .A1(n284), .A2(n152), .ZN(\ab[22][10] ) );
  NOR2_X1 U956 ( .A1(n314), .A2(n152), .ZN(\ab[22][0] ) );
  NOR2_X1 U957 ( .A1(n287), .A2(n157), .ZN(\ab[21][9] ) );
  NOR2_X1 U958 ( .A1(n290), .A2(n157), .ZN(\ab[21][8] ) );
  NOR2_X1 U959 ( .A1(n293), .A2(n157), .ZN(\ab[21][7] ) );
  NOR2_X1 U960 ( .A1(n296), .A2(n157), .ZN(\ab[21][6] ) );
  NOR2_X1 U961 ( .A1(n299), .A2(n157), .ZN(\ab[21][5] ) );
  NOR2_X1 U962 ( .A1(n302), .A2(n157), .ZN(\ab[21][4] ) );
  NOR2_X1 U963 ( .A1(n305), .A2(n157), .ZN(\ab[21][3] ) );
  NOR2_X1 U964 ( .A1(A[21]), .A2(n221), .ZN(\ab[21][31] ) );
  NOR2_X1 U965 ( .A1(n224), .A2(n156), .ZN(\ab[21][30] ) );
  NOR2_X1 U966 ( .A1(n308), .A2(n156), .ZN(\ab[21][2] ) );
  NOR2_X1 U967 ( .A1(n227), .A2(n156), .ZN(\ab[21][29] ) );
  NOR2_X1 U968 ( .A1(n230), .A2(n156), .ZN(\ab[21][28] ) );
  NOR2_X1 U969 ( .A1(n233), .A2(n156), .ZN(\ab[21][27] ) );
  NOR2_X1 U970 ( .A1(n236), .A2(n156), .ZN(\ab[21][26] ) );
  NOR2_X1 U971 ( .A1(n239), .A2(n156), .ZN(\ab[21][25] ) );
  NOR2_X1 U972 ( .A1(n242), .A2(n156), .ZN(\ab[21][24] ) );
  NOR2_X1 U973 ( .A1(n245), .A2(n156), .ZN(\ab[21][23] ) );
  NOR2_X1 U974 ( .A1(n248), .A2(n156), .ZN(\ab[21][22] ) );
  NOR2_X1 U975 ( .A1(n251), .A2(n156), .ZN(\ab[21][21] ) );
  NOR2_X1 U976 ( .A1(n254), .A2(n156), .ZN(\ab[21][20] ) );
  NOR2_X1 U977 ( .A1(n311), .A2(n155), .ZN(\ab[21][1] ) );
  NOR2_X1 U978 ( .A1(n257), .A2(n155), .ZN(\ab[21][19] ) );
  NOR2_X1 U979 ( .A1(n260), .A2(n155), .ZN(\ab[21][18] ) );
  NOR2_X1 U980 ( .A1(n263), .A2(n155), .ZN(\ab[21][17] ) );
  NOR2_X1 U981 ( .A1(n266), .A2(n155), .ZN(\ab[21][16] ) );
  NOR2_X1 U982 ( .A1(n269), .A2(n155), .ZN(\ab[21][15] ) );
  NOR2_X1 U983 ( .A1(n272), .A2(n155), .ZN(\ab[21][14] ) );
  NOR2_X1 U984 ( .A1(n275), .A2(n155), .ZN(\ab[21][13] ) );
  NOR2_X1 U985 ( .A1(n278), .A2(n155), .ZN(\ab[21][12] ) );
  NOR2_X1 U986 ( .A1(n281), .A2(n155), .ZN(\ab[21][11] ) );
  NOR2_X1 U987 ( .A1(n284), .A2(n155), .ZN(\ab[21][10] ) );
  NOR2_X1 U988 ( .A1(n314), .A2(n155), .ZN(\ab[21][0] ) );
  NOR2_X1 U989 ( .A1(n287), .A2(n160), .ZN(\ab[20][9] ) );
  NOR2_X1 U990 ( .A1(n290), .A2(n160), .ZN(\ab[20][8] ) );
  NOR2_X1 U991 ( .A1(n293), .A2(n160), .ZN(\ab[20][7] ) );
  NOR2_X1 U992 ( .A1(n296), .A2(n160), .ZN(\ab[20][6] ) );
  NOR2_X1 U993 ( .A1(n299), .A2(n160), .ZN(\ab[20][5] ) );
  NOR2_X1 U994 ( .A1(n302), .A2(n160), .ZN(\ab[20][4] ) );
  NOR2_X1 U995 ( .A1(n305), .A2(n160), .ZN(\ab[20][3] ) );
  NOR2_X1 U996 ( .A1(A[20]), .A2(n221), .ZN(\ab[20][31] ) );
  NOR2_X1 U997 ( .A1(n224), .A2(n159), .ZN(\ab[20][30] ) );
  NOR2_X1 U998 ( .A1(n308), .A2(n159), .ZN(\ab[20][2] ) );
  NOR2_X1 U999 ( .A1(n227), .A2(n159), .ZN(\ab[20][29] ) );
  NOR2_X1 U1000 ( .A1(n230), .A2(n159), .ZN(\ab[20][28] ) );
  NOR2_X1 U1001 ( .A1(n233), .A2(n159), .ZN(\ab[20][27] ) );
  NOR2_X1 U1002 ( .A1(n236), .A2(n159), .ZN(\ab[20][26] ) );
  NOR2_X1 U1003 ( .A1(n239), .A2(n159), .ZN(\ab[20][25] ) );
  NOR2_X1 U1004 ( .A1(n242), .A2(n159), .ZN(\ab[20][24] ) );
  NOR2_X1 U1005 ( .A1(n245), .A2(n159), .ZN(\ab[20][23] ) );
  NOR2_X1 U1006 ( .A1(n248), .A2(n159), .ZN(\ab[20][22] ) );
  NOR2_X1 U1007 ( .A1(n251), .A2(n159), .ZN(\ab[20][21] ) );
  NOR2_X1 U1008 ( .A1(n254), .A2(n159), .ZN(\ab[20][20] ) );
  NOR2_X1 U1009 ( .A1(n311), .A2(n158), .ZN(\ab[20][1] ) );
  NOR2_X1 U1010 ( .A1(n257), .A2(n158), .ZN(\ab[20][19] ) );
  NOR2_X1 U1011 ( .A1(n260), .A2(n158), .ZN(\ab[20][18] ) );
  NOR2_X1 U1012 ( .A1(n263), .A2(n158), .ZN(\ab[20][17] ) );
  NOR2_X1 U1013 ( .A1(n266), .A2(n158), .ZN(\ab[20][16] ) );
  NOR2_X1 U1014 ( .A1(n269), .A2(n158), .ZN(\ab[20][15] ) );
  NOR2_X1 U1015 ( .A1(n272), .A2(n158), .ZN(\ab[20][14] ) );
  NOR2_X1 U1016 ( .A1(n275), .A2(n158), .ZN(\ab[20][13] ) );
  NOR2_X1 U1017 ( .A1(n278), .A2(n158), .ZN(\ab[20][12] ) );
  NOR2_X1 U1018 ( .A1(n281), .A2(n158), .ZN(\ab[20][11] ) );
  NOR2_X1 U1019 ( .A1(n284), .A2(n158), .ZN(\ab[20][10] ) );
  NOR2_X1 U1020 ( .A1(n314), .A2(n158), .ZN(\ab[20][0] ) );
  NOR2_X1 U1021 ( .A1(n286), .A2(n217), .ZN(\ab[1][9] ) );
  NOR2_X1 U1022 ( .A1(n289), .A2(n217), .ZN(\ab[1][8] ) );
  NOR2_X1 U1023 ( .A1(n292), .A2(n217), .ZN(\ab[1][7] ) );
  NOR2_X1 U1024 ( .A1(n295), .A2(n217), .ZN(\ab[1][6] ) );
  NOR2_X1 U1025 ( .A1(n298), .A2(n217), .ZN(\ab[1][5] ) );
  NOR2_X1 U1026 ( .A1(n301), .A2(n217), .ZN(\ab[1][4] ) );
  NOR2_X1 U1027 ( .A1(n304), .A2(n217), .ZN(\ab[1][3] ) );
  NOR2_X1 U1028 ( .A1(A[1]), .A2(n221), .ZN(\ab[1][31] ) );
  NOR2_X1 U1029 ( .A1(n223), .A2(n216), .ZN(\ab[1][30] ) );
  NOR2_X1 U1030 ( .A1(n307), .A2(n216), .ZN(\ab[1][2] ) );
  NOR2_X1 U1031 ( .A1(n226), .A2(n216), .ZN(\ab[1][29] ) );
  NOR2_X1 U1032 ( .A1(n229), .A2(n216), .ZN(\ab[1][28] ) );
  NOR2_X1 U1033 ( .A1(n232), .A2(n216), .ZN(\ab[1][27] ) );
  NOR2_X1 U1034 ( .A1(n235), .A2(n216), .ZN(\ab[1][26] ) );
  NOR2_X1 U1035 ( .A1(n238), .A2(n216), .ZN(\ab[1][25] ) );
  NOR2_X1 U1036 ( .A1(n241), .A2(n216), .ZN(\ab[1][24] ) );
  NOR2_X1 U1037 ( .A1(n244), .A2(n216), .ZN(\ab[1][23] ) );
  NOR2_X1 U1038 ( .A1(n247), .A2(n216), .ZN(\ab[1][22] ) );
  NOR2_X1 U1039 ( .A1(n250), .A2(n216), .ZN(\ab[1][21] ) );
  NOR2_X1 U1040 ( .A1(n253), .A2(n216), .ZN(\ab[1][20] ) );
  NOR2_X1 U1041 ( .A1(n310), .A2(n215), .ZN(\ab[1][1] ) );
  NOR2_X1 U1042 ( .A1(n256), .A2(n215), .ZN(\ab[1][19] ) );
  NOR2_X1 U1043 ( .A1(n259), .A2(n215), .ZN(\ab[1][18] ) );
  NOR2_X1 U1044 ( .A1(n262), .A2(n215), .ZN(\ab[1][17] ) );
  NOR2_X1 U1045 ( .A1(n265), .A2(n215), .ZN(\ab[1][16] ) );
  NOR2_X1 U1046 ( .A1(n268), .A2(n215), .ZN(\ab[1][15] ) );
  NOR2_X1 U1047 ( .A1(n271), .A2(n215), .ZN(\ab[1][14] ) );
  NOR2_X1 U1048 ( .A1(n274), .A2(n215), .ZN(\ab[1][13] ) );
  NOR2_X1 U1049 ( .A1(n277), .A2(n215), .ZN(\ab[1][12] ) );
  NOR2_X1 U1050 ( .A1(n280), .A2(n215), .ZN(\ab[1][11] ) );
  NOR2_X1 U1051 ( .A1(n283), .A2(n215), .ZN(\ab[1][10] ) );
  NOR2_X1 U1052 ( .A1(n313), .A2(n215), .ZN(\ab[1][0] ) );
  NOR2_X1 U1053 ( .A1(n286), .A2(n163), .ZN(\ab[19][9] ) );
  NOR2_X1 U1054 ( .A1(n289), .A2(n163), .ZN(\ab[19][8] ) );
  NOR2_X1 U1055 ( .A1(n292), .A2(n163), .ZN(\ab[19][7] ) );
  NOR2_X1 U1056 ( .A1(n295), .A2(n163), .ZN(\ab[19][6] ) );
  NOR2_X1 U1057 ( .A1(n298), .A2(n163), .ZN(\ab[19][5] ) );
  NOR2_X1 U1058 ( .A1(n301), .A2(n163), .ZN(\ab[19][4] ) );
  NOR2_X1 U1059 ( .A1(n304), .A2(n163), .ZN(\ab[19][3] ) );
  NOR2_X1 U1060 ( .A1(A[19]), .A2(n221), .ZN(\ab[19][31] ) );
  NOR2_X1 U1061 ( .A1(n223), .A2(n162), .ZN(\ab[19][30] ) );
  NOR2_X1 U1062 ( .A1(n307), .A2(n162), .ZN(\ab[19][2] ) );
  NOR2_X1 U1063 ( .A1(n226), .A2(n162), .ZN(\ab[19][29] ) );
  NOR2_X1 U1064 ( .A1(n229), .A2(n162), .ZN(\ab[19][28] ) );
  NOR2_X1 U1065 ( .A1(n232), .A2(n162), .ZN(\ab[19][27] ) );
  NOR2_X1 U1066 ( .A1(n235), .A2(n162), .ZN(\ab[19][26] ) );
  NOR2_X1 U1067 ( .A1(n238), .A2(n162), .ZN(\ab[19][25] ) );
  NOR2_X1 U1068 ( .A1(n241), .A2(n162), .ZN(\ab[19][24] ) );
  NOR2_X1 U1069 ( .A1(n244), .A2(n162), .ZN(\ab[19][23] ) );
  NOR2_X1 U1070 ( .A1(n247), .A2(n162), .ZN(\ab[19][22] ) );
  NOR2_X1 U1071 ( .A1(n250), .A2(n162), .ZN(\ab[19][21] ) );
  NOR2_X1 U1072 ( .A1(n253), .A2(n162), .ZN(\ab[19][20] ) );
  NOR2_X1 U1073 ( .A1(n310), .A2(n161), .ZN(\ab[19][1] ) );
  NOR2_X1 U1074 ( .A1(n256), .A2(n161), .ZN(\ab[19][19] ) );
  NOR2_X1 U1075 ( .A1(n259), .A2(n161), .ZN(\ab[19][18] ) );
  NOR2_X1 U1076 ( .A1(n262), .A2(n161), .ZN(\ab[19][17] ) );
  NOR2_X1 U1077 ( .A1(n265), .A2(n161), .ZN(\ab[19][16] ) );
  NOR2_X1 U1078 ( .A1(n268), .A2(n161), .ZN(\ab[19][15] ) );
  NOR2_X1 U1079 ( .A1(n271), .A2(n161), .ZN(\ab[19][14] ) );
  NOR2_X1 U1080 ( .A1(n274), .A2(n161), .ZN(\ab[19][13] ) );
  NOR2_X1 U1081 ( .A1(n277), .A2(n161), .ZN(\ab[19][12] ) );
  NOR2_X1 U1082 ( .A1(n280), .A2(n161), .ZN(\ab[19][11] ) );
  NOR2_X1 U1083 ( .A1(n283), .A2(n161), .ZN(\ab[19][10] ) );
  NOR2_X1 U1084 ( .A1(n313), .A2(n161), .ZN(\ab[19][0] ) );
  NOR2_X1 U1085 ( .A1(n286), .A2(n166), .ZN(\ab[18][9] ) );
  NOR2_X1 U1086 ( .A1(n289), .A2(n166), .ZN(\ab[18][8] ) );
  NOR2_X1 U1087 ( .A1(n292), .A2(n166), .ZN(\ab[18][7] ) );
  NOR2_X1 U1088 ( .A1(n295), .A2(n166), .ZN(\ab[18][6] ) );
  NOR2_X1 U1089 ( .A1(n298), .A2(n166), .ZN(\ab[18][5] ) );
  NOR2_X1 U1090 ( .A1(n301), .A2(n166), .ZN(\ab[18][4] ) );
  NOR2_X1 U1091 ( .A1(n304), .A2(n166), .ZN(\ab[18][3] ) );
  NOR2_X1 U1092 ( .A1(A[18]), .A2(n221), .ZN(\ab[18][31] ) );
  NOR2_X1 U1093 ( .A1(n223), .A2(n165), .ZN(\ab[18][30] ) );
  NOR2_X1 U1094 ( .A1(n307), .A2(n165), .ZN(\ab[18][2] ) );
  NOR2_X1 U1095 ( .A1(n226), .A2(n165), .ZN(\ab[18][29] ) );
  NOR2_X1 U1096 ( .A1(n229), .A2(n165), .ZN(\ab[18][28] ) );
  NOR2_X1 U1097 ( .A1(n232), .A2(n165), .ZN(\ab[18][27] ) );
  NOR2_X1 U1098 ( .A1(n235), .A2(n165), .ZN(\ab[18][26] ) );
  NOR2_X1 U1099 ( .A1(n238), .A2(n165), .ZN(\ab[18][25] ) );
  NOR2_X1 U1100 ( .A1(n241), .A2(n165), .ZN(\ab[18][24] ) );
  NOR2_X1 U1101 ( .A1(n244), .A2(n165), .ZN(\ab[18][23] ) );
  NOR2_X1 U1102 ( .A1(n247), .A2(n165), .ZN(\ab[18][22] ) );
  NOR2_X1 U1103 ( .A1(n250), .A2(n165), .ZN(\ab[18][21] ) );
  NOR2_X1 U1104 ( .A1(n253), .A2(n165), .ZN(\ab[18][20] ) );
  NOR2_X1 U1105 ( .A1(n310), .A2(n164), .ZN(\ab[18][1] ) );
  NOR2_X1 U1106 ( .A1(n256), .A2(n164), .ZN(\ab[18][19] ) );
  NOR2_X1 U1107 ( .A1(n259), .A2(n164), .ZN(\ab[18][18] ) );
  NOR2_X1 U1108 ( .A1(n262), .A2(n164), .ZN(\ab[18][17] ) );
  NOR2_X1 U1109 ( .A1(n265), .A2(n164), .ZN(\ab[18][16] ) );
  NOR2_X1 U1110 ( .A1(n268), .A2(n164), .ZN(\ab[18][15] ) );
  NOR2_X1 U1111 ( .A1(n271), .A2(n164), .ZN(\ab[18][14] ) );
  NOR2_X1 U1112 ( .A1(n274), .A2(n164), .ZN(\ab[18][13] ) );
  NOR2_X1 U1113 ( .A1(n277), .A2(n164), .ZN(\ab[18][12] ) );
  NOR2_X1 U1114 ( .A1(n280), .A2(n164), .ZN(\ab[18][11] ) );
  NOR2_X1 U1115 ( .A1(n283), .A2(n164), .ZN(\ab[18][10] ) );
  NOR2_X1 U1116 ( .A1(n313), .A2(n164), .ZN(\ab[18][0] ) );
  NOR2_X1 U1117 ( .A1(n286), .A2(n169), .ZN(\ab[17][9] ) );
  NOR2_X1 U1118 ( .A1(n289), .A2(n169), .ZN(\ab[17][8] ) );
  NOR2_X1 U1119 ( .A1(n292), .A2(n169), .ZN(\ab[17][7] ) );
  NOR2_X1 U1120 ( .A1(n295), .A2(n169), .ZN(\ab[17][6] ) );
  NOR2_X1 U1121 ( .A1(n298), .A2(n169), .ZN(\ab[17][5] ) );
  NOR2_X1 U1122 ( .A1(n301), .A2(n169), .ZN(\ab[17][4] ) );
  NOR2_X1 U1123 ( .A1(n304), .A2(n169), .ZN(\ab[17][3] ) );
  NOR2_X1 U1124 ( .A1(A[17]), .A2(n221), .ZN(\ab[17][31] ) );
  NOR2_X1 U1125 ( .A1(n223), .A2(n168), .ZN(\ab[17][30] ) );
  NOR2_X1 U1126 ( .A1(n307), .A2(n168), .ZN(\ab[17][2] ) );
  NOR2_X1 U1127 ( .A1(n226), .A2(n168), .ZN(\ab[17][29] ) );
  NOR2_X1 U1128 ( .A1(n229), .A2(n168), .ZN(\ab[17][28] ) );
  NOR2_X1 U1129 ( .A1(n232), .A2(n168), .ZN(\ab[17][27] ) );
  NOR2_X1 U1130 ( .A1(n235), .A2(n168), .ZN(\ab[17][26] ) );
  NOR2_X1 U1131 ( .A1(n238), .A2(n168), .ZN(\ab[17][25] ) );
  NOR2_X1 U1132 ( .A1(n241), .A2(n168), .ZN(\ab[17][24] ) );
  NOR2_X1 U1133 ( .A1(n244), .A2(n168), .ZN(\ab[17][23] ) );
  NOR2_X1 U1134 ( .A1(n247), .A2(n168), .ZN(\ab[17][22] ) );
  NOR2_X1 U1135 ( .A1(n250), .A2(n168), .ZN(\ab[17][21] ) );
  NOR2_X1 U1136 ( .A1(n253), .A2(n168), .ZN(\ab[17][20] ) );
  NOR2_X1 U1137 ( .A1(n310), .A2(n167), .ZN(\ab[17][1] ) );
  NOR2_X1 U1138 ( .A1(n256), .A2(n167), .ZN(\ab[17][19] ) );
  NOR2_X1 U1139 ( .A1(n259), .A2(n167), .ZN(\ab[17][18] ) );
  NOR2_X1 U1140 ( .A1(n262), .A2(n167), .ZN(\ab[17][17] ) );
  NOR2_X1 U1141 ( .A1(n265), .A2(n167), .ZN(\ab[17][16] ) );
  NOR2_X1 U1142 ( .A1(n268), .A2(n167), .ZN(\ab[17][15] ) );
  NOR2_X1 U1143 ( .A1(n271), .A2(n167), .ZN(\ab[17][14] ) );
  NOR2_X1 U1144 ( .A1(n274), .A2(n167), .ZN(\ab[17][13] ) );
  NOR2_X1 U1145 ( .A1(n277), .A2(n167), .ZN(\ab[17][12] ) );
  NOR2_X1 U1146 ( .A1(n280), .A2(n167), .ZN(\ab[17][11] ) );
  NOR2_X1 U1147 ( .A1(n283), .A2(n167), .ZN(\ab[17][10] ) );
  NOR2_X1 U1148 ( .A1(n313), .A2(n167), .ZN(\ab[17][0] ) );
  NOR2_X1 U1149 ( .A1(n286), .A2(n172), .ZN(\ab[16][9] ) );
  NOR2_X1 U1150 ( .A1(n289), .A2(n172), .ZN(\ab[16][8] ) );
  NOR2_X1 U1151 ( .A1(n292), .A2(n172), .ZN(\ab[16][7] ) );
  NOR2_X1 U1152 ( .A1(n295), .A2(n172), .ZN(\ab[16][6] ) );
  NOR2_X1 U1153 ( .A1(n298), .A2(n172), .ZN(\ab[16][5] ) );
  NOR2_X1 U1154 ( .A1(n301), .A2(n172), .ZN(\ab[16][4] ) );
  NOR2_X1 U1155 ( .A1(n304), .A2(n172), .ZN(\ab[16][3] ) );
  NOR2_X1 U1156 ( .A1(A[16]), .A2(n221), .ZN(\ab[16][31] ) );
  NOR2_X1 U1157 ( .A1(n223), .A2(n171), .ZN(\ab[16][30] ) );
  NOR2_X1 U1158 ( .A1(n307), .A2(n171), .ZN(\ab[16][2] ) );
  NOR2_X1 U1159 ( .A1(n226), .A2(n171), .ZN(\ab[16][29] ) );
  NOR2_X1 U1160 ( .A1(n229), .A2(n171), .ZN(\ab[16][28] ) );
  NOR2_X1 U1161 ( .A1(n232), .A2(n171), .ZN(\ab[16][27] ) );
  NOR2_X1 U1162 ( .A1(n235), .A2(n171), .ZN(\ab[16][26] ) );
  NOR2_X1 U1163 ( .A1(n238), .A2(n171), .ZN(\ab[16][25] ) );
  NOR2_X1 U1164 ( .A1(n241), .A2(n171), .ZN(\ab[16][24] ) );
  NOR2_X1 U1165 ( .A1(n244), .A2(n171), .ZN(\ab[16][23] ) );
  NOR2_X1 U1166 ( .A1(n247), .A2(n171), .ZN(\ab[16][22] ) );
  NOR2_X1 U1167 ( .A1(n250), .A2(n171), .ZN(\ab[16][21] ) );
  NOR2_X1 U1168 ( .A1(n253), .A2(n171), .ZN(\ab[16][20] ) );
  NOR2_X1 U1169 ( .A1(n310), .A2(n170), .ZN(\ab[16][1] ) );
  NOR2_X1 U1170 ( .A1(n256), .A2(n170), .ZN(\ab[16][19] ) );
  NOR2_X1 U1171 ( .A1(n259), .A2(n170), .ZN(\ab[16][18] ) );
  NOR2_X1 U1172 ( .A1(n262), .A2(n170), .ZN(\ab[16][17] ) );
  NOR2_X1 U1173 ( .A1(n265), .A2(n170), .ZN(\ab[16][16] ) );
  NOR2_X1 U1174 ( .A1(n268), .A2(n170), .ZN(\ab[16][15] ) );
  NOR2_X1 U1175 ( .A1(n271), .A2(n170), .ZN(\ab[16][14] ) );
  NOR2_X1 U1176 ( .A1(n274), .A2(n170), .ZN(\ab[16][13] ) );
  NOR2_X1 U1177 ( .A1(n277), .A2(n170), .ZN(\ab[16][12] ) );
  NOR2_X1 U1178 ( .A1(n280), .A2(n170), .ZN(\ab[16][11] ) );
  NOR2_X1 U1179 ( .A1(n283), .A2(n170), .ZN(\ab[16][10] ) );
  NOR2_X1 U1180 ( .A1(n313), .A2(n170), .ZN(\ab[16][0] ) );
  NOR2_X1 U1181 ( .A1(n286), .A2(n175), .ZN(\ab[15][9] ) );
  NOR2_X1 U1182 ( .A1(n289), .A2(n175), .ZN(\ab[15][8] ) );
  NOR2_X1 U1183 ( .A1(n292), .A2(n175), .ZN(\ab[15][7] ) );
  NOR2_X1 U1184 ( .A1(n295), .A2(n175), .ZN(\ab[15][6] ) );
  NOR2_X1 U1185 ( .A1(n298), .A2(n175), .ZN(\ab[15][5] ) );
  NOR2_X1 U1186 ( .A1(n301), .A2(n175), .ZN(\ab[15][4] ) );
  NOR2_X1 U1187 ( .A1(n304), .A2(n175), .ZN(\ab[15][3] ) );
  NOR2_X1 U1188 ( .A1(A[15]), .A2(n221), .ZN(\ab[15][31] ) );
  NOR2_X1 U1189 ( .A1(n223), .A2(n174), .ZN(\ab[15][30] ) );
  NOR2_X1 U1190 ( .A1(n307), .A2(n174), .ZN(\ab[15][2] ) );
  NOR2_X1 U1191 ( .A1(n226), .A2(n174), .ZN(\ab[15][29] ) );
  NOR2_X1 U1192 ( .A1(n229), .A2(n174), .ZN(\ab[15][28] ) );
  NOR2_X1 U1193 ( .A1(n232), .A2(n174), .ZN(\ab[15][27] ) );
  NOR2_X1 U1194 ( .A1(n235), .A2(n174), .ZN(\ab[15][26] ) );
  NOR2_X1 U1195 ( .A1(n238), .A2(n174), .ZN(\ab[15][25] ) );
  NOR2_X1 U1196 ( .A1(n241), .A2(n174), .ZN(\ab[15][24] ) );
  NOR2_X1 U1197 ( .A1(n244), .A2(n174), .ZN(\ab[15][23] ) );
  NOR2_X1 U1198 ( .A1(n247), .A2(n174), .ZN(\ab[15][22] ) );
  NOR2_X1 U1199 ( .A1(n250), .A2(n174), .ZN(\ab[15][21] ) );
  NOR2_X1 U1200 ( .A1(n253), .A2(n174), .ZN(\ab[15][20] ) );
  NOR2_X1 U1201 ( .A1(n310), .A2(n173), .ZN(\ab[15][1] ) );
  NOR2_X1 U1202 ( .A1(n256), .A2(n173), .ZN(\ab[15][19] ) );
  NOR2_X1 U1203 ( .A1(n259), .A2(n173), .ZN(\ab[15][18] ) );
  NOR2_X1 U1204 ( .A1(n262), .A2(n173), .ZN(\ab[15][17] ) );
  NOR2_X1 U1205 ( .A1(n265), .A2(n173), .ZN(\ab[15][16] ) );
  NOR2_X1 U1206 ( .A1(n268), .A2(n173), .ZN(\ab[15][15] ) );
  NOR2_X1 U1207 ( .A1(n271), .A2(n173), .ZN(\ab[15][14] ) );
  NOR2_X1 U1208 ( .A1(n274), .A2(n173), .ZN(\ab[15][13] ) );
  NOR2_X1 U1209 ( .A1(n277), .A2(n173), .ZN(\ab[15][12] ) );
  NOR2_X1 U1210 ( .A1(n280), .A2(n173), .ZN(\ab[15][11] ) );
  NOR2_X1 U1211 ( .A1(n283), .A2(n173), .ZN(\ab[15][10] ) );
  NOR2_X1 U1212 ( .A1(n313), .A2(n173), .ZN(\ab[15][0] ) );
  NOR2_X1 U1213 ( .A1(n286), .A2(n178), .ZN(\ab[14][9] ) );
  NOR2_X1 U1214 ( .A1(n289), .A2(n178), .ZN(\ab[14][8] ) );
  NOR2_X1 U1215 ( .A1(n292), .A2(n178), .ZN(\ab[14][7] ) );
  NOR2_X1 U1216 ( .A1(n295), .A2(n178), .ZN(\ab[14][6] ) );
  NOR2_X1 U1217 ( .A1(n298), .A2(n178), .ZN(\ab[14][5] ) );
  NOR2_X1 U1218 ( .A1(n301), .A2(n178), .ZN(\ab[14][4] ) );
  NOR2_X1 U1219 ( .A1(n304), .A2(n178), .ZN(\ab[14][3] ) );
  NOR2_X1 U1220 ( .A1(A[14]), .A2(n221), .ZN(\ab[14][31] ) );
  NOR2_X1 U1221 ( .A1(n223), .A2(n177), .ZN(\ab[14][30] ) );
  NOR2_X1 U1222 ( .A1(n307), .A2(n177), .ZN(\ab[14][2] ) );
  NOR2_X1 U1223 ( .A1(n226), .A2(n177), .ZN(\ab[14][29] ) );
  NOR2_X1 U1224 ( .A1(n229), .A2(n177), .ZN(\ab[14][28] ) );
  NOR2_X1 U1225 ( .A1(n232), .A2(n177), .ZN(\ab[14][27] ) );
  NOR2_X1 U1226 ( .A1(n235), .A2(n177), .ZN(\ab[14][26] ) );
  NOR2_X1 U1227 ( .A1(n238), .A2(n177), .ZN(\ab[14][25] ) );
  NOR2_X1 U1228 ( .A1(n241), .A2(n177), .ZN(\ab[14][24] ) );
  NOR2_X1 U1229 ( .A1(n244), .A2(n177), .ZN(\ab[14][23] ) );
  NOR2_X1 U1230 ( .A1(n247), .A2(n177), .ZN(\ab[14][22] ) );
  NOR2_X1 U1231 ( .A1(n250), .A2(n177), .ZN(\ab[14][21] ) );
  NOR2_X1 U1232 ( .A1(n253), .A2(n177), .ZN(\ab[14][20] ) );
  NOR2_X1 U1233 ( .A1(n310), .A2(n176), .ZN(\ab[14][1] ) );
  NOR2_X1 U1234 ( .A1(n256), .A2(n176), .ZN(\ab[14][19] ) );
  NOR2_X1 U1235 ( .A1(n259), .A2(n176), .ZN(\ab[14][18] ) );
  NOR2_X1 U1236 ( .A1(n262), .A2(n176), .ZN(\ab[14][17] ) );
  NOR2_X1 U1237 ( .A1(n265), .A2(n176), .ZN(\ab[14][16] ) );
  NOR2_X1 U1238 ( .A1(n268), .A2(n176), .ZN(\ab[14][15] ) );
  NOR2_X1 U1239 ( .A1(n271), .A2(n176), .ZN(\ab[14][14] ) );
  NOR2_X1 U1240 ( .A1(n274), .A2(n176), .ZN(\ab[14][13] ) );
  NOR2_X1 U1241 ( .A1(n277), .A2(n176), .ZN(\ab[14][12] ) );
  NOR2_X1 U1242 ( .A1(n280), .A2(n176), .ZN(\ab[14][11] ) );
  NOR2_X1 U1243 ( .A1(n283), .A2(n176), .ZN(\ab[14][10] ) );
  NOR2_X1 U1244 ( .A1(n313), .A2(n176), .ZN(\ab[14][0] ) );
  NOR2_X1 U1245 ( .A1(n286), .A2(n181), .ZN(\ab[13][9] ) );
  NOR2_X1 U1246 ( .A1(n289), .A2(n181), .ZN(\ab[13][8] ) );
  NOR2_X1 U1247 ( .A1(n292), .A2(n181), .ZN(\ab[13][7] ) );
  NOR2_X1 U1248 ( .A1(n295), .A2(n181), .ZN(\ab[13][6] ) );
  NOR2_X1 U1249 ( .A1(n298), .A2(n181), .ZN(\ab[13][5] ) );
  NOR2_X1 U1250 ( .A1(n301), .A2(n181), .ZN(\ab[13][4] ) );
  NOR2_X1 U1251 ( .A1(n304), .A2(n181), .ZN(\ab[13][3] ) );
  NOR2_X1 U1252 ( .A1(A[13]), .A2(n221), .ZN(\ab[13][31] ) );
  NOR2_X1 U1253 ( .A1(n223), .A2(n180), .ZN(\ab[13][30] ) );
  NOR2_X1 U1254 ( .A1(n307), .A2(n180), .ZN(\ab[13][2] ) );
  NOR2_X1 U1255 ( .A1(n226), .A2(n180), .ZN(\ab[13][29] ) );
  NOR2_X1 U1256 ( .A1(n229), .A2(n180), .ZN(\ab[13][28] ) );
  NOR2_X1 U1257 ( .A1(n232), .A2(n180), .ZN(\ab[13][27] ) );
  NOR2_X1 U1258 ( .A1(n235), .A2(n180), .ZN(\ab[13][26] ) );
  NOR2_X1 U1259 ( .A1(n238), .A2(n180), .ZN(\ab[13][25] ) );
  NOR2_X1 U1260 ( .A1(n241), .A2(n180), .ZN(\ab[13][24] ) );
  NOR2_X1 U1261 ( .A1(n244), .A2(n180), .ZN(\ab[13][23] ) );
  NOR2_X1 U1262 ( .A1(n247), .A2(n180), .ZN(\ab[13][22] ) );
  NOR2_X1 U1263 ( .A1(n250), .A2(n180), .ZN(\ab[13][21] ) );
  NOR2_X1 U1264 ( .A1(n253), .A2(n180), .ZN(\ab[13][20] ) );
  NOR2_X1 U1265 ( .A1(n310), .A2(n179), .ZN(\ab[13][1] ) );
  NOR2_X1 U1266 ( .A1(n256), .A2(n179), .ZN(\ab[13][19] ) );
  NOR2_X1 U1267 ( .A1(n259), .A2(n179), .ZN(\ab[13][18] ) );
  NOR2_X1 U1268 ( .A1(n262), .A2(n179), .ZN(\ab[13][17] ) );
  NOR2_X1 U1269 ( .A1(n265), .A2(n179), .ZN(\ab[13][16] ) );
  NOR2_X1 U1270 ( .A1(n268), .A2(n179), .ZN(\ab[13][15] ) );
  NOR2_X1 U1271 ( .A1(n271), .A2(n179), .ZN(\ab[13][14] ) );
  NOR2_X1 U1272 ( .A1(n274), .A2(n179), .ZN(\ab[13][13] ) );
  NOR2_X1 U1273 ( .A1(n277), .A2(n179), .ZN(\ab[13][12] ) );
  NOR2_X1 U1274 ( .A1(n280), .A2(n179), .ZN(\ab[13][11] ) );
  NOR2_X1 U1275 ( .A1(n283), .A2(n179), .ZN(\ab[13][10] ) );
  NOR2_X1 U1276 ( .A1(n313), .A2(n179), .ZN(\ab[13][0] ) );
  NOR2_X1 U1277 ( .A1(n286), .A2(n184), .ZN(\ab[12][9] ) );
  NOR2_X1 U1278 ( .A1(n289), .A2(n184), .ZN(\ab[12][8] ) );
  NOR2_X1 U1279 ( .A1(n292), .A2(n184), .ZN(\ab[12][7] ) );
  NOR2_X1 U1280 ( .A1(n295), .A2(n184), .ZN(\ab[12][6] ) );
  NOR2_X1 U1281 ( .A1(n298), .A2(n184), .ZN(\ab[12][5] ) );
  NOR2_X1 U1282 ( .A1(n301), .A2(n184), .ZN(\ab[12][4] ) );
  NOR2_X1 U1283 ( .A1(n304), .A2(n184), .ZN(\ab[12][3] ) );
  NOR2_X1 U1284 ( .A1(A[12]), .A2(n221), .ZN(\ab[12][31] ) );
  NOR2_X1 U1285 ( .A1(n223), .A2(n183), .ZN(\ab[12][30] ) );
  NOR2_X1 U1286 ( .A1(n307), .A2(n183), .ZN(\ab[12][2] ) );
  NOR2_X1 U1287 ( .A1(n226), .A2(n183), .ZN(\ab[12][29] ) );
  NOR2_X1 U1288 ( .A1(n229), .A2(n183), .ZN(\ab[12][28] ) );
  NOR2_X1 U1289 ( .A1(n232), .A2(n183), .ZN(\ab[12][27] ) );
  NOR2_X1 U1290 ( .A1(n235), .A2(n183), .ZN(\ab[12][26] ) );
  NOR2_X1 U1291 ( .A1(n238), .A2(n183), .ZN(\ab[12][25] ) );
  NOR2_X1 U1292 ( .A1(n241), .A2(n183), .ZN(\ab[12][24] ) );
  NOR2_X1 U1293 ( .A1(n244), .A2(n183), .ZN(\ab[12][23] ) );
  NOR2_X1 U1294 ( .A1(n247), .A2(n183), .ZN(\ab[12][22] ) );
  NOR2_X1 U1295 ( .A1(n250), .A2(n183), .ZN(\ab[12][21] ) );
  NOR2_X1 U1296 ( .A1(n253), .A2(n183), .ZN(\ab[12][20] ) );
  NOR2_X1 U1297 ( .A1(n310), .A2(n182), .ZN(\ab[12][1] ) );
  NOR2_X1 U1298 ( .A1(n256), .A2(n182), .ZN(\ab[12][19] ) );
  NOR2_X1 U1299 ( .A1(n259), .A2(n182), .ZN(\ab[12][18] ) );
  NOR2_X1 U1300 ( .A1(n262), .A2(n182), .ZN(\ab[12][17] ) );
  NOR2_X1 U1301 ( .A1(n265), .A2(n182), .ZN(\ab[12][16] ) );
  NOR2_X1 U1302 ( .A1(n268), .A2(n182), .ZN(\ab[12][15] ) );
  NOR2_X1 U1303 ( .A1(n271), .A2(n182), .ZN(\ab[12][14] ) );
  NOR2_X1 U1304 ( .A1(n274), .A2(n182), .ZN(\ab[12][13] ) );
  NOR2_X1 U1305 ( .A1(n277), .A2(n182), .ZN(\ab[12][12] ) );
  NOR2_X1 U1306 ( .A1(n280), .A2(n182), .ZN(\ab[12][11] ) );
  NOR2_X1 U1307 ( .A1(n283), .A2(n182), .ZN(\ab[12][10] ) );
  NOR2_X1 U1308 ( .A1(n313), .A2(n182), .ZN(\ab[12][0] ) );
  NOR2_X1 U1309 ( .A1(n286), .A2(n187), .ZN(\ab[11][9] ) );
  NOR2_X1 U1310 ( .A1(n289), .A2(n187), .ZN(\ab[11][8] ) );
  NOR2_X1 U1311 ( .A1(n292), .A2(n187), .ZN(\ab[11][7] ) );
  NOR2_X1 U1312 ( .A1(n295), .A2(n187), .ZN(\ab[11][6] ) );
  NOR2_X1 U1313 ( .A1(n298), .A2(n187), .ZN(\ab[11][5] ) );
  NOR2_X1 U1314 ( .A1(n301), .A2(n187), .ZN(\ab[11][4] ) );
  NOR2_X1 U1315 ( .A1(n304), .A2(n187), .ZN(\ab[11][3] ) );
  NOR2_X1 U1316 ( .A1(A[11]), .A2(n221), .ZN(\ab[11][31] ) );
  NOR2_X1 U1317 ( .A1(n223), .A2(n186), .ZN(\ab[11][30] ) );
  NOR2_X1 U1318 ( .A1(n307), .A2(n186), .ZN(\ab[11][2] ) );
  NOR2_X1 U1319 ( .A1(n226), .A2(n186), .ZN(\ab[11][29] ) );
  NOR2_X1 U1320 ( .A1(n229), .A2(n186), .ZN(\ab[11][28] ) );
  NOR2_X1 U1321 ( .A1(n232), .A2(n186), .ZN(\ab[11][27] ) );
  NOR2_X1 U1322 ( .A1(n235), .A2(n186), .ZN(\ab[11][26] ) );
  NOR2_X1 U1323 ( .A1(n238), .A2(n186), .ZN(\ab[11][25] ) );
  NOR2_X1 U1324 ( .A1(n241), .A2(n186), .ZN(\ab[11][24] ) );
  NOR2_X1 U1325 ( .A1(n244), .A2(n186), .ZN(\ab[11][23] ) );
  NOR2_X1 U1326 ( .A1(n247), .A2(n186), .ZN(\ab[11][22] ) );
  NOR2_X1 U1327 ( .A1(n250), .A2(n186), .ZN(\ab[11][21] ) );
  NOR2_X1 U1328 ( .A1(n253), .A2(n186), .ZN(\ab[11][20] ) );
  NOR2_X1 U1329 ( .A1(n310), .A2(n185), .ZN(\ab[11][1] ) );
  NOR2_X1 U1330 ( .A1(n256), .A2(n185), .ZN(\ab[11][19] ) );
  NOR2_X1 U1331 ( .A1(n259), .A2(n185), .ZN(\ab[11][18] ) );
  NOR2_X1 U1332 ( .A1(n262), .A2(n185), .ZN(\ab[11][17] ) );
  NOR2_X1 U1333 ( .A1(n265), .A2(n185), .ZN(\ab[11][16] ) );
  NOR2_X1 U1334 ( .A1(n268), .A2(n185), .ZN(\ab[11][15] ) );
  NOR2_X1 U1335 ( .A1(n271), .A2(n185), .ZN(\ab[11][14] ) );
  NOR2_X1 U1336 ( .A1(n274), .A2(n185), .ZN(\ab[11][13] ) );
  NOR2_X1 U1337 ( .A1(n277), .A2(n185), .ZN(\ab[11][12] ) );
  NOR2_X1 U1338 ( .A1(n280), .A2(n185), .ZN(\ab[11][11] ) );
  NOR2_X1 U1339 ( .A1(n283), .A2(n185), .ZN(\ab[11][10] ) );
  NOR2_X1 U1340 ( .A1(n313), .A2(n185), .ZN(\ab[11][0] ) );
  NOR2_X1 U1341 ( .A1(n286), .A2(n190), .ZN(\ab[10][9] ) );
  NOR2_X1 U1342 ( .A1(n289), .A2(n190), .ZN(\ab[10][8] ) );
  NOR2_X1 U1343 ( .A1(n292), .A2(n190), .ZN(\ab[10][7] ) );
  NOR2_X1 U1344 ( .A1(n295), .A2(n190), .ZN(\ab[10][6] ) );
  NOR2_X1 U1345 ( .A1(n298), .A2(n190), .ZN(\ab[10][5] ) );
  NOR2_X1 U1346 ( .A1(n301), .A2(n190), .ZN(\ab[10][4] ) );
  NOR2_X1 U1347 ( .A1(n304), .A2(n190), .ZN(\ab[10][3] ) );
  NOR2_X1 U1348 ( .A1(A[10]), .A2(n221), .ZN(\ab[10][31] ) );
  NOR2_X1 U1349 ( .A1(n223), .A2(n189), .ZN(\ab[10][30] ) );
  NOR2_X1 U1350 ( .A1(n307), .A2(n189), .ZN(\ab[10][2] ) );
  NOR2_X1 U1351 ( .A1(n226), .A2(n189), .ZN(\ab[10][29] ) );
  NOR2_X1 U1352 ( .A1(n229), .A2(n189), .ZN(\ab[10][28] ) );
  NOR2_X1 U1353 ( .A1(n232), .A2(n189), .ZN(\ab[10][27] ) );
  NOR2_X1 U1354 ( .A1(n235), .A2(n189), .ZN(\ab[10][26] ) );
  NOR2_X1 U1355 ( .A1(n238), .A2(n189), .ZN(\ab[10][25] ) );
  NOR2_X1 U1356 ( .A1(n241), .A2(n189), .ZN(\ab[10][24] ) );
  NOR2_X1 U1357 ( .A1(n244), .A2(n189), .ZN(\ab[10][23] ) );
  NOR2_X1 U1358 ( .A1(n247), .A2(n189), .ZN(\ab[10][22] ) );
  NOR2_X1 U1359 ( .A1(n250), .A2(n189), .ZN(\ab[10][21] ) );
  NOR2_X1 U1360 ( .A1(n253), .A2(n189), .ZN(\ab[10][20] ) );
  NOR2_X1 U1361 ( .A1(n310), .A2(n188), .ZN(\ab[10][1] ) );
  NOR2_X1 U1362 ( .A1(n256), .A2(n188), .ZN(\ab[10][19] ) );
  NOR2_X1 U1363 ( .A1(n259), .A2(n188), .ZN(\ab[10][18] ) );
  NOR2_X1 U1364 ( .A1(n262), .A2(n188), .ZN(\ab[10][17] ) );
  NOR2_X1 U1365 ( .A1(n265), .A2(n188), .ZN(\ab[10][16] ) );
  NOR2_X1 U1366 ( .A1(n268), .A2(n188), .ZN(\ab[10][15] ) );
  NOR2_X1 U1367 ( .A1(n271), .A2(n188), .ZN(\ab[10][14] ) );
  NOR2_X1 U1368 ( .A1(n274), .A2(n188), .ZN(\ab[10][13] ) );
  NOR2_X1 U1369 ( .A1(n277), .A2(n188), .ZN(\ab[10][12] ) );
  NOR2_X1 U1370 ( .A1(n280), .A2(n188), .ZN(\ab[10][11] ) );
  NOR2_X1 U1371 ( .A1(n283), .A2(n188), .ZN(\ab[10][10] ) );
  NOR2_X1 U1372 ( .A1(n313), .A2(n188), .ZN(\ab[10][0] ) );
  NOR2_X1 U1373 ( .A1(n286), .A2(n220), .ZN(\ab[0][9] ) );
  NOR2_X1 U1374 ( .A1(n289), .A2(n220), .ZN(\ab[0][8] ) );
  NOR2_X1 U1375 ( .A1(n292), .A2(n220), .ZN(\ab[0][7] ) );
  NOR2_X1 U1376 ( .A1(n295), .A2(n220), .ZN(\ab[0][6] ) );
  NOR2_X1 U1377 ( .A1(n298), .A2(n220), .ZN(\ab[0][5] ) );
  NOR2_X1 U1378 ( .A1(n301), .A2(n220), .ZN(\ab[0][4] ) );
  NOR2_X1 U1379 ( .A1(n304), .A2(n220), .ZN(\ab[0][3] ) );
  NOR2_X1 U1380 ( .A1(A[0]), .A2(n221), .ZN(\ab[0][31] ) );
  NOR2_X1 U1381 ( .A1(n223), .A2(n219), .ZN(\ab[0][30] ) );
  NOR2_X1 U1382 ( .A1(n307), .A2(n219), .ZN(\ab[0][2] ) );
  NOR2_X1 U1383 ( .A1(n226), .A2(n219), .ZN(\ab[0][29] ) );
  NOR2_X1 U1384 ( .A1(n229), .A2(n219), .ZN(\ab[0][28] ) );
  NOR2_X1 U1385 ( .A1(n232), .A2(n219), .ZN(\ab[0][27] ) );
  NOR2_X1 U1386 ( .A1(n235), .A2(n219), .ZN(\ab[0][26] ) );
  NOR2_X1 U1387 ( .A1(n238), .A2(n219), .ZN(\ab[0][25] ) );
  NOR2_X1 U1388 ( .A1(n241), .A2(n219), .ZN(\ab[0][24] ) );
  NOR2_X1 U1389 ( .A1(n244), .A2(n219), .ZN(\ab[0][23] ) );
  NOR2_X1 U1390 ( .A1(n247), .A2(n219), .ZN(\ab[0][22] ) );
  NOR2_X1 U1391 ( .A1(n250), .A2(n219), .ZN(\ab[0][21] ) );
  NOR2_X1 U1392 ( .A1(n253), .A2(n219), .ZN(\ab[0][20] ) );
  NOR2_X1 U1393 ( .A1(n310), .A2(n218), .ZN(\ab[0][1] ) );
  NOR2_X1 U1394 ( .A1(n256), .A2(n218), .ZN(\ab[0][19] ) );
  NOR2_X1 U1395 ( .A1(n259), .A2(n218), .ZN(\ab[0][18] ) );
  NOR2_X1 U1396 ( .A1(n262), .A2(n218), .ZN(\ab[0][17] ) );
  NOR2_X1 U1397 ( .A1(n265), .A2(n218), .ZN(\ab[0][16] ) );
  NOR2_X1 U1398 ( .A1(n268), .A2(n218), .ZN(\ab[0][15] ) );
  NOR2_X1 U1399 ( .A1(n271), .A2(n218), .ZN(\ab[0][14] ) );
  NOR2_X1 U1400 ( .A1(n274), .A2(n218), .ZN(\ab[0][13] ) );
  NOR2_X1 U1401 ( .A1(n277), .A2(n218), .ZN(\ab[0][12] ) );
  NOR2_X1 U1402 ( .A1(n280), .A2(n218), .ZN(\ab[0][11] ) );
  NOR2_X1 U1403 ( .A1(n283), .A2(n218), .ZN(\ab[0][10] ) );
  NOR2_X1 U1404 ( .A1(n313), .A2(n218), .ZN(PRODUCT[0]) );
endmodule


module VerilogMultiplier ( clk, rst, A, B, P );
  input [31:0] A;
  input [31:0] B;
  output [63:0] P;
  input clk, rst;
  wire   N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13;
  wire   [31:0] B_reg;
  wire   [31:0] A_reg;

  DFFR_X1 \A_reg_reg[31]  ( .D(A[31]), .CK(clk), .RN(n12), .Q(A_reg[31]) );
  DFFR_X1 \A_reg_reg[30]  ( .D(A[30]), .CK(clk), .RN(n12), .Q(A_reg[30]) );
  DFFR_X1 \A_reg_reg[29]  ( .D(A[29]), .CK(clk), .RN(n12), .Q(A_reg[29]) );
  DFFR_X1 \A_reg_reg[28]  ( .D(A[28]), .CK(clk), .RN(n12), .Q(A_reg[28]) );
  DFFR_X1 \A_reg_reg[27]  ( .D(A[27]), .CK(clk), .RN(n12), .Q(A_reg[27]) );
  DFFR_X1 \A_reg_reg[26]  ( .D(A[26]), .CK(clk), .RN(n12), .Q(A_reg[26]) );
  DFFR_X1 \A_reg_reg[25]  ( .D(A[25]), .CK(clk), .RN(n12), .Q(A_reg[25]) );
  DFFR_X1 \A_reg_reg[24]  ( .D(A[24]), .CK(clk), .RN(n12), .Q(A_reg[24]) );
  DFFR_X1 \A_reg_reg[23]  ( .D(A[23]), .CK(clk), .RN(n11), .Q(A_reg[23]) );
  DFFR_X1 \A_reg_reg[22]  ( .D(A[22]), .CK(clk), .RN(n11), .Q(A_reg[22]) );
  DFFR_X1 \A_reg_reg[21]  ( .D(A[21]), .CK(clk), .RN(n11), .Q(A_reg[21]) );
  DFFR_X1 \A_reg_reg[20]  ( .D(A[20]), .CK(clk), .RN(n11), .Q(A_reg[20]) );
  DFFR_X1 \A_reg_reg[19]  ( .D(A[19]), .CK(clk), .RN(n11), .Q(A_reg[19]) );
  DFFR_X1 \A_reg_reg[18]  ( .D(A[18]), .CK(clk), .RN(n11), .Q(A_reg[18]) );
  DFFR_X1 \A_reg_reg[17]  ( .D(A[17]), .CK(clk), .RN(n11), .Q(A_reg[17]) );
  DFFR_X1 \A_reg_reg[16]  ( .D(A[16]), .CK(clk), .RN(n11), .Q(A_reg[16]) );
  DFFR_X1 \A_reg_reg[15]  ( .D(A[15]), .CK(clk), .RN(n11), .Q(A_reg[15]) );
  DFFR_X1 \A_reg_reg[14]  ( .D(A[14]), .CK(clk), .RN(n11), .Q(A_reg[14]) );
  DFFR_X1 \A_reg_reg[13]  ( .D(A[13]), .CK(clk), .RN(n11), .Q(A_reg[13]) );
  DFFR_X1 \A_reg_reg[12]  ( .D(A[12]), .CK(clk), .RN(n11), .Q(A_reg[12]) );
  DFFR_X1 \A_reg_reg[11]  ( .D(A[11]), .CK(clk), .RN(n10), .Q(A_reg[11]) );
  DFFR_X1 \A_reg_reg[10]  ( .D(A[10]), .CK(clk), .RN(n10), .Q(A_reg[10]) );
  DFFR_X1 \A_reg_reg[9]  ( .D(A[9]), .CK(clk), .RN(n10), .Q(A_reg[9]) );
  DFFR_X1 \A_reg_reg[8]  ( .D(A[8]), .CK(clk), .RN(n10), .Q(A_reg[8]) );
  DFFR_X1 \A_reg_reg[7]  ( .D(A[7]), .CK(clk), .RN(n10), .Q(A_reg[7]) );
  DFFR_X1 \A_reg_reg[6]  ( .D(A[6]), .CK(clk), .RN(n10), .Q(A_reg[6]) );
  DFFR_X1 \A_reg_reg[5]  ( .D(A[5]), .CK(clk), .RN(n10), .Q(A_reg[5]) );
  DFFR_X1 \A_reg_reg[4]  ( .D(A[4]), .CK(clk), .RN(n10), .Q(A_reg[4]) );
  DFFR_X1 \A_reg_reg[3]  ( .D(A[3]), .CK(clk), .RN(n10), .Q(A_reg[3]) );
  DFFR_X1 \A_reg_reg[2]  ( .D(A[2]), .CK(clk), .RN(n10), .Q(A_reg[2]) );
  DFFR_X1 \A_reg_reg[1]  ( .D(A[1]), .CK(clk), .RN(n10), .Q(A_reg[1]) );
  DFFR_X1 \A_reg_reg[0]  ( .D(A[0]), .CK(clk), .RN(n10), .Q(A_reg[0]) );
  DFFR_X1 \P_reg_reg[63]  ( .D(N64), .CK(clk), .RN(n9), .Q(P[63]) );
  DFFR_X1 \P_reg_reg[62]  ( .D(N63), .CK(clk), .RN(n9), .Q(P[62]) );
  DFFR_X1 \P_reg_reg[61]  ( .D(N62), .CK(clk), .RN(n9), .Q(P[61]) );
  DFFR_X1 \P_reg_reg[60]  ( .D(N61), .CK(clk), .RN(n9), .Q(P[60]) );
  DFFR_X1 \P_reg_reg[59]  ( .D(N60), .CK(clk), .RN(n9), .Q(P[59]) );
  DFFR_X1 \P_reg_reg[58]  ( .D(N59), .CK(clk), .RN(n9), .Q(P[58]) );
  DFFR_X1 \P_reg_reg[57]  ( .D(N58), .CK(clk), .RN(n9), .Q(P[57]) );
  DFFR_X1 \P_reg_reg[56]  ( .D(N57), .CK(clk), .RN(n9), .Q(P[56]) );
  DFFR_X1 \P_reg_reg[55]  ( .D(N56), .CK(clk), .RN(n9), .Q(P[55]) );
  DFFR_X1 \P_reg_reg[54]  ( .D(N55), .CK(clk), .RN(n9), .Q(P[54]) );
  DFFR_X1 \P_reg_reg[53]  ( .D(N54), .CK(clk), .RN(n9), .Q(P[53]) );
  DFFR_X1 \P_reg_reg[52]  ( .D(N53), .CK(clk), .RN(n9), .Q(P[52]) );
  DFFR_X1 \P_reg_reg[51]  ( .D(N52), .CK(clk), .RN(n8), .Q(P[51]) );
  DFFR_X1 \P_reg_reg[50]  ( .D(N51), .CK(clk), .RN(n8), .Q(P[50]) );
  DFFR_X1 \P_reg_reg[49]  ( .D(N50), .CK(clk), .RN(n8), .Q(P[49]) );
  DFFR_X1 \P_reg_reg[48]  ( .D(N49), .CK(clk), .RN(n8), .Q(P[48]) );
  DFFR_X1 \P_reg_reg[47]  ( .D(N48), .CK(clk), .RN(n8), .Q(P[47]) );
  DFFR_X1 \P_reg_reg[46]  ( .D(N47), .CK(clk), .RN(n8), .Q(P[46]) );
  DFFR_X1 \P_reg_reg[45]  ( .D(N46), .CK(clk), .RN(n8), .Q(P[45]) );
  DFFR_X1 \P_reg_reg[44]  ( .D(N45), .CK(clk), .RN(n8), .Q(P[44]) );
  DFFR_X1 \P_reg_reg[43]  ( .D(N44), .CK(clk), .RN(n8), .Q(P[43]) );
  DFFR_X1 \P_reg_reg[42]  ( .D(N43), .CK(clk), .RN(n8), .Q(P[42]) );
  DFFR_X1 \P_reg_reg[41]  ( .D(N42), .CK(clk), .RN(n8), .Q(P[41]) );
  DFFR_X1 \P_reg_reg[40]  ( .D(N41), .CK(clk), .RN(n8), .Q(P[40]) );
  DFFR_X1 \P_reg_reg[39]  ( .D(N40), .CK(clk), .RN(n7), .Q(P[39]) );
  DFFR_X1 \P_reg_reg[38]  ( .D(N39), .CK(clk), .RN(n7), .Q(P[38]) );
  DFFR_X1 \P_reg_reg[37]  ( .D(N38), .CK(clk), .RN(n7), .Q(P[37]) );
  DFFR_X1 \P_reg_reg[36]  ( .D(N37), .CK(clk), .RN(n7), .Q(P[36]) );
  DFFR_X1 \P_reg_reg[35]  ( .D(N36), .CK(clk), .RN(n7), .Q(P[35]) );
  DFFR_X1 \P_reg_reg[34]  ( .D(N35), .CK(clk), .RN(n7), .Q(P[34]) );
  DFFR_X1 \P_reg_reg[33]  ( .D(N34), .CK(clk), .RN(n7), .Q(P[33]) );
  DFFR_X1 \P_reg_reg[32]  ( .D(N33), .CK(clk), .RN(n7), .Q(P[32]) );
  DFFR_X1 \P_reg_reg[31]  ( .D(N32), .CK(clk), .RN(n7), .Q(P[31]) );
  DFFR_X1 \P_reg_reg[30]  ( .D(N31), .CK(clk), .RN(n7), .Q(P[30]) );
  DFFR_X1 \P_reg_reg[29]  ( .D(N30), .CK(clk), .RN(n7), .Q(P[29]) );
  DFFR_X1 \P_reg_reg[28]  ( .D(N29), .CK(clk), .RN(n7), .Q(P[28]) );
  DFFR_X1 \P_reg_reg[27]  ( .D(N28), .CK(clk), .RN(n6), .Q(P[27]) );
  DFFR_X1 \P_reg_reg[26]  ( .D(N27), .CK(clk), .RN(n6), .Q(P[26]) );
  DFFR_X1 \P_reg_reg[25]  ( .D(N26), .CK(clk), .RN(n6), .Q(P[25]) );
  DFFR_X1 \P_reg_reg[24]  ( .D(N25), .CK(clk), .RN(n6), .Q(P[24]) );
  DFFR_X1 \P_reg_reg[23]  ( .D(N24), .CK(clk), .RN(n6), .Q(P[23]) );
  DFFR_X1 \P_reg_reg[22]  ( .D(N23), .CK(clk), .RN(n6), .Q(P[22]) );
  DFFR_X1 \P_reg_reg[21]  ( .D(N22), .CK(clk), .RN(n6), .Q(P[21]) );
  DFFR_X1 \P_reg_reg[20]  ( .D(N21), .CK(clk), .RN(n6), .Q(P[20]) );
  DFFR_X1 \P_reg_reg[19]  ( .D(N20), .CK(clk), .RN(n6), .Q(P[19]) );
  DFFR_X1 \P_reg_reg[18]  ( .D(N19), .CK(clk), .RN(n6), .Q(P[18]) );
  DFFR_X1 \P_reg_reg[17]  ( .D(N18), .CK(clk), .RN(n6), .Q(P[17]) );
  DFFR_X1 \P_reg_reg[16]  ( .D(N17), .CK(clk), .RN(n6), .Q(P[16]) );
  DFFR_X1 \P_reg_reg[15]  ( .D(N16), .CK(clk), .RN(n5), .Q(P[15]) );
  DFFR_X1 \P_reg_reg[14]  ( .D(N15), .CK(clk), .RN(n5), .Q(P[14]) );
  DFFR_X1 \P_reg_reg[13]  ( .D(N14), .CK(clk), .RN(n5), .Q(P[13]) );
  DFFR_X1 \P_reg_reg[12]  ( .D(N13), .CK(clk), .RN(n5), .Q(P[12]) );
  DFFR_X1 \P_reg_reg[11]  ( .D(N12), .CK(clk), .RN(n5), .Q(P[11]) );
  DFFR_X1 \P_reg_reg[10]  ( .D(N11), .CK(clk), .RN(n5), .Q(P[10]) );
  DFFR_X1 \P_reg_reg[9]  ( .D(N10), .CK(clk), .RN(n5), .Q(P[9]) );
  DFFR_X1 \P_reg_reg[8]  ( .D(N9), .CK(clk), .RN(n5), .Q(P[8]) );
  DFFR_X1 \P_reg_reg[7]  ( .D(N8), .CK(clk), .RN(n5), .Q(P[7]) );
  DFFR_X1 \P_reg_reg[6]  ( .D(N7), .CK(clk), .RN(n5), .Q(P[6]) );
  DFFR_X1 \P_reg_reg[5]  ( .D(N6), .CK(clk), .RN(n5), .Q(P[5]) );
  DFFR_X1 \P_reg_reg[4]  ( .D(N5), .CK(clk), .RN(n5), .Q(P[4]) );
  DFFR_X1 \P_reg_reg[3]  ( .D(N4), .CK(clk), .RN(n4), .Q(P[3]) );
  DFFR_X1 \P_reg_reg[2]  ( .D(N3), .CK(clk), .RN(n4), .Q(P[2]) );
  DFFR_X1 \P_reg_reg[1]  ( .D(N2), .CK(clk), .RN(n4), .Q(P[1]) );
  DFFR_X1 \P_reg_reg[0]  ( .D(N1), .CK(clk), .RN(n4), .Q(P[0]) );
  DFFR_X1 \B_reg_reg[31]  ( .D(B[31]), .CK(clk), .RN(n4), .Q(B_reg[31]) );
  DFFR_X1 \B_reg_reg[30]  ( .D(B[30]), .CK(clk), .RN(n4), .Q(B_reg[30]) );
  DFFR_X1 \B_reg_reg[29]  ( .D(B[29]), .CK(clk), .RN(n4), .Q(B_reg[29]) );
  DFFR_X1 \B_reg_reg[28]  ( .D(B[28]), .CK(clk), .RN(n4), .Q(B_reg[28]) );
  DFFR_X1 \B_reg_reg[27]  ( .D(B[27]), .CK(clk), .RN(n4), .Q(B_reg[27]) );
  DFFR_X1 \B_reg_reg[26]  ( .D(B[26]), .CK(clk), .RN(n4), .Q(B_reg[26]) );
  DFFR_X1 \B_reg_reg[25]  ( .D(B[25]), .CK(clk), .RN(n4), .Q(B_reg[25]) );
  DFFR_X1 \B_reg_reg[24]  ( .D(B[24]), .CK(clk), .RN(n4), .Q(B_reg[24]) );
  DFFR_X1 \B_reg_reg[23]  ( .D(B[23]), .CK(clk), .RN(n3), .Q(B_reg[23]) );
  DFFR_X1 \B_reg_reg[22]  ( .D(B[22]), .CK(clk), .RN(n3), .Q(B_reg[22]) );
  DFFR_X1 \B_reg_reg[21]  ( .D(B[21]), .CK(clk), .RN(n3), .Q(B_reg[21]) );
  DFFR_X1 \B_reg_reg[20]  ( .D(B[20]), .CK(clk), .RN(n3), .Q(B_reg[20]) );
  DFFR_X1 \B_reg_reg[19]  ( .D(B[19]), .CK(clk), .RN(n3), .Q(B_reg[19]) );
  DFFR_X1 \B_reg_reg[18]  ( .D(B[18]), .CK(clk), .RN(n3), .Q(B_reg[18]) );
  DFFR_X1 \B_reg_reg[17]  ( .D(B[17]), .CK(clk), .RN(n3), .Q(B_reg[17]) );
  DFFR_X1 \B_reg_reg[16]  ( .D(B[16]), .CK(clk), .RN(n3), .Q(B_reg[16]) );
  DFFR_X1 \B_reg_reg[15]  ( .D(B[15]), .CK(clk), .RN(n3), .Q(B_reg[15]) );
  DFFR_X1 \B_reg_reg[14]  ( .D(B[14]), .CK(clk), .RN(n3), .Q(B_reg[14]) );
  DFFR_X1 \B_reg_reg[13]  ( .D(B[13]), .CK(clk), .RN(n3), .Q(B_reg[13]) );
  DFFR_X1 \B_reg_reg[12]  ( .D(B[12]), .CK(clk), .RN(n3), .Q(B_reg[12]) );
  DFFR_X1 \B_reg_reg[11]  ( .D(B[11]), .CK(clk), .RN(n2), .Q(B_reg[11]) );
  DFFR_X1 \B_reg_reg[10]  ( .D(B[10]), .CK(clk), .RN(n2), .Q(B_reg[10]) );
  DFFR_X1 \B_reg_reg[9]  ( .D(B[9]), .CK(clk), .RN(n2), .Q(B_reg[9]) );
  DFFR_X1 \B_reg_reg[8]  ( .D(B[8]), .CK(clk), .RN(n2), .Q(B_reg[8]) );
  DFFR_X1 \B_reg_reg[7]  ( .D(B[7]), .CK(clk), .RN(n2), .Q(B_reg[7]) );
  DFFR_X1 \B_reg_reg[6]  ( .D(B[6]), .CK(clk), .RN(n2), .Q(B_reg[6]) );
  DFFR_X1 \B_reg_reg[5]  ( .D(B[5]), .CK(clk), .RN(n2), .Q(B_reg[5]) );
  DFFR_X1 \B_reg_reg[4]  ( .D(B[4]), .CK(clk), .RN(n2), .Q(B_reg[4]) );
  DFFR_X1 \B_reg_reg[3]  ( .D(B[3]), .CK(clk), .RN(n2), .Q(B_reg[3]) );
  DFFR_X1 \B_reg_reg[2]  ( .D(B[2]), .CK(clk), .RN(n2), .Q(B_reg[2]) );
  DFFR_X1 \B_reg_reg[1]  ( .D(B[1]), .CK(clk), .RN(n2), .Q(B_reg[1]) );
  DFFR_X1 \B_reg_reg[0]  ( .D(B[0]), .CK(clk), .RN(n2), .Q(B_reg[0]) );
  VerilogMultiplier_DW02_mult_0 mult_21 ( .A(A_reg), .B(B_reg), .TC(1'b1), 
        .PRODUCT({N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  INV_X1 U4 ( .A(rst), .ZN(n13) );
  BUF_X1 U5 ( .A(n13), .Z(n2) );
  BUF_X1 U6 ( .A(n13), .Z(n3) );
  BUF_X1 U7 ( .A(n13), .Z(n4) );
  BUF_X1 U8 ( .A(n13), .Z(n5) );
  BUF_X1 U9 ( .A(n13), .Z(n6) );
  BUF_X1 U10 ( .A(n13), .Z(n7) );
  BUF_X1 U11 ( .A(n13), .Z(n8) );
  BUF_X1 U12 ( .A(n13), .Z(n9) );
  BUF_X1 U13 ( .A(n13), .Z(n10) );
  BUF_X1 U14 ( .A(n13), .Z(n11) );
  BUF_X1 U15 ( .A(n13), .Z(n12) );
endmodule

