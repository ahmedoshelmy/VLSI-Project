
module BoothMultiplier_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n13, n15, n16, n17, n19, n21,
         n23, n27, n28, n29, n30, n32, n33, n35, n36, n39, n40, n42, n43, n44,
         n46, n47, n48, n50, n53, n54, n55, n56, n57, n58, n59, n61, n62, n65,
         n66, n68, n69, n71, n72, n74, n75, n76, n78, n79, n81, n84, n86, n90,
         n91, n94, n95, n96, n97, n99, n100, n101, n103, n104, n105, n106,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n119,
         n120, n121, n122, n123, n124, n126, n127, n128, n129, n130, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n147, n148, n151, n154, n155, n156, n157, n158, n159, n160, n164,
         n165, n166, n169, n170, n171, n172, n175, n176, n177, n178, n181,
         n182, n183, n186, n187, n188, n189, n191, n194, n195, n196, n197,
         n199, n200, n201, n202, n203, n204, n205, n207, n208, n209, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n222, n226, n227,
         n229, n230, n231, n232, n233, n234, n235, n236, n238, n241, n242,
         n243, n244, n245, n247, n248, n251, n252, n253, n254, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n270, n271,
         n272, n273, n274, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n289, n290, n291, n292, n293, n294, n295, n298,
         n301, n302, n305, n306, n308, n311, n312, n313, n315, n316, n317,
         n319, n320, n321, n322, n323, n325, n327, n328, n329, n330, n331,
         n333, n334, n335, n336, n338, n339, n341, n342, n344, n345, n346,
         n350, n351, n353, n357, n358, n361, n362, n364, n365, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491;

  NAND4X0 U3 ( .IN1(n262), .IN2(n260), .IN3(n261), .IN4(n259), .QN(n55) );
  AND2X1 U8 ( .IN1(n175), .IN2(n176), .Q(n3) );
  XOR3X1 U9 ( .IN1(n467), .IN2(B[29]), .IN3(n57), .Q(DIFF[29]) );
  AND2X1 U10 ( .IN1(n422), .IN2(n207), .Q(n1) );
  AND2X1 U11 ( .IN1(n272), .IN2(n305), .Q(n2) );
  AND2X1 U12 ( .IN1(n169), .IN2(n170), .Q(n4) );
  AND2X1 U17 ( .IN1(n8), .IN2(n9), .Q(n301) );
  OR2X1 U18 ( .IN1(n435), .IN2(n272), .Q(n9) );
  OR2X1 U23 ( .IN1(n395), .IN2(n148), .Q(n13) );
  AND2X1 U25 ( .IN1(n158), .IN2(n147), .Q(n15) );
  XOR3X1 U26 ( .IN1(n466), .IN2(B[30]), .IN3(n144), .Q(DIFF[30]) );
  OR2X1 U30 ( .IN1(n402), .IN2(n165), .Q(n17) );
  AND2X1 U32 ( .IN1(n169), .IN2(n164), .Q(n19) );
  AND2X1 U36 ( .IN1(n186), .IN2(n181), .Q(n23) );
  AND2X1 U40 ( .IN1(n1), .IN2(n202), .Q(n27) );
  AND2X1 U43 ( .IN1(n61), .IN2(n44), .Q(n28) );
  AND2X1 U46 ( .IN1(n46), .IN2(n76), .Q(n30) );
  XOR3X1 U49 ( .IN1(A[31]), .IN2(n392), .IN3(n140), .Q(DIFF[31]) );
  AND2X1 U56 ( .IN1(n205), .IN2(n72), .Q(n35) );
  AND2X1 U60 ( .IN1(n42), .IN2(n66), .Q(n39) );
  OR2X1 U64 ( .IN1(n397), .IN2(n48), .Q(n44) );
  AND2X1 U66 ( .IN1(n50), .IN2(n158), .Q(n46) );
  AND2X1 U71 ( .IN1(n53), .IN2(n79), .Q(n50) );
  AND2X1 U74 ( .IN1(n175), .IN2(n69), .Q(n53) );
  AND2X1 U76 ( .IN1(n134), .IN2(n338), .Q(n56) );
  AND2X1 U81 ( .IN1(n58), .IN2(n59), .Q(n142) );
  OR2X1 U82 ( .IN1(n394), .IN2(n147), .Q(n59) );
  AND2X1 U84 ( .IN1(n148), .IN2(n143), .Q(n61) );
  OR2X1 U85 ( .IN1(n410), .IN2(n200), .Q(n62) );
  OR2X1 U89 ( .IN1(n409), .IN2(n194), .Q(n66) );
  AND2X1 U91 ( .IN1(n197), .IN2(n74), .Q(n68) );
  OR2X1 U92 ( .IN1(n401), .IN2(n169), .Q(n69) );
  AND2X1 U94 ( .IN1(n171), .IN2(n81), .Q(n71) );
  OR2X1 U95 ( .IN1(n407), .IN2(n186), .Q(n72) );
  AND2X1 U97 ( .IN1(n189), .IN2(n78), .Q(n74) );
  AND2X1 U98 ( .IN1(n75), .IN2(n76), .Q(n176) );
  OR2X1 U99 ( .IN1(n406), .IN2(n181), .Q(n76) );
  AND2X1 U101 ( .IN1(n182), .IN2(n177), .Q(n78) );
  OR2X1 U102 ( .IN1(n399), .IN2(n164), .Q(n79) );
  AND2X1 U104 ( .IN1(n165), .IN2(n160), .Q(n81) );
  AND2X1 U156 ( .IN1(n219), .IN2(n207), .Q(n99) );
  AND2X1 U184 ( .IN1(n278), .IN2(n320), .Q(n84) );
  AND2X1 U190 ( .IN1(n112), .IN2(n113), .Q(n86) );
  OR2X1 U199 ( .IN1(n439), .IN2(A[12]), .Q(n294) );
  OR2X1 U204 ( .IN1(n450), .IN2(A[6]), .Q(n117) );
  NAND3X0 U209 ( .IN1(A[0]), .IN2(n157), .IN3(n139), .QN(n345) );
  OR2X1 U214 ( .IN1(n441), .IN2(A[11]), .Q(n278) );
  OR2X1 U225 ( .IN1(n418), .IN2(A[21]), .Q(n202) );
  OR2X1 U226 ( .IN1(n415), .IN2(A[22]), .Q(n197) );
  AND2X1 U265 ( .IN1(n279), .IN2(n94), .Q(n263) );
  OR2X1 U270 ( .IN1(n464), .IN2(A[0]), .Q(n229) );
  OR2X1 U284 ( .IN1(n420), .IN2(n217), .Q(n97) );
  XOR2X1 U375 ( .IN1(n101), .IN2(n446), .Q(DIFF[9]) );
  XOR2X1 U376 ( .IN1(n106), .IN2(n448), .Q(DIFF[8]) );
  XOR2X1 U377 ( .IN1(n111), .IN2(n86), .Q(DIFF[7]) );
  XOR2X1 U378 ( .IN1(n451), .IN2(n119), .Q(DIFF[6]) );
  XOR2X1 U379 ( .IN1(n124), .IN2(n453), .Q(DIFF[5]) );
  XOR2X1 U380 ( .IN1(n130), .IN2(n455), .Q(DIFF[4]) );
  XOR2X1 U382 ( .IN1(n138), .IN2(n151), .Q(DIFF[2]) );
  XOR2X1 U383 ( .IN1(n4), .IN2(n166), .Q(DIFF[27]) );
  XOR2X1 U384 ( .IN1(n3), .IN2(n172), .Q(DIFF[26]) );
  XOR2X1 U385 ( .IN1(n7), .IN2(n178), .Q(DIFF[25]) );
  XOR2X1 U386 ( .IN1(n5), .IN2(n183), .Q(DIFF[24]) );
  XOR2X1 U387 ( .IN1(n414), .IN2(n191), .Q(DIFF[23]) );
  XOR2X1 U388 ( .IN1(n416), .IN2(n199), .Q(DIFF[22]) );
  XOR2X1 U389 ( .IN1(n203), .IN2(n6), .Q(DIFF[21]) );
  XOR2X1 U390 ( .IN1(n213), .IN2(n214), .Q(DIFF[20]) );
  XOR2X1 U391 ( .IN1(n463), .IN2(n226), .Q(DIFF[1]) );
  XOR2X1 U392 ( .IN1(n230), .IN2(n231), .Q(DIFF[19]) );
  XOR2X1 U393 ( .IN1(n241), .IN2(n242), .Q(DIFF[18]) );
  XOR2X1 U394 ( .IN1(n251), .IN2(n252), .Q(DIFF[17]) );
  XOR2X1 U395 ( .IN1(n258), .IN2(n430), .Q(DIFF[16]) );
  NAND4X0 U396 ( .IN1(n262), .IN2(n260), .IN3(n261), .IN4(n259), .QN(n208) );
  XOR2X1 U399 ( .IN1(n2), .IN2(n302), .Q(DIFF[14]) );
  XOR2X1 U400 ( .IN1(n437), .IN2(n308), .Q(DIFF[13]) );
  XOR2X1 U401 ( .IN1(n313), .IN2(n440), .Q(DIFF[12]) );
  NAND3X0 U402 ( .IN1(n321), .IN2(n320), .IN3(n319), .QN(n279) );
  NAND4X0 U403 ( .IN1(A[8]), .IN2(n325), .IN3(n104), .IN4(n447), .QN(n319) );
  XOR2X1 U404 ( .IN1(n327), .IN2(n84), .Q(DIFF[11]) );
  XOR2X1 U405 ( .IN1(n331), .IN2(n444), .Q(DIFF[10]) );
  NAND4X0 U406 ( .IN1(A[4]), .IN2(n117), .IN3(n123), .IN4(n454), .QN(n362) );
  INVX0 U4 ( (n66), (n408) );
  INVX0 U5 ( (n55), (n430) );
  NOR2X0 U6 ( .IN1(n430), .IN2(n222), .QN(n232) );
  NOR2X0 U7 ( .IN1(n430), .IN2(n238), .QN(n243) );
  AND2X1 U13 ( .IN1(n204), .IN2(n62), .Q(n42) );
  AND2X1 U14 ( .IN1(n54), .IN2(n204), .Q(n6) );
  INVX0 U15 ( (n116), (n451) );
  INVX0 U16 ( (n188), (n414) );
  INVX0 U19 ( (n196), (n416) );
  INVX0 U20 ( (n330), (n444) );
  INVX0 U21 ( (n129), (n455) );
  INVX0 U22 ( (n103), (n446) );
  NAND2X1 U24 ( .IN1(n72), .IN2(n373), .QN(n33) );
  NOR2X0 U27 ( .IN1(n408), .IN2(n40), .QN(n373) );
  INVX0 U28 ( (n122), (n453) );
  INVX0 U29 ( (n277), (n438) );
  INVX0 U31 ( (n69), (n400) );
  INVX0 U33 ( (n156), (n463) );
  NAND2X1 U34 ( .IN1(n122), .IN2(n123), .QN(n121) );
  NOR2X0 U35 ( .IN1(n215), .IN2(n212), .QN(n214) );
  NAND2X1 U37 ( .IN1(n216), .IN2(n217), .QN(n212) );
  AND2X1 U38 ( .IN1(n374), .IN2(n211), .Q(n204) );
  AND2X1 U39 ( .IN1(n96), .IN2(n97), .Q(n374) );
  NAND2X1 U41 ( .IN1(n100), .IN2(n112), .QN(n335) );
  NAND2X1 U42 ( .IN1(n104), .IN2(n103), .QN(n333) );
  NAND2X1 U44 ( .IN1(n285), .IN2(n112), .QN(n282) );
  NOR2X0 U45 ( .IN1(n456), .IN2(n344), .QN(n342) );
  NOR2X0 U47 ( .IN1(n458), .IN2(n136), .QN(n351) );
  NAND2X1 U48 ( .IN1(n279), .IN2(n278), .QN(n315) );
  INVX0 U50 ( (n164), (n402) );
  NOR2X0 U51 ( .IN1(n375), .IN2(n376), .QN(n201) );
  AND2X1 U52 ( .IN1(n55), .IN2(n27), .Q(n375) );
  NOR2X0 U53 ( .IN1(n417), .IN2(n204), .QN(n376) );
  OR2X1 U54 ( .IN1(n291), .IN2(n377), .Q(n129) );
  AND2X1 U55 ( .IN1(n134), .IN2(n338), .Q(n377) );
  NOR2X0 U57 ( .IN1(n378), .IN2(n379), .QN(n7) );
  AND2X1 U58 ( .IN1(n188), .IN2(n391), .Q(n378) );
  NOR2X0 U59 ( .IN1(n390), .IN2(n23), .QN(n379) );
  NAND2X1 U61 ( .IN1(n110), .IN2(n334), .QN(n103) );
  NAND2X1 U62 ( .IN1(n154), .IN2(n155), .QN(n138) );
  NAND2X1 U63 ( .IN1(n126), .IN2(n127), .QN(n122) );
  NAND2X1 U65 ( .IN1(A[12]), .IN2(n439), .QN(n277) );
  NOR2X0 U67 ( .IN1(n154), .IN2(n353), .QN(n350) );
  INVX0 U68 ( (n254), (n427) );
  NAND2X1 U69 ( .IN1(n426), .IN2(n236), .QN(n222) );
  INVX0 U70 ( (n134), (n458) );
  NOR2X0 U72 ( .IN1(n253), .IN2(n427), .QN(n252) );
  NOR2X0 U73 ( .IN1(n429), .IN2(n430), .QN(n253) );
  INVX0 U75 ( (n248), (n429) );
  NOR2X0 U77 ( .IN1(n357), .IN2(n358), .QN(n289) );
  NAND2X1 U78 ( .IN1(n128), .IN2(n123), .QN(n357) );
  NAND2X1 U79 ( .IN1(n112), .IN2(n117), .QN(n358) );
  NOR2X0 U80 ( .IN1(n459), .IN2(n461), .QN(n151) );
  XNOR2X1 U83 ( .IN1(n133), .IN2(n380), .Q(DIFF[3]) );
  NAND2X1 U86 ( .IN1(n134), .IN2(n135), .QN(n380) );
  NAND2X1 U87 ( .IN1(n128), .IN2(n126), .QN(n130) );
  NAND2X1 U88 ( .IN1(n169), .IN2(n171), .QN(n172) );
  NAND2X1 U90 ( .IN1(n164), .IN2(n165), .QN(n166) );
  NAND2X1 U93 ( .IN1(n202), .IN2(n200), .QN(n203) );
  NAND2X1 U96 ( .IN1(n109), .IN2(n110), .QN(n106) );
  XNOR2X1 U100 ( .IN1(n298), .IN2(n381), .Q(DIFF[15]) );
  NAND2X1 U103 ( .IN1(n271), .IN2(n260), .QN(n381) );
  NAND2X1 U105 ( .IN1(n294), .IN2(n277), .QN(n313) );
  NAND2X1 U106 ( .IN1(n248), .IN2(n254), .QN(n258) );
  NOR2X0 U107 ( .IN1(n267), .IN2(n268), .QN(n266) );
  NOR2X0 U108 ( .IN1(n432), .IN2(n270), .QN(n268) );
  NAND2X1 U109 ( .IN1(n114), .IN2(n115), .QN(n111) );
  NAND2X1 U110 ( .IN1(n116), .IN2(n117), .QN(n114) );
  NAND2X1 U111 ( .IN1(n227), .IN2(n465), .QN(n156) );
  INVX0 U112 ( (n95), (n465) );
  INVX0 U113 ( (n81), (n401) );
  INVX0 U114 ( (n74), (n409) );
  INVX0 U115 ( (n135), (n456) );
  INVX0 U116 ( (n271), (n432) );
  NAND2X1 U117 ( .IN1(A[11]), .IN2(n441), .QN(n320) );
  NAND2X1 U118 ( .IN1(n270), .IN2(n301), .QN(n298) );
  NAND2X1 U119 ( .IN1(n136), .IN2(n137), .QN(n133) );
  NAND2X1 U120 ( .IN1(n138), .IN2(n139), .QN(n137) );
  INVX0 U121 ( (n207), (n420) );
  INVX0 U122 ( (n202), (n417) );
  NAND2X1 U123 ( .IN1(n79), .IN2(n382), .QN(n48) );
  NOR2X0 U124 ( .IN1(n400), .IN2(n71), .QN(n382) );
  NAND2X1 U125 ( .IN1(n62), .IN2(n383), .QN(n40) );
  NAND2X1 U126 ( .IN1(n202), .IN2(n68), .QN(n383) );
  INVX0 U127 ( (n160), (n399) );
  INVX0 U128 ( (n158), (n397) );
  NAND2X1 U129 ( .IN1(A[4]), .IN2(n454), .QN(n126) );
  NAND2X1 U130 ( .IN1(A[8]), .IN2(n447), .QN(n110) );
  AND2X1 U131 ( .IN1(n295), .IN2(n274), .Q(n11) );
  AND2X1 U132 ( .IN1(n189), .IN2(n21), .Q(n391) );
  OR2X1 U133 ( .IN1(n411), .IN2(n182), .Q(n21) );
  INVX0 U134 ( (n181), (n411) );
  NAND2X1 U135 ( .IN1(n115), .IN2(n117), .QN(n119) );
  INVX0 U136 ( (n136), (n459) );
  NAND2X1 U137 ( .IN1(n219), .IN2(n217), .QN(n230) );
  NAND2X1 U138 ( .IN1(n236), .IN2(n234), .QN(n241) );
  NAND2X1 U139 ( .IN1(n186), .IN2(n189), .QN(n191) );
  NAND2X1 U140 ( .IN1(n272), .IN2(n295), .QN(n308) );
  NAND2X1 U141 ( .IN1(n104), .IN2(n105), .QN(n101) );
  NAND2X1 U142 ( .IN1(n207), .IN2(n211), .QN(n213) );
  NAND2X1 U143 ( .IN1(n194), .IN2(n197), .QN(n199) );
  INVX0 U144 ( (n147), (n395) );
  INVX0 U145 ( (n274), (n435) );
  INVX0 U146 ( (n143), (n394) );
  INVX0 U147 ( (B[25]), (n405) );
  NOR2X0 U148 ( .IN1(B[10]), .IN2(n482), .QN(n323) );
  INVX0 U149 ( (B[5]), (n452) );
  INVX0 U150 ( (A[16]), (n478) );
  NOR2X0 U151 ( .IN1(n450), .IN2(A[6]), .QN(n36) );
  INVX0 U152 ( (B[7]), (n449) );
  INVX0 U153 ( (B[16]), (n428) );
  NAND2X1 U154 ( .IN1(A[30]), .IN2(n393), .QN(n141) );
  INVX0 U155 ( (B[30]), (n393) );
  NAND2X1 U157 ( .IN1(B[7]), .IN2(n485), .QN(n112) );
  INVX0 U158 ( (A[7]), (n485) );
  NAND2X1 U159 ( .IN1(B[5]), .IN2(n486), .QN(n123) );
  NOR2X0 U160 ( .IN1(n90), .IN2(n91), .QN(n284) );
  NAND2X1 U161 ( .IN1(n317), .IN2(n278), .QN(n91) );
  NAND2X1 U162 ( .IN1(B[10]), .IN2(n482), .QN(n317) );
  NAND2X1 U163 ( .IN1(B[9]), .IN2(n483), .QN(n104) );
  NAND2X1 U164 ( .IN1(A[6]), .IN2(n450), .QN(n115) );
  INVX0 U165 ( (A[10]), (n482) );
  NAND2X1 U166 ( .IN1(A[14]), .IN2(n434), .QN(n270) );
  INVX0 U167 ( (B[14]), (n434) );
  NAND2X1 U168 ( .IN1(A[2]), .IN2(n460), .QN(n136) );
  INVX0 U169 ( (B[2]), (n460) );
  NAND2X1 U170 ( .IN1(A[19]), .IN2(n421), .QN(n217) );
  INVX0 U171 ( (B[19]), (n421) );
  NAND2X1 U172 ( .IN1(A[27]), .IN2(n403), .QN(n164) );
  INVX0 U173 ( (B[27]), (n403) );
  NAND2X1 U174 ( .IN1(B[4]), .IN2(n487), .QN(n128) );
  INVX0 U175 ( (A[4]), (n487) );
  NAND2X1 U176 ( .IN1(B[19]), .IN2(n475), .QN(n219) );
  INVX0 U177 ( (A[19]), (n475) );
  NAND2X1 U178 ( .IN1(B[18]), .IN2(n476), .QN(n236) );
  INVX0 U179 ( (A[18]), (n476) );
  NAND2X1 U180 ( .IN1(A[1]), .IN2(n462), .QN(n154) );
  INVX0 U181 ( (B[1]), (n462) );
  NAND2X1 U182 ( .IN1(A[23]), .IN2(n413), .QN(n186) );
  INVX0 U183 ( (B[23]), (n413) );
  NAND2X1 U185 ( .IN1(A[26]), .IN2(n404), .QN(n169) );
  INVX0 U186 ( (B[26]), (n404) );
  NAND2X1 U187 ( .IN1(A[21]), .IN2(n418), .QN(n200) );
  NAND2X1 U188 ( .IN1(B[20]), .IN2(n474), .QN(n207) );
  INVX0 U189 ( (A[20]), (n474) );
  NAND2X1 U191 ( .IN1(A[13]), .IN2(n436), .QN(n272) );
  INVX0 U192 ( (B[13]), (n436) );
  NAND2X1 U193 ( .IN1(B[14]), .IN2(n480), .QN(n274) );
  INVX0 U194 ( (A[14]), (n480) );
  NAND2X1 U195 ( .IN1(B[27]), .IN2(n469), .QN(n165) );
  NAND2X1 U196 ( .IN1(B[8]), .IN2(n484), .QN(n109) );
  NAND2X1 U197 ( .IN1(B[23]), .IN2(n473), .QN(n189) );
  INVX0 U198 ( (A[23]), (n473) );
  NAND2X1 U200 ( .IN1(A[22]), .IN2(n415), .QN(n194) );
  NAND2X1 U201 ( .IN1(B[13]), .IN2(n481), .QN(n295) );
  INVX0 U202 ( (A[13]), (n481) );
  NAND2X1 U203 ( .IN1(B[0]), .IN2(n491), .QN(n95) );
  INVX0 U205 ( (A[0]), (n491) );
  NAND2X1 U206 ( .IN1(A[9]), .IN2(n445), .QN(n105) );
  INVX0 U207 ( (B[9]), (n445) );
  NAND2X1 U208 ( .IN1(A[18]), .IN2(n423), .QN(n234) );
  INVX0 U210 ( (B[18]), (n423) );
  NAND2X1 U211 ( .IN1(B[26]), .IN2(n470), .QN(n171) );
  INVX0 U212 ( (A[26]), (n470) );
  NAND2X1 U213 ( .IN1(A[20]), .IN2(n419), .QN(n211) );
  INVX0 U215 ( (B[20]), (n419) );
  NAND2X1 U216 ( .IN1(B[15]), .IN2(n479), .QN(n271) );
  INVX0 U217 ( (A[15]), (n479) );
  NAND2X1 U218 ( .IN1(n95), .IN2(n227), .QN(DIFF[0]) );
  NAND2X1 U219 ( .IN1(A[3]), .IN2(n457), .QN(n135) );
  INVX0 U220 ( (B[3]), (n457) );
  NAND2X1 U221 ( .IN1(B[28]), .IN2(n468), .QN(n160) );
  INVX0 U222 ( (A[28]), (n468) );
  NAND2X1 U223 ( .IN1(A[15]), .IN2(n431), .QN(n260) );
  INVX0 U224 ( (B[15]), (n431) );
  NAND2X0 U227 ( .IN1(B[17]), .IN2(n477), .QN(n247) );
  INVX0 U228 ( (A[17]), (n477) );
  NAND2X1 U229 ( .IN1(A[17]), .IN2(n425), .QN(n245) );
  INVX0 U230 ( (B[17]), (n425) );
  INVX0 U231 ( (B[24]), (n412) );
  INVX0 U232 ( (B[10]), (n442) );
  INVX0 U233 ( (A[29]), (n467) );
  INVX0 U234 ( (A[30]), (n466) );
  NAND2X1 U235 ( .IN1(A[0]), .IN2(n464), .QN(n227) );
  NAND2X1 U236 ( .IN1(A[28]), .IN2(n398), .QN(n158) );
  INVX0 U237 ( (B[28]), (n398) );
  NAND2X1 U238 ( .IN1(A[29]), .IN2(n396), .QN(n147) );
  INVX0 U239 ( (B[29]), (n396) );
  NAND2X1 U240 ( .IN1(B[30]), .IN2(n466), .QN(n143) );
  NAND2X1 U241 ( .IN1(B[29]), .IN2(n467), .QN(n148) );
  INVX0 U242 ( (B[6]), (n450) );
  INVX0 U243 ( (B[0]), (n464) );
  INVX0 U244 ( (B[8]), (n447) );
  INVX0 U245 ( (B[4]), (n454) );
  INVX0 U246 ( (B[21]), (n418) );
  INVX0 U247 ( (B[11]), (n441) );
  INVX0 U248 ( (B[22]), (n415) );
  INVX0 U249 ( (B[12]), (n439) );
  INVX0 U250 ( (B[31]), (n392) );
  NAND2X0 U251 ( .IN1(n233), .IN2(n234), .QN(n384) );
  INVX0 U252 ( (A[27]), (n469) );
  NAND2X1 U253 ( .IN1(n311), .IN2(n277), .QN(n306) );
  INVX0 U254 ( (n68), (n410) );
  NOR2X0 U255 ( .IN1(n430), .IN2(n209), .QN(n215) );
  INVX0 U256 ( (n209), (n422) );
  INVX0 U257 ( (n177), (n406) );
  INVX0 U258 ( (n78), (n407) );
  NAND2X0 U259 ( .IN1(B[25]), .IN2(n471), .QN(n177) );
  INVX0 U260 ( (n312), (n440) );
  INVX0 U261 ( (n108), (n448) );
  NAND2X0 U262 ( .IN1(n181), .IN2(n182), .QN(n183) );
  NAND2X1 U263 ( .IN1(n47), .IN2(n388), .QN(n385) );
  NAND2X0 U264 ( .IN1(n385), .IN2(n386), .QN(n144) );
  OR2X1 U266 ( .IN1(n387), .IN2(n15), .Q(n386) );
  INVX0 U267 ( (n13), (n387) );
  AND2X1 U268 ( .IN1(n48), .IN2(n13), .Q(n388) );
  NOR2X0 U269 ( .IN1(n243), .IN2(n235), .QN(n242) );
  NAND2X0 U271 ( .IN1(n233), .IN2(n234), .QN(n218) );
  NAND2X1 U272 ( .IN1(A[16]), .IN2(n428), .QN(n254) );
  NOR2X0 U273 ( .IN1(n263), .IN2(n264), .QN(n262) );
  INVX0 U274 ( (n238), (n426) );
  NAND2X0 U275 ( .IN1(n200), .IN2(n201), .QN(n196) );
  NAND2X0 U276 ( .IN1(n175), .IN2(n177), .QN(n178) );
  XOR3X1 U277 ( .IN1(A[28]), .IN2(B[28]), .IN3(n389), .Q(DIFF[28]) );
  NAND2X0 U278 ( .IN1(n16), .IN2(n17), .QN(n389) );
  NAND2X0 U279 ( .IN1(n123), .IN2(n120), .QN(n124) );
  NAND2X0 U280 ( .IN1(n120), .IN2(n121), .QN(n116) );
  NAND2X0 U281 ( .IN1(n361), .IN2(n362), .QN(n100) );
  NAND2X1 U282 ( .IN1(n361), .IN2(n362), .QN(n285) );
  NOR2X0 U283 ( .IN1(n339), .IN2(n461), .QN(n338) );
  INVX0 U285 ( (n139), (n461) );
  NAND4X0 U286 ( .IN1(n294), .IN2(n295), .IN3(n274), .IN4(n271), .QN(n290) );
  NAND2X0 U287 ( .IN1(n156), .IN2(n157), .QN(n155) );
  NAND2X0 U288 ( .IN1(n154), .IN2(n157), .QN(n226) );
  NAND2X0 U289 ( .IN1(n157), .IN2(n229), .QN(n339) );
  NAND2X0 U290 ( .IN1(n265), .IN2(n266), .QN(n264) );
  NAND2X0 U291 ( .IN1(n244), .IN2(n245), .QN(n235) );
  NOR2X0 U292 ( .IN1(n350), .IN2(n351), .QN(n341) );
  NAND2X0 U293 ( .IN1(n341), .IN2(n342), .QN(n291) );
  NAND2X0 U294 ( .IN1(A[25]), .IN2(n405), .QN(n175) );
  NOR2X0 U295 ( .IN1(n272), .IN2(n273), .QN(n267) );
  NAND2X0 U296 ( .IN1(n109), .IN2(n104), .QN(n90) );
  NOR2X0 U297 ( .IN1(n282), .IN2(n283), .QN(n281) );
  INVX0 U298 ( (A[9]), (n483) );
  INVX0 U299 ( (A[24]), (n472) );
  NAND2X1 U300 ( .IN1(B[24]), .IN2(n472), .QN(n182) );
  NAND2X0 U301 ( .IN1(A[24]), .IN2(n412), .QN(n181) );
  NAND2X0 U302 ( .IN1(n139), .IN2(n134), .QN(n353) );
  NAND2X0 U303 ( .IN1(n105), .IN2(n333), .QN(n330) );
  NAND2X0 U304 ( .IN1(n335), .IN2(n336), .QN(n108) );
  NAND2X0 U305 ( .IN1(n141), .IN2(n142), .QN(n140) );
  INVX0 U306 ( (A[25]), (n471) );
  NAND2X1 U307 ( .IN1(n424), .IN2(n219), .QN(n209) );
  INVX0 U308 ( (n222), (n424) );
  NAND2X1 U309 ( .IN1(B[16]), .IN2(n478), .QN(n248) );
  NAND2X0 U310 ( .IN1(n196), .IN2(n197), .QN(n195) );
  AND2X1 U311 ( .IN1(n433), .IN2(n278), .Q(n94) );
  INVX0 U312 ( (n290), (n433) );
  NAND2X0 U313 ( .IN1(n194), .IN2(n195), .QN(n188) );
  INVX0 U314 ( (n325), (n443) );
  NOR2X0 U315 ( .IN1(n443), .IN2(n105), .QN(n322) );
  NOR2X0 U316 ( .IN1(n322), .IN2(n323), .QN(n321) );
  NAND2X0 U317 ( .IN1(B[10]), .IN2(n482), .QN(n325) );
  NAND2X0 U318 ( .IN1(n284), .IN2(n56), .QN(n287) );
  NAND2X1 U319 ( .IN1(B[1]), .IN2(n490), .QN(n157) );
  INVX0 U320 ( (A[1]), (n490) );
  NAND2X0 U321 ( .IN1(n270), .IN2(n274), .QN(n302) );
  NOR2X0 U322 ( .IN1(n293), .IN2(n290), .QN(n292) );
  NAND2X0 U323 ( .IN1(n284), .IN2(n433), .QN(n283) );
  NAND2X0 U324 ( .IN1(n438), .IN2(n433), .QN(n265) );
  NAND2X0 U325 ( .IN1(n274), .IN2(n271), .QN(n273) );
  NAND2X0 U326 ( .IN1(n109), .IN2(n108), .QN(n334) );
  NAND2X0 U327 ( .IN1(n128), .IN2(n129), .QN(n127) );
  NOR2X0 U328 ( .IN1(n345), .IN2(n346), .QN(n344) );
  NAND2X0 U329 ( .IN1(n170), .IN2(n19), .QN(n16) );
  NAND2X0 U330 ( .IN1(n325), .IN2(n328), .QN(n331) );
  NAND2X0 U331 ( .IN1(n158), .IN2(n159), .QN(n57) );
  NAND2X0 U332 ( .IN1(A[10]), .IN2(n442), .QN(n328) );
  NAND2X0 U333 ( .IN1(n47), .IN2(n48), .QN(n159) );
  INVX0 U334 ( (A[5]), (n486) );
  NAND2X0 U335 ( .IN1(A[5]), .IN2(n452), .QN(n120) );
  INVX0 U336 ( (n21), (n390) );
  NAND2X0 U337 ( .IN1(n43), .IN2(n28), .QN(n58) );
  AND2X1 U338 ( .IN1(n186), .IN2(n187), .Q(n5) );
  NAND2X0 U339 ( .IN1(n188), .IN2(n189), .QN(n187) );
  NOR2X0 U340 ( .IN1(n280), .IN2(n281), .QN(n261) );
  NOR2X0 U341 ( .IN1(n365), .IN2(n364), .QN(n361) );
  NOR2X0 U342 ( .IN1(n36), .IN2(n120), .QN(n365) );
  NAND2X1 U343 ( .IN1(n113), .IN2(n115), .QN(n364) );
  INVX0 U344 ( (n306), (n437) );
  NAND2X0 U345 ( .IN1(n306), .IN2(n11), .QN(n8) );
  NAND2X0 U346 ( .IN1(n306), .IN2(n295), .QN(n305) );
  NAND2X1 U347 ( .IN1(B[2]), .IN2(n489), .QN(n139) );
  INVX0 U348 ( (A[2]), (n489) );
  NAND2X0 U349 ( .IN1(n330), .IN2(n325), .QN(n329) );
  NAND2X0 U350 ( .IN1(n65), .IN2(n171), .QN(n170) );
  NAND2X0 U351 ( .IN1(n175), .IN2(n176), .QN(n65) );
  NAND2X0 U352 ( .IN1(n291), .IN2(n292), .QN(n259) );
  NAND2X0 U353 ( .IN1(n433), .IN2(n289), .QN(n286) );
  NAND2X0 U354 ( .IN1(n284), .IN2(n289), .QN(n293) );
  NAND2X0 U355 ( .IN1(A[7]), .IN2(n449), .QN(n113) );
  NAND2X0 U356 ( .IN1(n247), .IN2(n245), .QN(n251) );
  NAND2X0 U357 ( .IN1(n427), .IN2(n247), .QN(n244) );
  NAND2X1 U358 ( .IN1(n248), .IN2(n247), .QN(n238) );
  NOR2X0 U359 ( .IN1(n232), .IN2(n384), .QN(n231) );
  NAND2X0 U360 ( .IN1(n384), .IN2(n219), .QN(n216) );
  NAND2X0 U361 ( .IN1(n29), .IN2(n30), .QN(n43) );
  NAND2X0 U362 ( .IN1(n33), .IN2(n32), .QN(n29) );
  NAND2X0 U363 ( .IN1(n218), .IN2(n99), .QN(n96) );
  NAND2X0 U364 ( .IN1(n39), .IN2(n35), .QN(n32) );
  NOR2X0 U365 ( .IN1(n287), .IN2(n286), .QN(n280) );
  NAND2X0 U366 ( .IN1(n1), .IN2(n55), .QN(n54) );
  NAND2X0 U367 ( .IN1(n328), .IN2(n329), .QN(n327) );
  NAND2X0 U368 ( .IN1(n289), .IN2(n129), .QN(n336) );
  NAND2X0 U369 ( .IN1(n134), .IN2(n464), .QN(n346) );
  NAND2X0 U370 ( .IN1(n1), .IN2(n208), .QN(n205) );
  INVX0 U371 ( (A[8]), (n484) );
  NAND2X0 U372 ( .IN1(n176), .IN2(n50), .QN(n47) );
  NAND2X0 U373 ( .IN1(n32), .IN2(n33), .QN(n75) );
  NAND2X0 U374 ( .IN1(n236), .IN2(n235), .QN(n233) );
  NAND2X0 U381 ( .IN1(n315), .IN2(n316), .QN(n312) );
  NAND2X0 U397 ( .IN1(n284), .IN2(n108), .QN(n316) );
  NAND2X0 U398 ( .IN1(n312), .IN2(n294), .QN(n311) );
  NAND2X1 U407 ( .IN1(B[3]), .IN2(n488), .QN(n134) );
  INVX0 U408 ( (A[3]), (n488) );
endmodule


module BoothMultiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17,
         n18, n21, n22, n26, n27, n29, n30, n31, n32, n34, n36, n39, n40, n42,
         n43, n46, n48, n50, n51, n54, n56, n58, n59, n61, n62, n63, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n76, n77, n79, n80, n82, n83,
         n84, n85, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n99,
         n100, n101, n102, n103, n105, n106, n107, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n120, n121, n122, n123, n126,
         n127, n128, n131, n132, n135, n136, n137, n138, n139, n140, n142,
         n143, n146, n147, n148, n149, n152, n155, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n172,
         n173, n174, n175, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n255,
         n256, n257, n259, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n276, n277, n278, n279, n280,
         n281, n282, n283, n286, n287, n288, n289, n290, n291, n292, n293,
         n295, n296, n297, n298, n299, n300, n303, n304, n305, n306, n307,
         n310, n311, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366;

  AND2X1 U2 ( .IN1(B[28]), .IN2(A[28]), .Q(n22) );
  AND2X1 U5 ( .IN1(n165), .IN2(n162), .Q(n58) );
  AND2X1 U7 ( .IN1(B[16]), .IN2(A[16]), .Q(n66) );
  AND2X1 U11 ( .IN1(n31), .IN2(n282), .Q(n289) );
  XOR3X1 U13 ( .IN1(B[30]), .IN2(A[30]), .IN3(n143), .Q(SUM[30]) );
  AND2X1 U15 ( .IN1(n182), .IN2(n183), .Q(n2) );
  AND2X1 U16 ( .IN1(B[1]), .IN2(A[1]), .Q(n3) );
  AND2X1 U17 ( .IN1(n212), .IN2(n211), .Q(SUM[0]) );
  OR2X1 U20 ( .IN1(B[8]), .IN2(A[8]), .Q(n109) );
  AND2X1 U27 ( .IN1(n165), .IN2(n170), .Q(n10) );
  AND2X1 U31 ( .IN1(n54), .IN2(n22), .Q(n13) );
  OR2X1 U35 ( .IN1(B[28]), .IN2(A[28]), .Q(n158) );
  AND2X1 U38 ( .IN1(n178), .IN2(n85), .Q(n16) );
  OR2X1 U53 ( .IN1(n345), .IN2(n165), .Q(n27) );
  AND2X1 U54 ( .IN1(n167), .IN2(n164), .Q(n29) );
  XOR3X1 U55 ( .IN1(B[28]), .IN2(A[28]), .IN3(n159), .Q(SUM[28]) );
  AND2X1 U56 ( .IN1(n30), .IN2(n31), .Q(n281) );
  AND2X1 U63 ( .IN1(n39), .IN2(n80), .Q(n36) );
  AND2X1 U66 ( .IN1(n42), .IN2(n74), .Q(n39) );
  AND2X1 U69 ( .IN1(n46), .IN2(n68), .Q(n42) );
  AND2X1 U71 ( .IN1(n303), .IN2(n139), .Q(n298) );
  AND2X1 U74 ( .IN1(n178), .IN2(n63), .Q(n46) );
  XOR3X1 U75 ( .IN1(B[31]), .IN2(A[31]), .IN3(n140), .Q(SUM[31]) );
  OR2X1 U79 ( .IN1(n344), .IN2(n167), .Q(n48) );
  AND2X1 U81 ( .IN1(n170), .IN2(n58), .Q(n50) );
  AND2X1 U84 ( .IN1(n148), .IN2(n142), .Q(n54) );
  OR2X1 U86 ( .IN1(n343), .IN2(n164), .Q(n56) );
  OR2X1 U90 ( .IN1(n342), .IN2(n173), .Q(n63) );
  AND2X1 U92 ( .IN1(n175), .IN2(n69), .Q(n65) );
  OR2X1 U94 ( .IN1(n11), .IN2(n167), .Q(n68) );
  AND2X1 U95 ( .IN1(n82), .IN2(n10), .Q(n69) );
  OR2X1 U97 ( .IN1(n18), .IN2(n217), .Q(n71) );
  AND2X1 U98 ( .IN1(n219), .IN2(n99), .Q(n72) );
  OR2X1 U100 ( .IN1(n340), .IN2(n164), .Q(n74) );
  AND2X1 U104 ( .IN1(n194), .IN2(n350), .Q(n77) );
  OR2X1 U106 ( .IN1(B[21]), .IN2(A[21]), .Q(n190) );
  OR2X1 U108 ( .IN1(n338), .IN2(n160), .Q(n80) );
  AND2X1 U110 ( .IN1(n162), .IN2(n158), .Q(n82) );
  AND2X1 U124 ( .IN1(n84), .IN2(n85), .Q(n179) );
  OR2X1 U125 ( .IN1(n348), .IN2(n182), .Q(n85) );
  AND2X1 U127 ( .IN1(n185), .IN2(n180), .Q(n87) );
  AND2X1 U129 ( .IN1(n251), .IN2(n252), .Q(n89) );
  AND2X1 U134 ( .IN1(n208), .IN2(n198), .Q(n99) );
  OR2X1 U139 ( .IN1(n209), .IN2(n88), .Q(n201) );
  NAND3X0 U142 ( .IN1(n257), .IN2(n355), .IN3(n259), .QN(n256) );
  AND2X1 U171 ( .IN1(n238), .IN2(n257), .Q(n262) );
  AND2X1 U182 ( .IN1(n112), .IN2(n113), .Q(n92) );
  AND2X1 U183 ( .IN1(n246), .IN2(n280), .Q(n93) );
  OR2X1 U186 ( .IN1(B[13]), .IN2(A[13]), .Q(n270) );
  OR2X1 U188 ( .IN1(B[4]), .IN2(A[4]), .Q(n128) );
  OR2X1 U189 ( .IN1(B[16]), .IN2(A[16]), .Q(n228) );
  OR2X1 U195 ( .IN1(B[12]), .IN2(A[12]), .Q(n274) );
  OR2X1 U198 ( .IN1(B[7]), .IN2(A[7]), .Q(n112) );
  OR2X1 U200 ( .IN1(B[11]), .IN2(A[11]), .Q(n246) );
  OR2X1 U201 ( .IN1(B[18]), .IN2(A[18]), .Q(n219) );
  OR2X1 U202 ( .IN1(B[19]), .IN2(A[19]), .Q(n208) );
  OR2X1 U204 ( .IN1(A[17]), .IN2(B[17]), .Q(n227) );
  OR2X1 U211 ( .IN1(B[26]), .IN2(A[26]), .Q(n165) );
  OR2X1 U213 ( .IN1(B[23]), .IN2(A[23]), .Q(n180) );
  OR2X1 U214 ( .IN1(B[27]), .IN2(A[27]), .Q(n162) );
  OR2X1 U215 ( .IN1(B[22]), .IN2(A[22]), .Q(n185) );
  OR2X1 U216 ( .IN1(B[0]), .IN2(A[0]), .Q(n212) );
  NAND3X0 U223 ( .IN1(n243), .IN2(n244), .IN3(n242), .QN(n235) );
  AND2X1 U238 ( .IN1(n257), .IN2(n259), .Q(n252) );
  AND2X1 U253 ( .IN1(n270), .IN2(n274), .Q(n251) );
  XOR2X1 U312 ( .IN1(n102), .IN2(n103), .Q(SUM[9]) );
  XOR2X1 U314 ( .IN1(n111), .IN2(n92), .Q(SUM[7]) );
  XOR2X1 U315 ( .IN1(n116), .IN2(n118), .Q(SUM[6]) );
  XOR2X1 U318 ( .IN1(n131), .IN2(n132), .Q(SUM[3]) );
  XOR2X1 U319 ( .IN1(n138), .IN2(n152), .Q(SUM[2]) );
  XOR2X1 U320 ( .IN1(n32), .IN2(n163), .Q(SUM[27]) );
  XOR2X1 U321 ( .IN1(n1), .IN2(n166), .Q(SUM[26]) );
  XOR2X1 U322 ( .IN1(n346), .IN2(n172), .Q(SUM[25]) );
  XOR2X1 U323 ( .IN1(n347), .IN2(n177), .Q(SUM[24]) );
  XOR2X1 U324 ( .IN1(n2), .IN2(n181), .Q(SUM[23]) );
  XOR2X1 U325 ( .IN1(n186), .IN2(n349), .Q(SUM[22]) );
  XOR2X1 U326 ( .IN1(n192), .IN2(n191), .Q(SUM[21]) );
  XOR2X1 U327 ( .IN1(n202), .IN2(n203), .Q(SUM[20]) );
  XOR2X1 U328 ( .IN1(n210), .IN2(n211), .Q(SUM[1]) );
  XOR2X1 U329 ( .IN1(n213), .IN2(n214), .Q(SUM[19]) );
  XOR2X1 U330 ( .IN1(n222), .IN2(n223), .Q(SUM[18]) );
  XOR2X1 U331 ( .IN1(n229), .IN2(n230), .Q(SUM[17]) );
  XOR2X1 U332 ( .IN1(n234), .IN2(n94), .Q(SUM[16]) );
  NAND4X0 U333 ( .IN1(n241), .IN2(n89), .IN3(n17), .IN4(n239), .QN(n237) );
  NAND4X0 U334 ( .IN1(n245), .IN2(n89), .IN3(n240), .IN4(n112), .QN(n244) );
  NAND3X0 U335 ( .IN1(n89), .IN2(n246), .IN3(n247), .QN(n243) );
  XOR2X1 U336 ( .IN1(n261), .IN2(n262), .Q(SUM[15]) );
  NAND3X0 U340 ( .IN1(n281), .IN2(n280), .IN3(n279), .QN(n247) );
  NAND3X0 U341 ( .IN1(n282), .IN2(n105), .IN3(n283), .QN(n279) );
  XOR2X1 U342 ( .IN1(n286), .IN2(n93), .Q(SUM[11]) );
  XOR2X1 U343 ( .IN1(n288), .IN2(n289), .Q(SUM[10]) );
  NAND4X0 U344 ( .IN1(n297), .IN2(n296), .IN3(n295), .IN4(n135), .QN(n241) );
  NAND4X0 U345 ( .IN1(B[4]), .IN2(A[4]), .IN3(n96), .IN4(n117), .QN(n307) );
  INVX0 U3 ( (n74), (n339) );
  INVX0 U4 ( (n142), (n337) );
  XNOR2X1 U6 ( .IN1(n317), .IN2(n314), .Q(SUM[4]) );
  NAND2X1 U8 ( .IN1(n126), .IN2(n128), .QN(n314) );
  XNOR2X1 U9 ( .IN1(n122), .IN2(n315), .Q(SUM[5]) );
  NAND2X1 U10 ( .IN1(n120), .IN2(n96), .QN(n315) );
  NAND2X0 U12 ( .IN1(n173), .IN2(n174), .QN(n316) );
  NBUFFX2 U14 ( (n241), (n317) );
  NOR2X0 U18 ( .IN1(n94), .IN2(n221), .QN(n224) );
  NOR2X0 U19 ( .IN1(n215), .IN2(n207), .QN(n214) );
  NOR2X0 U21 ( .IN1(n94), .IN2(n209), .QN(n215) );
  INVX0 U22 ( (n316), (n346) );
  INVX0 U23 ( (n67), (n349) );
  NAND2X1 U24 ( .IN1(n80), .IN2(n318), .QN(n34) );
  NOR2X0 U25 ( .IN1(n339), .IN2(n40), .QN(n318) );
  INVX0 U26 ( (n63), (n341) );
  NBUFFX2 U28 ( (n115), (n332) );
  NAND3X0 U29 ( .IN1(n139), .IN2(n6), .IN3(n3), .QN(n296) );
  NOR2X0 U30 ( .IN1(n94), .IN2(n200), .QN(n193) );
  NOR2X0 U32 ( .IN1(n365), .IN2(n358), .QN(n283) );
  NAND2X1 U33 ( .IN1(n123), .IN2(n128), .QN(n304) );
  NAND2X1 U34 ( .IN1(n292), .IN2(n293), .QN(n107) );
  NOR2X0 U36 ( .IN1(n351), .IN2(n206), .QN(n9) );
  INVX0 U37 ( (n332), (n359) );
  NOR2X0 U39 ( .IN1(n319), .IN2(n320), .QN(n161) );
  NAND2X1 U40 ( .IN1(n56), .IN2(n48), .QN(n319) );
  AND2X1 U41 ( .IN1(n169), .IN2(n50), .Q(n320) );
  INVX0 U42 ( (n83), (n350) );
  AND2X1 U43 ( .IN1(n190), .IN2(n198), .Q(n62) );
  NAND2X1 U44 ( .IN1(n114), .IN2(n332), .QN(n111) );
  NOR2X0 U45 ( .IN1(n231), .IN2(n66), .QN(n230) );
  NOR2X0 U46 ( .IN1(n352), .IN2(n94), .QN(n231) );
  INVX0 U47 ( (n228), (n352) );
  NAND2X1 U48 ( .IN1(n126), .IN2(n127), .QN(n122) );
  NAND2X1 U49 ( .IN1(n216), .IN2(n217), .QN(n207) );
  NOR2X0 U50 ( .IN1(n204), .IN2(n197), .QN(n203) );
  NAND2X1 U51 ( .IN1(n205), .IN2(n206), .QN(n197) );
  NOR2X0 U52 ( .IN1(n94), .IN2(n201), .QN(n204) );
  NAND2X1 U57 ( .IN1(n207), .IN2(n208), .QN(n205) );
  NAND2X1 U58 ( .IN1(n164), .IN2(n165), .QN(n166) );
  AND2X1 U59 ( .IN1(n167), .IN2(n168), .Q(n1) );
  AND2X1 U60 ( .IN1(n179), .IN2(n36), .Q(n330) );
  NAND2X1 U61 ( .IN1(n273), .IN2(n274), .QN(n272) );
  INVX0 U62 ( (n267), (n355) );
  NOR2X0 U64 ( .IN1(n209), .IN2(n88), .QN(n61) );
  NAND2X1 U65 ( .IN1(n276), .IN2(n277), .QN(n273) );
  NAND2X1 U67 ( .IN1(n334), .IN2(n107), .QN(n277) );
  XOR2X1 U68 ( .IN1(n269), .IN2(n271), .Q(SUM[13]) );
  NAND2X1 U70 ( .IN1(n120), .IN2(n121), .QN(n116) );
  NAND2X1 U72 ( .IN1(n122), .IN2(n97), .QN(n121) );
  NOR2X0 U73 ( .IN1(n321), .IN2(n322), .QN(n149) );
  AND2X1 U76 ( .IN1(n179), .IN2(n328), .Q(n321) );
  NOR2X0 U77 ( .IN1(n22), .IN2(n34), .QN(n322) );
  NAND2X1 U78 ( .IN1(n110), .IN2(n291), .QN(n102) );
  NAND2X1 U80 ( .IN1(n109), .IN2(n107), .QN(n291) );
  NAND2X1 U82 ( .IN1(n67), .IN2(n185), .QN(n183) );
  NAND2X1 U83 ( .IN1(n165), .IN2(n82), .QN(n11) );
  XOR2X1 U85 ( .IN1(n265), .IN2(n266), .Q(SUM[14]) );
  NAND2X1 U87 ( .IN1(n190), .IN2(n188), .QN(n192) );
  NOR2X0 U88 ( .IN1(n193), .IN2(n43), .QN(n191) );
  XNOR2X1 U89 ( .IN1(n273), .IN2(n323), .Q(SUM[12]) );
  NAND2X1 U91 ( .IN1(n250), .IN2(n274), .QN(n323) );
  NAND2X1 U93 ( .IN1(n160), .IN2(n162), .QN(n163) );
  NAND2X1 U96 ( .IN1(n263), .IN2(n264), .QN(n261) );
  INVX0 U99 ( (n82), (n340) );
  NAND2X1 U101 ( .IN1(n68), .IN2(n324), .QN(n40) );
  NOR2X0 U102 ( .IN1(n341), .IN2(n65), .QN(n324) );
  INVX0 U103 ( (n180), (n348) );
  INVX0 U105 ( (n58), (n344) );
  INVX0 U107 ( (n158), (n338) );
  INVX0 U109 ( (n259), (n354) );
  NOR2X0 U111 ( .IN1(n73), .IN2(n357), .QN(n103) );
  NAND2X1 U112 ( .IN1(n157), .IN2(n5), .QN(n210) );
  NAND2X1 U113 ( .IN1(n167), .IN2(n170), .QN(n172) );
  NAND2X1 U114 ( .IN1(n198), .IN2(n196), .QN(n202) );
  NAND2X1 U115 ( .IN1(n173), .IN2(n175), .QN(n177) );
  NOR2X0 U116 ( .IN1(n355), .IN2(n356), .QN(n271) );
  INVX0 U117 ( (n270), (n356) );
  NAND2X1 U118 ( .IN1(n208), .IN2(n206), .QN(n213) );
  NAND2X1 U119 ( .IN1(n219), .IN2(n217), .QN(n222) );
  NAND2X1 U120 ( .IN1(n5), .IN2(n155), .QN(n138) );
  NAND2X1 U121 ( .IN1(n364), .IN2(n157), .QN(n155) );
  INVX0 U122 ( (n211), (n364) );
  NAND2X1 U123 ( .IN1(n185), .IN2(n182), .QN(n186) );
  NAND2X1 U126 ( .IN1(n178), .IN2(n180), .QN(n181) );
  XNOR2X1 U128 ( .IN1(n107), .IN2(n325), .Q(SUM[8]) );
  NAND2X1 U130 ( .IN1(n110), .IN2(n109), .QN(n325) );
  INVX0 U131 ( (n164), (n345) );
  INVX0 U132 ( (n162), (n343) );
  NAND2X1 U133 ( .IN1(n106), .IN2(n290), .QN(n288) );
  NOR2X0 U135 ( .IN1(B[19]), .IN2(A[19]), .QN(n88) );
  NAND2X1 U136 ( .IN1(B[26]), .IN2(A[26]), .QN(n164) );
  NAND2X1 U137 ( .IN1(B[19]), .IN2(A[19]), .QN(n206) );
  NAND2X1 U138 ( .IN1(B[18]), .IN2(A[18]), .QN(n217) );
  NAND2X1 U140 ( .IN1(B[21]), .IN2(A[21]), .QN(n188) );
  NAND2X1 U141 ( .IN1(B[22]), .IN2(A[22]), .QN(n182) );
  NAND2X1 U143 ( .IN1(B[27]), .IN2(A[27]), .QN(n160) );
  NAND2X1 U144 ( .IN1(B[23]), .IN2(A[23]), .QN(n178) );
  NOR2X0 U145 ( .IN1(B[21]), .IN2(A[21]), .QN(n83) );
  AND2X1 U146 ( .IN1(A[2]), .IN2(B[2]), .Q(n335) );
  OR2X1 U147 ( .IN1(B[25]), .IN2(A[25]), .Q(n170) );
  OR2X1 U148 ( .IN1(B[9]), .IN2(A[9]), .Q(n105) );
  OR2X1 U149 ( .IN1(B[24]), .IN2(A[24]), .Q(n175) );
  OR2X1 U150 ( .IN1(A[10]), .IN2(B[10]), .Q(n282) );
  NAND2X0 U151 ( .IN1(B[16]), .IN2(A[16]), .QN(n232) );
  NAND2X1 U152 ( .IN1(B[12]), .IN2(A[12]), .QN(n250) );
  OR2X1 U153 ( .IN1(A[20]), .IN2(B[20]), .Q(n198) );
  XOR3X1 U154 ( .IN1(B[29]), .IN2(A[29]), .IN3(n149), .Q(SUM[29]) );
  NAND2X1 U155 ( .IN1(B[11]), .IN2(A[11]), .QN(n280) );
  AND2X1 U156 ( .IN1(A[9]), .IN2(B[9]), .Q(n73) );
  OR2X1 U157 ( .IN1(A[2]), .IN2(B[2]), .Q(n139) );
  OR2X1 U158 ( .IN1(A[3]), .IN2(B[3]), .Q(n6) );
  OR2X1 U159 ( .IN1(B[6]), .IN2(A[6]), .Q(n117) );
  OR2X1 U160 ( .IN1(A[3]), .IN2(B[3]), .Q(n303) );
  NAND2X1 U161 ( .IN1(B[4]), .IN2(A[4]), .QN(n126) );
  OR2X1 U162 ( .IN1(B[1]), .IN2(A[1]), .Q(n157) );
  NAND2X1 U163 ( .IN1(B[29]), .IN2(A[29]), .QN(n146) );
  NAND2X1 U164 ( .IN1(B[0]), .IN2(A[0]), .QN(n211) );
  OR2X1 U165 ( .IN1(B[29]), .IN2(A[29]), .Q(n148) );
  NAND2X1 U166 ( .IN1(B[8]), .IN2(A[8]), .QN(n110) );
  OR2X1 U167 ( .IN1(B[30]), .IN2(A[30]), .Q(n142) );
  NOR2X0 U168 ( .IN1(n326), .IN2(n327), .QN(n21) );
  AND2X1 U169 ( .IN1(B[30]), .IN2(A[30]), .Q(n326) );
  NOR2X0 U170 ( .IN1(n337), .IN2(n146), .QN(n327) );
  INVX0 U172 ( (B[8]), (n358) );
  INVX0 U173 ( (B[5]), (n360) );
  INVX0 U174 ( (n69), (n342) );
  AND2X1 U175 ( .IN1(n36), .IN2(n329), .Q(n328) );
  INVX0 U176 ( (n22), (n329) );
  NAND2X0 U177 ( .IN1(B[24]), .IN2(A[24]), .QN(n173) );
  NOR2X0 U178 ( .IN1(n330), .IN2(n331), .QN(n12) );
  NAND2X0 U179 ( .IN1(n54), .IN2(n34), .QN(n331) );
  OR2X1 U180 ( .IN1(A[10]), .IN2(B[10]), .Q(n278) );
  NAND2X1 U181 ( .IN1(n26), .IN2(n27), .QN(n32) );
  NAND2X0 U184 ( .IN1(B[13]), .IN2(A[13]), .QN(n267) );
  INVX0 U185 ( (n6), (n362) );
  INVX0 U187 ( (n135), (n361) );
  NOR2X0 U190 ( .IN1(n361), .IN2(n362), .QN(n132) );
  NAND2X0 U191 ( .IN1(B[15]), .IN2(A[15]), .QN(n238) );
  OR2X1 U192 ( .IN1(B[15]), .IN2(A[15]), .Q(n257) );
  OR2X1 U193 ( .IN1(B[14]), .IN2(A[14]), .Q(n259) );
  NAND2X0 U194 ( .IN1(B[14]), .IN2(A[14]), .QN(n263) );
  NAND2X1 U196 ( .IN1(n138), .IN2(n139), .QN(n137) );
  INVX0 U197 ( (n139), (n363) );
  NAND2X1 U199 ( .IN1(n136), .IN2(n137), .QN(n131) );
  NAND2X0 U203 ( .IN1(n225), .IN2(n226), .QN(n218) );
  INVX0 U205 ( (n333), (n221) );
  NAND2X1 U206 ( .IN1(n333), .IN2(n219), .QN(n209) );
  AND2X1 U207 ( .IN1(n228), .IN2(n227), .Q(n333) );
  NAND2X0 U208 ( .IN1(B[20]), .IN2(A[20]), .QN(n196) );
  NAND2X0 U209 ( .IN1(B[3]), .IN2(A[3]), .QN(n135) );
  NAND2X0 U210 ( .IN1(B[25]), .IN2(A[25]), .QN(n167) );
  NOR2X0 U212 ( .IN1(A[6]), .IN2(B[6]), .QN(n100) );
  NAND2X0 U217 ( .IN1(n208), .IN2(n198), .QN(n18) );
  INVX0 U218 ( (n198), (n351) );
  NOR2X0 U219 ( .IN1(A[1]), .IN2(B[1]), .QN(n95) );
  NAND2X0 U220 ( .IN1(B[1]), .IN2(A[1]), .QN(n5) );
  NAND2X0 U221 ( .IN1(B[6]), .IN2(A[6]), .QN(n115) );
  NAND2X1 U222 ( .IN1(n288), .IN2(n282), .QN(n287) );
  NAND2X0 U224 ( .IN1(n31), .IN2(n287), .QN(n286) );
  NAND2X0 U225 ( .IN1(n278), .IN2(n73), .QN(n30) );
  NAND2X0 U226 ( .IN1(B[9]), .IN2(A[9]), .QN(n106) );
  NOR2X0 U227 ( .IN1(n7), .IN2(n91), .QN(n240) );
  INVX0 U228 ( (n335), (n136) );
  NAND2X0 U229 ( .IN1(n335), .IN2(n6), .QN(n295) );
  NOR2X0 U230 ( .IN1(n335), .IN2(n363), .QN(n152) );
  NAND2X0 U231 ( .IN1(n360), .IN2(n366), .QN(n97) );
  NAND2X0 U232 ( .IN1(n360), .IN2(n366), .QN(n96) );
  NOR2X0 U233 ( .IN1(n90), .IN2(n91), .QN(n334) );
  NOR2X0 U234 ( .IN1(n90), .IN2(n91), .QN(n17) );
  NAND2X0 U235 ( .IN1(n278), .IN2(n246), .QN(n91) );
  NAND2X0 U236 ( .IN1(n105), .IN2(n109), .QN(n90) );
  NAND2X0 U237 ( .IN1(n105), .IN2(n102), .QN(n290) );
  NAND2X0 U239 ( .IN1(n105), .IN2(n109), .QN(n7) );
  INVX0 U240 ( (n105), (n357) );
  NAND2X0 U241 ( .IN1(n227), .IN2(n226), .QN(n229) );
  NAND2X0 U242 ( .IN1(n66), .IN2(n227), .QN(n225) );
  NAND2X0 U243 ( .IN1(B[17]), .IN2(A[17]), .QN(n226) );
  NOR2X0 U244 ( .IN1(n249), .IN2(n248), .QN(n242) );
  NAND2X1 U245 ( .IN1(n255), .IN2(n256), .QN(n248) );
  NAND2X0 U246 ( .IN1(n116), .IN2(n117), .QN(n114) );
  NOR2X0 U247 ( .IN1(n304), .IN2(n305), .QN(n239) );
  NAND2X0 U248 ( .IN1(n353), .IN2(n257), .QN(n255) );
  NOR2X0 U249 ( .IN1(n353), .IN2(n354), .QN(n266) );
  INVX0 U250 ( (n263), (n353) );
  NAND2X0 U251 ( .IN1(B[10]), .IN2(A[10]), .QN(n31) );
  NAND2X0 U252 ( .IN1(n247), .IN2(n246), .QN(n276) );
  NAND2X0 U254 ( .IN1(n113), .IN2(n115), .QN(n310) );
  NAND2X0 U255 ( .IN1(n307), .IN2(n306), .QN(n336) );
  NOR2X0 U256 ( .IN1(n95), .IN2(n300), .QN(n299) );
  NOR2X0 U257 ( .IN1(n359), .IN2(n100), .QN(n118) );
  NAND2X0 U258 ( .IN1(n29), .IN2(n168), .QN(n26) );
  NAND2X0 U259 ( .IN1(n336), .IN2(n112), .QN(n292) );
  NOR2X0 U260 ( .IN1(n120), .IN2(n100), .QN(n311) );
  NAND2X0 U261 ( .IN1(n160), .IN2(n161), .QN(n159) );
  INVX0 U262 ( (A[5]), (n366) );
  NAND2X0 U263 ( .IN1(n360), .IN2(n366), .QN(n123) );
  NAND2X0 U264 ( .IN1(n265), .IN2(n259), .QN(n264) );
  NAND2X0 U265 ( .IN1(n267), .IN2(n268), .QN(n265) );
  NAND2X0 U266 ( .IN1(n269), .IN2(n270), .QN(n268) );
  NAND2X1 U267 ( .IN1(n272), .IN2(n250), .QN(n269) );
  NOR2X0 U268 ( .IN1(n101), .IN2(n250), .QN(n249) );
  NAND2X0 U269 ( .IN1(n251), .IN2(n252), .QN(n101) );
  NOR2X0 U270 ( .IN1(n199), .IN2(n79), .QN(n76) );
  NAND2X0 U271 ( .IN1(n146), .IN2(n147), .QN(n143) );
  NAND2X0 U272 ( .IN1(n195), .IN2(n196), .QN(n43) );
  NAND2X0 U273 ( .IN1(n195), .IN2(n196), .QN(n194) );
  NOR2X0 U274 ( .IN1(n8), .IN2(n9), .QN(n195) );
  INVX0 U275 ( (n59), (n347) );
  NAND2X0 U276 ( .IN1(n112), .IN2(n117), .QN(n305) );
  NAND2X0 U277 ( .IN1(n15), .IN2(n16), .QN(n59) );
  NOR2X0 U278 ( .IN1(n12), .IN2(n13), .QN(n51) );
  NAND2X0 U279 ( .IN1(B[7]), .IN2(A[7]), .QN(n113) );
  NAND2X0 U280 ( .IN1(n228), .IN2(n232), .QN(n234) );
  NAND2X0 U281 ( .IN1(n61), .IN2(n198), .QN(n200) );
  NAND2X0 U282 ( .IN1(n184), .IN2(n87), .QN(n84) );
  NAND2X0 U283 ( .IN1(n184), .IN2(n87), .QN(n15) );
  NAND2X0 U284 ( .IN1(n61), .IN2(n62), .QN(n79) );
  NAND2X0 U285 ( .IN1(n70), .IN2(n71), .QN(n8) );
  NAND2X0 U286 ( .IN1(n188), .IN2(n189), .QN(n184) );
  NAND2X0 U287 ( .IN1(n51), .IN2(n21), .QN(n140) );
  NOR2X0 U288 ( .IN1(n235), .IN2(n236), .QN(n94) );
  NOR2X0 U289 ( .IN1(n235), .IN2(n236), .QN(n199) );
  NAND2X1 U290 ( .IN1(B[5]), .IN2(A[5]), .QN(n120) );
  NAND2X0 U291 ( .IN1(n306), .IN2(n307), .QN(n245) );
  NOR2X0 U292 ( .IN1(n311), .IN2(n310), .QN(n306) );
  NOR2X0 U293 ( .IN1(n76), .IN2(n77), .QN(n189) );
  NAND2X0 U294 ( .IN1(B[0]), .IN2(A[0]), .QN(n300) );
  INVX0 U295 ( (A[8]), (n365) );
  NOR2X0 U296 ( .IN1(n224), .IN2(n218), .QN(n223) );
  NAND2X0 U297 ( .IN1(n148), .IN2(n149), .QN(n147) );
  NAND2X0 U298 ( .IN1(n188), .IN2(n189), .QN(n67) );
  NAND2X0 U299 ( .IN1(n218), .IN2(n219), .QN(n216) );
  NAND2X0 U300 ( .IN1(n218), .IN2(n72), .QN(n70) );
  NAND2X0 U301 ( .IN1(n173), .IN2(n174), .QN(n169) );
  NAND2X0 U302 ( .IN1(n316), .IN2(n170), .QN(n168) );
  NAND2X0 U303 ( .IN1(n128), .IN2(n317), .QN(n127) );
  NAND2X0 U304 ( .IN1(n239), .IN2(n317), .QN(n293) );
  NAND2X1 U305 ( .IN1(n237), .IN2(n238), .QN(n236) );
  NAND2X0 U306 ( .IN1(n59), .IN2(n175), .QN(n174) );
  NAND2X0 U307 ( .IN1(n298), .IN2(n299), .QN(n297) );
endmodule


module BoothMultiplier ( clk, oClk, rst, oRst, M, Q, P );
  input [31:0] M;
  input [31:0] Q;
  output [63:0] P;
  input clk, oClk, rst, oRst;
  wire   n141, n142, n143, n148, n149, n150, n152, n153, n154, n155, n159,
         n160, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n310, n312, n314, n315, n318, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n618, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678;
  wire   [31:0] Acc;
  wire   [31:0] Q_reg;
  wire   [31:0] M_reg;
  wire   [64:33] case_add;
  wire   [64:33] case_sub;

  LATCHX1 \M_reg_reg[31]  ( .CLK(n663), .D(M[31]), .Q(M_reg[31]) );
  LATCHX1 \M_reg_reg[30]  ( .CLK(n663), .D(M[30]), .Q(M_reg[30]) );
  LATCHX1 \M_reg_reg[29]  ( .CLK(n663), .D(M[29]), .Q(M_reg[29]) );
  LATCHX1 \M_reg_reg[28]  ( .CLK(n663), .D(M[28]), .Q(M_reg[28]) );
  LATCHX1 \M_reg_reg[27]  ( .CLK(n663), .D(M[27]), .Q(M_reg[27]) );
  LATCHX1 \M_reg_reg[26]  ( .CLK(n663), .D(M[26]), .Q(M_reg[26]) );
  LATCHX1 \M_reg_reg[25]  ( .CLK(n663), .D(M[25]), .Q(M_reg[25]) );
  LATCHX1 \M_reg_reg[24]  ( .CLK(n663), .D(M[24]), .Q(M_reg[24]) );
  LATCHX1 \M_reg_reg[23]  ( .CLK(n663), .D(M[23]), .Q(M_reg[23]) );
  LATCHX1 \M_reg_reg[22]  ( .CLK(n663), .D(M[22]), .Q(M_reg[22]) );
  LATCHX1 \M_reg_reg[21]  ( .CLK(n663), .D(M[21]), .Q(M_reg[21]) );
  LATCHX1 \M_reg_reg[20]  ( .CLK(n663), .D(M[20]), .Q(M_reg[20]) );
  LATCHX1 \M_reg_reg[19]  ( .CLK(n663), .D(M[19]), .Q(M_reg[19]) );
  LATCHX1 \M_reg_reg[18]  ( .CLK(n663), .D(M[18]), .Q(M_reg[18]) );
  LATCHX1 \M_reg_reg[17]  ( .CLK(n663), .D(M[17]), .Q(M_reg[17]) );
  LATCHX1 \M_reg_reg[16]  ( .CLK(n663), .D(M[16]), .Q(M_reg[16]) );
  LATCHX1 \M_reg_reg[15]  ( .CLK(n663), .D(M[15]), .Q(M_reg[15]) );
  LATCHX1 \M_reg_reg[14]  ( .CLK(n663), .D(M[14]), .Q(M_reg[14]) );
  LATCHX1 \M_reg_reg[13]  ( .CLK(n663), .D(M[13]), .Q(M_reg[13]) );
  LATCHX1 \M_reg_reg[12]  ( .CLK(n663), .D(M[12]), .Q(M_reg[12]) );
  LATCHX1 \M_reg_reg[11]  ( .CLK(n663), .D(M[11]), .Q(M_reg[11]) );
  LATCHX1 \M_reg_reg[10]  ( .CLK(n663), .D(M[10]), .Q(M_reg[10]) );
  LATCHX1 \M_reg_reg[9]  ( .CLK(n663), .D(M[9]), .Q(M_reg[9]) );
  LATCHX1 \M_reg_reg[8]  ( .CLK(n662), .D(M[8]), .Q(M_reg[8]) );
  LATCHX1 \M_reg_reg[7]  ( .CLK(n662), .D(M[7]), .Q(M_reg[7]) );
  LATCHX1 \M_reg_reg[6]  ( .CLK(n662), .D(M[6]), .Q(M_reg[6]) );
  LATCHX1 \M_reg_reg[5]  ( .CLK(n662), .D(M[5]), .Q(M_reg[5]) );
  LATCHX1 \M_reg_reg[4]  ( .CLK(n662), .D(M[4]), .Q(M_reg[4]) );
  LATCHX1 \M_reg_reg[3]  ( .CLK(n662), .D(M[3]), .Q(M_reg[3]) );
  LATCHX1 \M_reg_reg[2]  ( .CLK(n662), .D(M[2]), .Q(M_reg[2]) );
  LATCHX1 \M_reg_reg[1]  ( .CLK(n662), .D(M[1]), .Q(M_reg[1]) );
  LATCHX1 \M_reg_reg[0]  ( .CLK(n662), .D(M[0]), .Q(M_reg[0]) );
  DFFARX1 \P_reg[63]  ( .D(Acc[31]), .CLK(oClk), .RSTB(n629), .Q(P[63]) );
  DFFARX1 \P_reg[62]  ( .D(Acc[31]), .CLK(oClk), .RSTB(n629), .Q(P[62]) );
  DFFARX1 \P_reg[61]  ( .D(Acc[30]), .CLK(oClk), .RSTB(n629), .Q(P[61]) );
  DFFARX1 \P_reg[60]  ( .D(Acc[29]), .CLK(oClk), .RSTB(n629), .Q(P[60]) );
  DFFARX1 \P_reg[59]  ( .D(Acc[28]), .CLK(oClk), .RSTB(n630), .Q(P[59]) );
  DFFARX1 \P_reg[58]  ( .D(Acc[27]), .CLK(oClk), .RSTB(n630), .Q(P[58]) );
  DFFARX1 \P_reg[57]  ( .D(Acc[26]), .CLK(oClk), .RSTB(n630), .Q(P[57]) );
  DFFARX1 \P_reg[56]  ( .D(Acc[25]), .CLK(oClk), .RSTB(n630), .Q(P[56]) );
  DFFARX1 \P_reg[55]  ( .D(Acc[24]), .CLK(oClk), .RSTB(n629), .Q(P[55]) );
  DFFARX1 \P_reg[54]  ( .D(Acc[23]), .CLK(oClk), .RSTB(n631), .Q(P[54]) );
  DFFARX1 \P_reg[53]  ( .D(Acc[22]), .CLK(oClk), .RSTB(n631), .Q(P[53]) );
  DFFARX1 \P_reg[52]  ( .D(Acc[21]), .CLK(oClk), .RSTB(n631), .Q(P[52]) );
  DFFARX1 \P_reg[51]  ( .D(Acc[20]), .CLK(oClk), .RSTB(n631), .Q(P[51]) );
  DFFARX1 \P_reg[50]  ( .D(n668), .CLK(oClk), .RSTB(n630), .Q(P[50]) );
  DFFARX1 \P_reg[49]  ( .D(Acc[18]), .CLK(oClk), .RSTB(n632), .Q(P[49]) );
  DFFARX1 \P_reg[48]  ( .D(Acc[17]), .CLK(oClk), .RSTB(n632), .Q(P[48]) );
  DFFARX1 \P_reg[47]  ( .D(Acc[16]), .CLK(oClk), .RSTB(n632), .Q(P[47]) );
  DFFARX1 \P_reg[46]  ( .D(Acc[15]), .CLK(oClk), .RSTB(n632), .Q(P[46]) );
  DFFARX1 \P_reg[45]  ( .D(n670), .CLK(oClk), .RSTB(n631), .Q(P[45]) );
  DFFARX1 \P_reg[44]  ( .D(n671), .CLK(oClk), .RSTB(n633), .Q(P[44]) );
  DFFARX1 \P_reg[43]  ( .D(n672), .CLK(oClk), .RSTB(n633), .Q(P[43]) );
  DFFARX1 \P_reg[42]  ( .D(Acc[11]), .CLK(oClk), .RSTB(n633), .Q(P[42]) );
  DFFARX1 \P_reg[41]  ( .D(n673), .CLK(oClk), .RSTB(n632), .Q(P[41]) );
  DFFARX1 \P_reg[40]  ( .D(n674), .CLK(oClk), .RSTB(n633), .Q(P[40]) );
  DFFARX1 \P_reg[39]  ( .D(n628), .CLK(oClk), .RSTB(n634), .Q(P[39]) );
  DFFARX1 \P_reg[38]  ( .D(Acc[7]), .CLK(oClk), .RSTB(n634), .Q(P[38]) );
  DFFARX1 \P_reg[37]  ( .D(Acc[6]), .CLK(oClk), .RSTB(n633), .Q(P[37]) );
  DFFARX1 \P_reg[36]  ( .D(Acc[5]), .CLK(oClk), .RSTB(n634), .Q(P[36]) );
  DFFARX1 \P_reg[35]  ( .D(n627), .CLK(oClk), .RSTB(n634), .Q(P[35]) );
  DFFARX1 \P_reg[34]  ( .D(n675), .CLK(oClk), .RSTB(n635), .Q(P[34]) );
  DFFARX1 \P_reg[33]  ( .D(Acc[2]), .CLK(oClk), .RSTB(n635), .Q(P[33]) );
  DFFARX1 \P_reg[32]  ( .D(n677), .CLK(oClk), .RSTB(n635), .Q(P[32]) );
  DFFARX1 \P_reg[31]  ( .D(Acc[0]), .CLK(oClk), .RSTB(n635), .Q(P[31]) );
  DFFARX1 \P_reg[30]  ( .D(Q_reg[31]), .CLK(oClk), .RSTB(n634), .Q(P[30]) );
  DFFARX1 \P_reg[29]  ( .D(Q_reg[30]), .CLK(oClk), .RSTB(n636), .Q(P[29]) );
  DFFARX1 \P_reg[28]  ( .D(Q_reg[29]), .CLK(oClk), .RSTB(n636), .Q(P[28]) );
  DFFARX1 \P_reg[27]  ( .D(Q_reg[28]), .CLK(oClk), .RSTB(n636), .Q(P[27]) );
  DFFARX1 \P_reg[26]  ( .D(Q_reg[27]), .CLK(oClk), .RSTB(n636), .Q(P[26]) );
  DFFARX1 \P_reg[25]  ( .D(Q_reg[26]), .CLK(oClk), .RSTB(n635), .Q(P[25]) );
  DFFARX1 \P_reg[24]  ( .D(Q_reg[25]), .CLK(oClk), .RSTB(n637), .Q(P[24]) );
  DFFARX1 \P_reg[23]  ( .D(Q_reg[24]), .CLK(oClk), .RSTB(n637), .Q(P[23]) );
  DFFARX1 \P_reg[22]  ( .D(Q_reg[23]), .CLK(oClk), .RSTB(n637), .Q(P[22]) );
  DFFARX1 \P_reg[21]  ( .D(Q_reg[22]), .CLK(oClk), .RSTB(n637), .Q(P[21]) );
  DFFARX1 \P_reg[20]  ( .D(Q_reg[21]), .CLK(oClk), .RSTB(n636), .Q(P[20]) );
  DFFARX1 \P_reg[19]  ( .D(Q_reg[20]), .CLK(oClk), .RSTB(n638), .Q(P[19]) );
  DFFARX1 \P_reg[18]  ( .D(Q_reg[19]), .CLK(oClk), .RSTB(n638), .Q(P[18]) );
  DFFARX1 \P_reg[17]  ( .D(Q_reg[18]), .CLK(oClk), .RSTB(n638), .Q(P[17]) );
  DFFARX1 \P_reg[16]  ( .D(Q_reg[17]), .CLK(oClk), .RSTB(n638), .Q(P[16]) );
  DFFARX1 \P_reg[15]  ( .D(Q_reg[16]), .CLK(oClk), .RSTB(n637), .Q(P[15]) );
  DFFARX1 \P_reg[14]  ( .D(Q_reg[15]), .CLK(oClk), .RSTB(n639), .Q(P[14]) );
  DFFARX1 \P_reg[13]  ( .D(Q_reg[14]), .CLK(oClk), .RSTB(n639), .Q(P[13]) );
  DFFARX1 \P_reg[12]  ( .D(Q_reg[13]), .CLK(oClk), .RSTB(n639), .Q(P[12]) );
  DFFARX1 \P_reg[11]  ( .D(Q_reg[12]), .CLK(oClk), .RSTB(n639), .Q(P[11]) );
  DFFARX1 \P_reg[10]  ( .D(Q_reg[11]), .CLK(oClk), .RSTB(n638), .Q(P[10]) );
  DFFARX1 \P_reg[9]  ( .D(Q_reg[10]), .CLK(oClk), .RSTB(n640), .Q(P[9]) );
  DFFARX1 \P_reg[8]  ( .D(Q_reg[9]), .CLK(oClk), .RSTB(n640), .Q(P[8]) );
  DFFARX1 \P_reg[7]  ( .D(Q_reg[8]), .CLK(oClk), .RSTB(n640), .Q(P[7]) );
  DFFARX1 \P_reg[6]  ( .D(Q_reg[7]), .CLK(oClk), .RSTB(n640), .Q(P[6]) );
  DFFARX1 \P_reg[5]  ( .D(Q_reg[6]), .CLK(oClk), .RSTB(n639), .Q(P[5]) );
  DFFARX1 \P_reg[4]  ( .D(Q_reg[5]), .CLK(oClk), .RSTB(n641), .Q(P[4]) );
  DFFARX1 \P_reg[3]  ( .D(Q_reg[4]), .CLK(oClk), .RSTB(n641), .Q(P[3]) );
  DFFARX1 \P_reg[2]  ( .D(Q_reg[3]), .CLK(oClk), .RSTB(n641), .Q(P[2]) );
  DFFARX1 \P_reg[1]  ( .D(Q_reg[2]), .CLK(oClk), .RSTB(n641), .Q(P[1]) );
  DFFARX1 \P_reg[0]  ( .D(Q_reg[1]), .CLK(oClk), .RSTB(n640), .Q(P[0]) );
  DFFASX1 \count_reg[0]  ( .D(n310), .CLK(clk), .SETB(n667), .QN(n312) );
  DFFASX1 \count_reg[1]  ( .D(n308), .CLK(clk), .SETB(n667), .QN(n315) );
  DFFASX1 \count_reg[2]  ( .D(n307), .CLK(clk), .SETB(n667), .QN(n620) );
  DFFASX1 \count_reg[3]  ( .D(n306), .CLK(clk), .SETB(n667), .Q(n624), .QN(
        n621) );
  DFFASX1 \count_reg[4]  ( .D(n305), .CLK(clk), .SETB(n667), .QN(n622) );
  DFFASRX1 \Q_reg_reg[0]  ( .D(n304), .CLK(clk), .RSTB(n238), .SETB(n237), .Q(
        n314) );
  DFFARX1 Q_prev_reg ( .D(n303), .CLK(clk), .RSTB(n664), .Q(n623), .QN(n318)
         );
  DFFARX1 \Acc_reg[31]  ( .D(n302), .CLK(clk), .RSTB(n665), .Q(Acc[31]) );
  DFFARX1 \Acc_reg[30]  ( .D(n301), .CLK(clk), .RSTB(n664), .Q(Acc[30]) );
  DFFARX1 \Acc_reg[29]  ( .D(n300), .CLK(clk), .RSTB(n664), .Q(Acc[29]) );
  DFFARX1 \Acc_reg[28]  ( .D(n299), .CLK(clk), .RSTB(n664), .Q(Acc[28]) );
  DFFARX1 \Acc_reg[27]  ( .D(n298), .CLK(clk), .RSTB(n664), .Q(Acc[27]) );
  DFFARX1 \Acc_reg[26]  ( .D(n297), .CLK(clk), .RSTB(n664), .Q(Acc[26]) );
  DFFARX1 \Acc_reg[25]  ( .D(n296), .CLK(clk), .RSTB(n664), .Q(Acc[25]) );
  DFFARX1 \Acc_reg[24]  ( .D(n295), .CLK(clk), .RSTB(n664), .Q(Acc[24]) );
  DFFARX1 \Acc_reg[23]  ( .D(n294), .CLK(clk), .RSTB(n664), .Q(Acc[23]) );
  DFFARX1 \Acc_reg[22]  ( .D(n293), .CLK(clk), .RSTB(n664), .Q(Acc[22]) );
  DFFARX1 \Acc_reg[21]  ( .D(n292), .CLK(clk), .RSTB(n664), .Q(Acc[21]) );
  DFFARX1 \Acc_reg[20]  ( .D(n291), .CLK(clk), .RSTB(n664), .Q(Acc[20]), .QN(
        n160) );
  DFFARX1 \Acc_reg[19]  ( .D(n290), .CLK(clk), .RSTB(n666), .Q(Acc[19]), .QN(
        n159) );
  DFFARX1 \Acc_reg[18]  ( .D(n289), .CLK(clk), .RSTB(n664), .Q(Acc[18]) );
  DFFARX1 \Acc_reg[17]  ( .D(n288), .CLK(clk), .RSTB(n667), .Q(Acc[17]) );
  DFFARX1 \Acc_reg[16]  ( .D(n287), .CLK(clk), .RSTB(n665), .Q(Acc[16]) );
  DFFARX1 \Acc_reg[15]  ( .D(n286), .CLK(clk), .RSTB(n666), .Q(Acc[15]), .QN(
        n155) );
  DFFARX1 \Acc_reg[14]  ( .D(n285), .CLK(clk), .RSTB(n664), .Q(Acc[14]), .QN(
        n154) );
  DFFARX1 \Acc_reg[13]  ( .D(n284), .CLK(clk), .RSTB(n667), .Q(Acc[13]), .QN(
        n153) );
  DFFARX1 \Acc_reg[12]  ( .D(n283), .CLK(clk), .RSTB(n665), .Q(Acc[12]), .QN(
        n152) );
  DFFARX1 \Acc_reg[11]  ( .D(n282), .CLK(clk), .RSTB(n666), .Q(Acc[11]) );
  DFFARX1 \Acc_reg[10]  ( .D(n281), .CLK(clk), .RSTB(n664), .Q(Acc[10]), .QN(
        n150) );
  DFFARX1 \Acc_reg[9]  ( .D(n280), .CLK(clk), .RSTB(n667), .Q(Acc[9]), .QN(
        n149) );
  DFFARX1 \Acc_reg[8]  ( .D(n279), .CLK(clk), .RSTB(n665), .Q(Acc[8]), .QN(
        n148) );
  DFFARX1 \Acc_reg[7]  ( .D(n278), .CLK(clk), .RSTB(n665), .Q(Acc[7]) );
  DFFARX1 \Acc_reg[6]  ( .D(n277), .CLK(clk), .RSTB(n665), .Q(Acc[6]) );
  DFFARX1 \Acc_reg[5]  ( .D(n276), .CLK(clk), .RSTB(n665), .Q(Acc[5]) );
  DFFARX1 \Acc_reg[4]  ( .D(n275), .CLK(clk), .RSTB(n665), .Q(Acc[4]), .QN(
        n618) );
  DFFARX1 \Acc_reg[3]  ( .D(n274), .CLK(clk), .RSTB(n665), .Q(Acc[3]), .QN(
        n143) );
  DFFARX1 \Acc_reg[2]  ( .D(n273), .CLK(clk), .RSTB(n665), .Q(Acc[2]), .QN(
        n142) );
  DFFARX1 \Acc_reg[1]  ( .D(n272), .CLK(clk), .RSTB(n665), .Q(Acc[1]), .QN(
        n141) );
  DFFARX1 \Acc_reg[0]  ( .D(n271), .CLK(clk), .RSTB(n665), .Q(Acc[0]) );
  DFFASRX1 \Q_reg_reg[31]  ( .D(n270), .CLK(clk), .RSTB(n236), .SETB(n235), 
        .Q(Q_reg[31]) );
  DFFASRX1 \Q_reg_reg[30]  ( .D(n269), .CLK(clk), .RSTB(n234), .SETB(n233), 
        .Q(Q_reg[30]) );
  DFFASRX1 \Q_reg_reg[29]  ( .D(n268), .CLK(clk), .RSTB(n232), .SETB(n231), 
        .Q(Q_reg[29]) );
  DFFASRX1 \Q_reg_reg[28]  ( .D(n267), .CLK(clk), .RSTB(n230), .SETB(n229), 
        .Q(Q_reg[28]) );
  DFFASRX1 \Q_reg_reg[27]  ( .D(n266), .CLK(clk), .RSTB(n228), .SETB(n227), 
        .Q(Q_reg[27]) );
  DFFASRX1 \Q_reg_reg[26]  ( .D(n265), .CLK(clk), .RSTB(n226), .SETB(n225), 
        .Q(Q_reg[26]) );
  DFFASRX1 \Q_reg_reg[25]  ( .D(n264), .CLK(clk), .RSTB(n224), .SETB(n223), 
        .Q(Q_reg[25]) );
  DFFASRX1 \Q_reg_reg[24]  ( .D(n263), .CLK(clk), .RSTB(n222), .SETB(n221), 
        .Q(Q_reg[24]) );
  DFFASRX1 \Q_reg_reg[23]  ( .D(n262), .CLK(clk), .RSTB(n220), .SETB(n219), 
        .Q(Q_reg[23]) );
  DFFASRX1 \Q_reg_reg[22]  ( .D(n261), .CLK(clk), .RSTB(n218), .SETB(n217), 
        .Q(Q_reg[22]) );
  DFFASRX1 \Q_reg_reg[21]  ( .D(n260), .CLK(clk), .RSTB(n216), .SETB(n215), 
        .Q(Q_reg[21]) );
  DFFASRX1 \Q_reg_reg[20]  ( .D(n259), .CLK(clk), .RSTB(n214), .SETB(n213), 
        .Q(Q_reg[20]) );
  DFFASRX1 \Q_reg_reg[19]  ( .D(n258), .CLK(clk), .RSTB(n212), .SETB(n211), 
        .Q(Q_reg[19]) );
  DFFASRX1 \Q_reg_reg[18]  ( .D(n257), .CLK(clk), .RSTB(n210), .SETB(n209), 
        .Q(Q_reg[18]) );
  DFFASRX1 \Q_reg_reg[17]  ( .D(n256), .CLK(clk), .RSTB(n208), .SETB(n207), 
        .Q(Q_reg[17]) );
  DFFASRX1 \Q_reg_reg[16]  ( .D(n255), .CLK(clk), .RSTB(n206), .SETB(n205), 
        .Q(Q_reg[16]) );
  DFFASRX1 \Q_reg_reg[15]  ( .D(n254), .CLK(clk), .RSTB(n204), .SETB(n203), 
        .Q(Q_reg[15]) );
  DFFASRX1 \Q_reg_reg[14]  ( .D(n253), .CLK(clk), .RSTB(n202), .SETB(n201), 
        .Q(Q_reg[14]) );
  DFFASRX1 \Q_reg_reg[13]  ( .D(n252), .CLK(clk), .RSTB(n200), .SETB(n199), 
        .Q(Q_reg[13]) );
  DFFASRX1 \Q_reg_reg[12]  ( .D(n251), .CLK(clk), .RSTB(n198), .SETB(n197), 
        .Q(Q_reg[12]) );
  DFFASRX1 \Q_reg_reg[11]  ( .D(n250), .CLK(clk), .RSTB(n196), .SETB(n195), 
        .Q(Q_reg[11]) );
  DFFASRX1 \Q_reg_reg[10]  ( .D(n249), .CLK(clk), .RSTB(n194), .SETB(n193), 
        .Q(Q_reg[10]) );
  DFFASRX1 \Q_reg_reg[9]  ( .D(n248), .CLK(clk), .RSTB(n192), .SETB(n191), .Q(
        Q_reg[9]) );
  DFFASRX1 \Q_reg_reg[8]  ( .D(n247), .CLK(clk), .RSTB(n190), .SETB(n189), .Q(
        Q_reg[8]) );
  DFFASRX1 \Q_reg_reg[7]  ( .D(n246), .CLK(clk), .RSTB(n188), .SETB(n187), .Q(
        Q_reg[7]) );
  DFFASRX1 \Q_reg_reg[6]  ( .D(n245), .CLK(clk), .RSTB(n186), .SETB(n185), .Q(
        Q_reg[6]) );
  DFFASRX1 \Q_reg_reg[5]  ( .D(n244), .CLK(clk), .RSTB(n184), .SETB(n183), .Q(
        Q_reg[5]) );
  DFFASRX1 \Q_reg_reg[4]  ( .D(n243), .CLK(clk), .RSTB(n182), .SETB(n181), .Q(
        Q_reg[4]) );
  DFFASRX1 \Q_reg_reg[3]  ( .D(n242), .CLK(clk), .RSTB(n180), .SETB(n179), .Q(
        Q_reg[3]) );
  DFFASRX1 \Q_reg_reg[2]  ( .D(n241), .CLK(clk), .RSTB(n178), .SETB(n177), .Q(
        Q_reg[2]) );
  DFFASRX1 \Q_reg_reg[1]  ( .D(n240), .CLK(clk), .RSTB(n176), .SETB(n175), .Q(
        Q_reg[1]) );
  AND2X1 U351 ( .IN1(n655), .IN2(n312), .Q(n310) );
  OA21X1 U353 ( .IN1(n538), .IN2(n539), .IN3(n659), .Q(n308) );
  OAI21X1 U354 ( .IN1(n539), .IN2(n620), .IN3(n540), .QN(n307) );
  AO21X1 U355 ( .IN1(n540), .IN2(n624), .IN3(n537), .Q(n306) );
  XNOR2X1 U356 ( .IN1(n622), .IN2(n537), .Q(n305) );
  AO22X1 U357 ( .IN1(n655), .IN2(Q_reg[1]), .IN3(n314), .IN4(n651), .Q(n304)
         );
  AO22X1 U358 ( .IN1(n314), .IN2(n655), .IN3(n651), .IN4(n623), .Q(n303) );
  OR2X1 U360 ( .IN1(n544), .IN2(n651), .Q(n542) );
  AO22X1 U362 ( .IN1(case_add[64]), .IN2(n647), .IN3(case_sub[64]), .IN4(n644), 
        .Q(n543) );
  AO221X1 U363 ( .IN1(n648), .IN2(Acc[30]), .IN3(case_sub[63]), .IN4(n644), 
        .IN5(n548), .Q(n300) );
  AO22X1 U364 ( .IN1(n652), .IN2(Acc[29]), .IN3(n647), .IN4(case_add[63]), .Q(
        n548) );
  AO221X1 U365 ( .IN1(n648), .IN2(Acc[29]), .IN3(case_sub[62]), .IN4(n644), 
        .IN5(n549), .Q(n299) );
  AO22X1 U366 ( .IN1(n653), .IN2(Acc[28]), .IN3(case_add[62]), .IN4(n647), .Q(
        n549) );
  AO221X1 U367 ( .IN1(n648), .IN2(Acc[28]), .IN3(case_sub[61]), .IN4(n644), 
        .IN5(n550), .Q(n298) );
  AO22X1 U368 ( .IN1(n652), .IN2(Acc[27]), .IN3(case_add[61]), .IN4(n647), .Q(
        n550) );
  AO221X1 U369 ( .IN1(n648), .IN2(Acc[27]), .IN3(case_sub[60]), .IN4(n644), 
        .IN5(n551), .Q(n297) );
  AO22X1 U370 ( .IN1(n652), .IN2(Acc[26]), .IN3(case_add[60]), .IN4(n647), .Q(
        n551) );
  AO221X1 U371 ( .IN1(n648), .IN2(Acc[26]), .IN3(case_sub[59]), .IN4(n644), 
        .IN5(n552), .Q(n296) );
  AO22X1 U372 ( .IN1(n653), .IN2(Acc[25]), .IN3(case_add[59]), .IN4(n647), .Q(
        n552) );
  AO221X1 U373 ( .IN1(n648), .IN2(Acc[25]), .IN3(case_sub[58]), .IN4(n644), 
        .IN5(n553), .Q(n295) );
  AO22X1 U374 ( .IN1(n652), .IN2(Acc[24]), .IN3(case_add[58]), .IN4(n647), .Q(
        n553) );
  AO221X1 U375 ( .IN1(n648), .IN2(Acc[24]), .IN3(case_sub[57]), .IN4(n644), 
        .IN5(n554), .Q(n294) );
  AO22X1 U376 ( .IN1(n653), .IN2(Acc[23]), .IN3(case_add[57]), .IN4(n647), .Q(
        n554) );
  AO221X1 U377 ( .IN1(n648), .IN2(Acc[23]), .IN3(case_sub[56]), .IN4(n643), 
        .IN5(n555), .Q(n293) );
  AO22X1 U378 ( .IN1(n653), .IN2(Acc[22]), .IN3(case_add[56]), .IN4(n646), .Q(
        n555) );
  AO221X1 U379 ( .IN1(n648), .IN2(Acc[22]), .IN3(case_sub[55]), .IN4(n643), 
        .IN5(n556), .Q(n292) );
  AO22X1 U380 ( .IN1(n653), .IN2(Acc[21]), .IN3(case_add[55]), .IN4(n646), .Q(
        n556) );
  AO221X1 U381 ( .IN1(n648), .IN2(Acc[21]), .IN3(case_sub[54]), .IN4(n643), 
        .IN5(n557), .Q(n291) );
  AO22X1 U382 ( .IN1(n653), .IN2(Acc[20]), .IN3(case_add[54]), .IN4(n646), .Q(
        n557) );
  AO221X1 U383 ( .IN1(n648), .IN2(Acc[20]), .IN3(case_sub[53]), .IN4(n643), 
        .IN5(n558), .Q(n290) );
  AO22X1 U384 ( .IN1(n653), .IN2(n668), .IN3(case_add[53]), .IN4(n646), .Q(
        n558) );
  AO221X1 U385 ( .IN1(n649), .IN2(n668), .IN3(case_sub[52]), .IN4(n643), .IN5(
        n559), .Q(n289) );
  AO22X1 U386 ( .IN1(n653), .IN2(Acc[18]), .IN3(case_add[52]), .IN4(n646), .Q(
        n559) );
  AO221X1 U387 ( .IN1(n649), .IN2(Acc[18]), .IN3(case_sub[51]), .IN4(n643), 
        .IN5(n560), .Q(n288) );
  AO22X1 U388 ( .IN1(n652), .IN2(Acc[17]), .IN3(case_add[51]), .IN4(n646), .Q(
        n560) );
  AO221X1 U389 ( .IN1(n649), .IN2(Acc[17]), .IN3(case_sub[50]), .IN4(n643), 
        .IN5(n561), .Q(n287) );
  AO22X1 U390 ( .IN1(n653), .IN2(Acc[16]), .IN3(case_add[50]), .IN4(n646), .Q(
        n561) );
  AO221X1 U391 ( .IN1(n649), .IN2(Acc[16]), .IN3(case_sub[49]), .IN4(n643), 
        .IN5(n562), .Q(n286) );
  AO22X1 U392 ( .IN1(n653), .IN2(n669), .IN3(case_add[49]), .IN4(n646), .Q(
        n562) );
  AO221X1 U393 ( .IN1(n649), .IN2(n669), .IN3(case_sub[48]), .IN4(n643), .IN5(
        n563), .Q(n285) );
  AO22X1 U394 ( .IN1(n653), .IN2(n670), .IN3(case_add[48]), .IN4(n646), .Q(
        n563) );
  AO221X1 U395 ( .IN1(n649), .IN2(n670), .IN3(case_sub[47]), .IN4(n643), .IN5(
        n564), .Q(n284) );
  AO22X1 U396 ( .IN1(n653), .IN2(n671), .IN3(case_add[47]), .IN4(n646), .Q(
        n564) );
  AO221X1 U397 ( .IN1(n649), .IN2(n671), .IN3(case_sub[46]), .IN4(n643), .IN5(
        n565), .Q(n283) );
  AO22X1 U398 ( .IN1(n653), .IN2(n672), .IN3(case_add[46]), .IN4(n646), .Q(
        n565) );
  AO221X1 U399 ( .IN1(n649), .IN2(n672), .IN3(case_sub[45]), .IN4(n643), .IN5(
        n566), .Q(n282) );
  AO22X1 U400 ( .IN1(n653), .IN2(Acc[11]), .IN3(case_add[45]), .IN4(n646), .Q(
        n566) );
  AO221X1 U401 ( .IN1(n649), .IN2(Acc[11]), .IN3(case_sub[44]), .IN4(n642), 
        .IN5(n567), .Q(n281) );
  AO22X1 U402 ( .IN1(n653), .IN2(n673), .IN3(case_add[44]), .IN4(n645), .Q(
        n567) );
  AO221X1 U403 ( .IN1(n649), .IN2(n673), .IN3(case_sub[43]), .IN4(n642), .IN5(
        n568), .Q(n280) );
  AO22X1 U404 ( .IN1(n653), .IN2(n674), .IN3(case_add[43]), .IN4(n645), .Q(
        n568) );
  AO221X1 U405 ( .IN1(n649), .IN2(n674), .IN3(case_sub[42]), .IN4(n642), .IN5(
        n569), .Q(n279) );
  AO22X1 U406 ( .IN1(n653), .IN2(n628), .IN3(case_add[42]), .IN4(n645), .Q(
        n569) );
  AO221X1 U407 ( .IN1(n649), .IN2(n628), .IN3(case_sub[41]), .IN4(n642), .IN5(
        n570), .Q(n278) );
  AO22X1 U408 ( .IN1(n653), .IN2(Acc[7]), .IN3(case_add[41]), .IN4(n645), .Q(
        n570) );
  AO221X1 U409 ( .IN1(n650), .IN2(Acc[7]), .IN3(case_sub[40]), .IN4(n642), 
        .IN5(n571), .Q(n277) );
  AO22X1 U410 ( .IN1(n653), .IN2(Acc[6]), .IN3(case_add[40]), .IN4(n645), .Q(
        n571) );
  AO221X1 U411 ( .IN1(n650), .IN2(Acc[6]), .IN3(case_sub[39]), .IN4(n642), 
        .IN5(n572), .Q(n276) );
  AO22X1 U412 ( .IN1(n653), .IN2(Acc[5]), .IN3(case_add[39]), .IN4(n645), .Q(
        n572) );
  AO221X1 U413 ( .IN1(n650), .IN2(Acc[5]), .IN3(case_sub[38]), .IN4(n642), 
        .IN5(n573), .Q(n275) );
  AO22X1 U414 ( .IN1(n653), .IN2(n627), .IN3(case_add[38]), .IN4(n645), .Q(
        n573) );
  AO221X1 U415 ( .IN1(n650), .IN2(n627), .IN3(case_sub[37]), .IN4(n642), .IN5(
        n574), .Q(n274) );
  AO22X1 U416 ( .IN1(n653), .IN2(n675), .IN3(case_add[37]), .IN4(n645), .Q(
        n574) );
  AO221X1 U417 ( .IN1(n650), .IN2(n675), .IN3(case_sub[36]), .IN4(n642), .IN5(
        n575), .Q(n273) );
  AO22X1 U418 ( .IN1(n653), .IN2(n626), .IN3(case_add[36]), .IN4(n645), .Q(
        n575) );
  AO221X1 U419 ( .IN1(n650), .IN2(n626), .IN3(case_sub[35]), .IN4(n642), .IN5(
        n576), .Q(n272) );
  AO22X1 U420 ( .IN1(n653), .IN2(n677), .IN3(case_add[35]), .IN4(n645), .Q(
        n576) );
  AO221X1 U421 ( .IN1(n650), .IN2(n677), .IN3(case_sub[34]), .IN4(n642), .IN5(
        n577), .Q(n271) );
  AO22X1 U422 ( .IN1(n652), .IN2(Acc[0]), .IN3(case_add[34]), .IN4(n645), .Q(
        n577) );
  AO221X1 U423 ( .IN1(n650), .IN2(Acc[0]), .IN3(case_sub[33]), .IN4(n642), 
        .IN5(n578), .Q(n270) );
  AO22X1 U424 ( .IN1(n652), .IN2(Q_reg[31]), .IN3(case_add[33]), .IN4(n645), 
        .Q(n578) );
  NOR3X0 U425 ( .IN1(n314), .IN2(n318), .IN3(n651), .QN(n546) );
  AND3X1 U426 ( .IN1(n314), .IN2(n659), .IN3(n318), .Q(n547) );
  AND2X1 U427 ( .IN1(n544), .IN2(n655), .Q(n545) );
  XNOR2X1 U428 ( .IN1(n314), .IN2(n623), .Q(n544) );
  AO22X1 U429 ( .IN1(n655), .IN2(Q_reg[31]), .IN3(n652), .IN4(Q_reg[30]), .Q(
        n269) );
  AO22X1 U430 ( .IN1(n655), .IN2(Q_reg[30]), .IN3(n652), .IN4(Q_reg[29]), .Q(
        n268) );
  AO22X1 U431 ( .IN1(n655), .IN2(Q_reg[29]), .IN3(n652), .IN4(Q_reg[28]), .Q(
        n267) );
  AO22X1 U432 ( .IN1(n656), .IN2(Q_reg[28]), .IN3(n652), .IN4(Q_reg[27]), .Q(
        n266) );
  AO22X1 U433 ( .IN1(n656), .IN2(Q_reg[27]), .IN3(n652), .IN4(Q_reg[26]), .Q(
        n265) );
  AO22X1 U434 ( .IN1(n656), .IN2(Q_reg[26]), .IN3(n652), .IN4(Q_reg[25]), .Q(
        n264) );
  AO22X1 U435 ( .IN1(n656), .IN2(Q_reg[25]), .IN3(n652), .IN4(Q_reg[24]), .Q(
        n263) );
  AO22X1 U436 ( .IN1(n656), .IN2(Q_reg[24]), .IN3(n652), .IN4(Q_reg[23]), .Q(
        n262) );
  AO22X1 U437 ( .IN1(n656), .IN2(Q_reg[23]), .IN3(n652), .IN4(Q_reg[22]), .Q(
        n261) );
  AO22X1 U438 ( .IN1(n656), .IN2(Q_reg[22]), .IN3(n652), .IN4(Q_reg[21]), .Q(
        n260) );
  AO22X1 U439 ( .IN1(n656), .IN2(Q_reg[21]), .IN3(n652), .IN4(Q_reg[20]), .Q(
        n259) );
  AO22X1 U440 ( .IN1(n657), .IN2(Q_reg[20]), .IN3(n652), .IN4(Q_reg[19]), .Q(
        n258) );
  AO22X1 U441 ( .IN1(n657), .IN2(Q_reg[19]), .IN3(n652), .IN4(Q_reg[18]), .Q(
        n257) );
  AO22X1 U442 ( .IN1(n657), .IN2(Q_reg[18]), .IN3(n652), .IN4(Q_reg[17]), .Q(
        n256) );
  AO22X1 U443 ( .IN1(n657), .IN2(Q_reg[17]), .IN3(n652), .IN4(Q_reg[16]), .Q(
        n255) );
  AO22X1 U444 ( .IN1(n657), .IN2(Q_reg[16]), .IN3(n651), .IN4(Q_reg[15]), .Q(
        n254) );
  AO22X1 U445 ( .IN1(n657), .IN2(Q_reg[15]), .IN3(n651), .IN4(Q_reg[14]), .Q(
        n253) );
  AO22X1 U446 ( .IN1(n657), .IN2(Q_reg[14]), .IN3(n651), .IN4(Q_reg[13]), .Q(
        n252) );
  AO22X1 U447 ( .IN1(n658), .IN2(Q_reg[13]), .IN3(n651), .IN4(Q_reg[12]), .Q(
        n251) );
  AO22X1 U448 ( .IN1(n658), .IN2(Q_reg[12]), .IN3(n651), .IN4(Q_reg[11]), .Q(
        n250) );
  AO22X1 U449 ( .IN1(n658), .IN2(Q_reg[11]), .IN3(n651), .IN4(Q_reg[10]), .Q(
        n249) );
  AO22X1 U450 ( .IN1(n658), .IN2(Q_reg[10]), .IN3(n651), .IN4(Q_reg[9]), .Q(
        n248) );
  AO22X1 U451 ( .IN1(n658), .IN2(Q_reg[9]), .IN3(n651), .IN4(Q_reg[8]), .Q(
        n247) );
  AO22X1 U452 ( .IN1(n658), .IN2(Q_reg[8]), .IN3(n651), .IN4(Q_reg[7]), .Q(
        n246) );
  AO22X1 U453 ( .IN1(n657), .IN2(Q_reg[7]), .IN3(n651), .IN4(Q_reg[6]), .Q(
        n245) );
  AO22X1 U454 ( .IN1(n658), .IN2(Q_reg[6]), .IN3(n651), .IN4(Q_reg[5]), .Q(
        n244) );
  AO22X1 U455 ( .IN1(n658), .IN2(Q_reg[5]), .IN3(n651), .IN4(Q_reg[4]), .Q(
        n243) );
  AO22X1 U456 ( .IN1(n659), .IN2(Q_reg[4]), .IN3(n651), .IN4(Q_reg[3]), .Q(
        n242) );
  AO22X1 U457 ( .IN1(n659), .IN2(Q_reg[3]), .IN3(n652), .IN4(Q_reg[2]), .Q(
        n241) );
  AO22X1 U458 ( .IN1(n655), .IN2(Q_reg[2]), .IN3(n651), .IN4(Q_reg[1]), .Q(
        n240) );
  AND2X1 U460 ( .IN1(n620), .IN2(n539), .Q(n541) );
  AND2X1 U461 ( .IN1(n315), .IN2(n312), .Q(n539) );
  OR2X1 U462 ( .IN1(n666), .IN2(Q[0]), .Q(n238) );
  OR2X1 U463 ( .IN1(n665), .IN2(Q[31]), .Q(n236) );
  OR2X1 U464 ( .IN1(n665), .IN2(Q[30]), .Q(n234) );
  OR2X1 U465 ( .IN1(n665), .IN2(Q[29]), .Q(n232) );
  OR2X1 U466 ( .IN1(n666), .IN2(Q[28]), .Q(n230) );
  OR2X1 U467 ( .IN1(n666), .IN2(Q[27]), .Q(n228) );
  OR2X1 U468 ( .IN1(n666), .IN2(Q[26]), .Q(n226) );
  OR2X1 U469 ( .IN1(n666), .IN2(Q[25]), .Q(n224) );
  OR2X1 U470 ( .IN1(n666), .IN2(Q[24]), .Q(n222) );
  OR2X1 U471 ( .IN1(n666), .IN2(Q[23]), .Q(n220) );
  OR2X1 U472 ( .IN1(n666), .IN2(Q[22]), .Q(n218) );
  OR2X1 U473 ( .IN1(n666), .IN2(Q[21]), .Q(n216) );
  OR2X1 U474 ( .IN1(n666), .IN2(Q[20]), .Q(n214) );
  OR2X1 U475 ( .IN1(n666), .IN2(Q[19]), .Q(n212) );
  OR2X1 U476 ( .IN1(n666), .IN2(Q[18]), .Q(n210) );
  OR2X1 U477 ( .IN1(n666), .IN2(Q[17]), .Q(n208) );
  OR2X1 U478 ( .IN1(n666), .IN2(Q[16]), .Q(n206) );
  OR2X1 U479 ( .IN1(n666), .IN2(Q[15]), .Q(n204) );
  OR2X1 U480 ( .IN1(n666), .IN2(Q[14]), .Q(n202) );
  OR2X1 U481 ( .IN1(n666), .IN2(Q[13]), .Q(n200) );
  OR2X1 U482 ( .IN1(n667), .IN2(Q[12]), .Q(n198) );
  OR2X1 U483 ( .IN1(n667), .IN2(Q[11]), .Q(n196) );
  OR2X1 U484 ( .IN1(n667), .IN2(Q[10]), .Q(n194) );
  OR2X1 U485 ( .IN1(n667), .IN2(Q[9]), .Q(n192) );
  OR2X1 U486 ( .IN1(n667), .IN2(Q[8]), .Q(n190) );
  OR2X1 U487 ( .IN1(n667), .IN2(Q[7]), .Q(n188) );
  OR2X1 U488 ( .IN1(n667), .IN2(Q[6]), .Q(n186) );
  OR2X1 U489 ( .IN1(n667), .IN2(Q[5]), .Q(n184) );
  OR2X1 U490 ( .IN1(n667), .IN2(Q[4]), .Q(n182) );
  OR2X1 U491 ( .IN1(n667), .IN2(Q[3]), .Q(n180) );
  OR2X1 U492 ( .IN1(n667), .IN2(Q[2]), .Q(n178) );
  OR2X1 U493 ( .IN1(n667), .IN2(Q[1]), .Q(n176) );
  BoothMultiplier_DW01_sub_1 sub_61 ( .A({Acc[31:20], n668, Acc[18:15], n670, 
        n671, n672, Acc[11:10], n674, n628, Acc[7:5], n627, n675, Acc[2], n677, 
        Acc[0]}), .B(M_reg), .CI(1'b0), .DIFF(case_sub) );
  BoothMultiplier_DW01_add_1 add_57 ( .A({Acc[31:21], n625, Acc[19:16], n669, 
        Acc[14:11], n673, Acc[9:3], n676, Acc[1:0]}), .B(M_reg), .CI(1'b0), 
        .SUM(case_add) );
  NAND3X0 U494 ( .IN1(n622), .IN2(n541), .IN3(n621), .QN(n536) );
  INVX0 U495 ( (n654), (n651) );
  INVX0 U496 ( (n654), (n652) );
  INVX0 U497 ( (n654), (n653) );
  NBUFFX2 U498 ( (n545), (n650) );
  NBUFFX2 U499 ( (n536), (n654) );
  NBUFFX2 U500 ( (n547), (n644) );
  NBUFFX2 U501 ( (n546), (n647) );
  NBUFFX2 U502 ( (n536), (n655) );
  NBUFFX2 U503 ( (n536), (n659) );
  NAND2X1 U504 ( .IN1(n541), .IN2(n654), .QN(n540) );
  NOR2X0 U505 ( .IN1(n540), .IN2(n624), .QN(n537) );
  AO221X1 U506 ( .IN1(n648), .IN2(Acc[31]), .IN3(n651), .IN4(Acc[30]), .IN5(
        n543), .Q(n301) );
  AO21X1 U507 ( .IN1(n542), .IN2(Acc[31]), .IN3(n543), .Q(n302) );
  NBUFFX2 U508 ( (n536), (n658) );
  NBUFFX2 U509 ( (n536), (n657) );
  NBUFFX2 U510 ( (n536), (n656) );
  NBUFFX2 U511 ( (n678), (n640) );
  NBUFFX2 U512 ( (n678), (n639) );
  NBUFFX2 U513 ( (n678), (n638) );
  NBUFFX2 U514 ( (n678), (n637) );
  NBUFFX2 U515 ( (n678), (n636) );
  NBUFFX2 U516 ( (n678), (n635) );
  NBUFFX2 U517 ( (n678), (n634) );
  NBUFFX2 U518 ( (n678), (n633) );
  NBUFFX2 U519 ( (n678), (n632) );
  NBUFFX2 U520 ( (n678), (n631) );
  NBUFFX2 U521 ( (n678), (n630) );
  NBUFFX2 U522 ( (n678), (n629) );
  NBUFFX2 U523 ( (n678), (n641) );
  INVX0 U524 ( (n153), (n671) );
  INVX0 U525 ( (n159), (n668) );
  INVX0 U526 ( (n152), (n672) );
  INVX0 U527 ( (n149), (n674) );
  INVX0 U528 ( (n141), (n677) );
  INVX0 U529 ( (n150), (n673) );
  INVX0 U530 ( (n155), (n669) );
  NBUFFX2 U531 ( (Acc[2]), (n626) );
  NOR2X0 U532 ( .IN1(n315), .IN2(n312), .QN(n538) );
  INVX0 U533 ( (oRst), (n678) );
  NBUFFX2 U534 ( (rst), (n662) );
  NBUFFX2 U535 ( (rst), (n660) );
  NBUFFX2 U536 ( (rst), (n661) );
  NBUFFX2 U537 ( (rst), (n663) );
  NAND2X1 U538 ( .IN1(Q[25]), .IN2(n662), .QN(n223) );
  NAND2X1 U539 ( .IN1(Q[26]), .IN2(n662), .QN(n225) );
  NAND2X1 U540 ( .IN1(Q[27]), .IN2(n662), .QN(n227) );
  NAND2X1 U541 ( .IN1(Q[28]), .IN2(n662), .QN(n229) );
  NAND2X1 U542 ( .IN1(Q[29]), .IN2(n662), .QN(n231) );
  NAND2X1 U543 ( .IN1(Q[30]), .IN2(n662), .QN(n233) );
  NAND2X1 U544 ( .IN1(Q[31]), .IN2(n662), .QN(n235) );
  NAND2X1 U545 ( .IN1(Q[0]), .IN2(n662), .QN(n237) );
  NAND2X1 U546 ( .IN1(Q[1]), .IN2(n660), .QN(n175) );
  NAND2X1 U547 ( .IN1(Q[2]), .IN2(n660), .QN(n177) );
  NAND2X1 U548 ( .IN1(Q[3]), .IN2(n660), .QN(n179) );
  NAND2X1 U549 ( .IN1(Q[4]), .IN2(n660), .QN(n181) );
  NAND2X1 U550 ( .IN1(Q[5]), .IN2(n660), .QN(n183) );
  NAND2X1 U551 ( .IN1(Q[6]), .IN2(n660), .QN(n185) );
  NAND2X1 U552 ( .IN1(Q[7]), .IN2(n660), .QN(n187) );
  NAND2X1 U553 ( .IN1(Q[8]), .IN2(n660), .QN(n189) );
  NAND2X1 U554 ( .IN1(Q[9]), .IN2(n660), .QN(n191) );
  NAND2X1 U555 ( .IN1(Q[10]), .IN2(n660), .QN(n193) );
  NAND2X1 U556 ( .IN1(Q[11]), .IN2(n660), .QN(n195) );
  NAND2X1 U557 ( .IN1(Q[12]), .IN2(n660), .QN(n197) );
  NAND2X1 U558 ( .IN1(Q[13]), .IN2(n661), .QN(n199) );
  NAND2X1 U559 ( .IN1(Q[14]), .IN2(n661), .QN(n201) );
  NAND2X1 U560 ( .IN1(Q[15]), .IN2(n661), .QN(n203) );
  NAND2X1 U561 ( .IN1(Q[16]), .IN2(n661), .QN(n205) );
  NAND2X1 U562 ( .IN1(Q[17]), .IN2(n661), .QN(n207) );
  NAND2X1 U563 ( .IN1(Q[18]), .IN2(n661), .QN(n209) );
  NAND2X1 U564 ( .IN1(Q[19]), .IN2(n661), .QN(n211) );
  NAND2X1 U565 ( .IN1(Q[20]), .IN2(n661), .QN(n213) );
  NAND2X1 U566 ( .IN1(Q[21]), .IN2(n661), .QN(n215) );
  NAND2X1 U567 ( .IN1(Q[22]), .IN2(n661), .QN(n217) );
  NAND2X1 U568 ( .IN1(Q[23]), .IN2(n661), .QN(n219) );
  NAND2X1 U569 ( .IN1(Q[24]), .IN2(n661), .QN(n221) );
  INVX0 U570 ( (n143), (n675) );
  INVX0 U571 ( (n160), (n625) );
  INVX0 U572 ( (n618), (n627) );
  INVX0 U573 ( (n154), (n670) );
  INVX0 U574 ( (n148), (n628) );
  INVX0 U575 ( (n142), (n676) );
  NBUFFX2 U576 ( (n547), (n642) );
  NBUFFX2 U577 ( (n547), (n643) );
  NBUFFX2 U578 ( (n546), (n645) );
  NBUFFX2 U579 ( (n546), (n646) );
  NBUFFX2 U580 ( (n545), (n648) );
  NBUFFX2 U581 ( (n545), (n649) );
  INVX0 U582 ( (n662), (n664) );
  INVX0 U583 ( (n662), (n665) );
  INVX0 U584 ( (n662), (n666) );
  INVX0 U585 ( (n662), (n667) );
endmodule
