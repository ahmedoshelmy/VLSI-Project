
module BoothMultiplier_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391;

  AND2X1 U3 ( .IN1(n213), .IN2(n206), .Q(n55) );
  AND2X1 U4 ( .IN1(n213), .IN2(n221), .Q(n48) );
  AND2X1 U5 ( .IN1(n221), .IN2(n229), .Q(n46) );
  AND2X1 U6 ( .IN1(n60), .IN2(n10), .Q(n24) );
  AND2X1 U7 ( .IN1(n199), .IN2(n192), .Q(n35) );
  XOR3X1 U8 ( .IN1(n175), .IN2(B[28]), .IN3(n66), .Q(DIFF[28]) );
  AND2X1 U9 ( .IN1(n210), .IN2(n211), .Q(n1) );
  AND2X1 U10 ( .IN1(n196), .IN2(n197), .Q(n2) );
  AND2X1 U11 ( .IN1(n190), .IN2(n191), .Q(n3) );
  NOR2X0 U12 ( .IN1(n13), .IN2(n14), .QN(n4) );
  NOR2X0 U13 ( .IN1(n27), .IN2(n28), .QN(n5) );
  NAND2X1 U14 ( .IN1(B[2]), .IN2(n376), .QN(n153) );
  NOR2X0 U15 ( .IN1(n6), .IN2(n7), .QN(n60) );
  NAND2X1 U16 ( .IN1(n58), .IN2(n56), .QN(n6) );
  AND2X1 U17 ( .IN1(n228), .IN2(n57), .Q(n7) );
  OR2X1 U18 ( .IN1(n8), .IN2(n9), .Q(n66) );
  NAND2X1 U19 ( .IN1(n23), .IN2(n67), .QN(n8) );
  NAND2X0 U20 ( .IN1(n60), .IN2(n11), .QN(n9) );
  AND2X1 U21 ( .IN1(n61), .IN2(n4), .Q(n10) );
  AND2X1 U22 ( .IN1(n61), .IN2(n12), .Q(n11) );
  INVX0 U23 ( .INP(n14), .ZN(n12) );
  INVX0 U24 ( .INP(n67), .ZN(n13) );
  NOR2X0 U25 ( .IN1(n64), .IN2(n204), .QN(n14) );
  NAND2X0 U26 ( .IN1(n205), .IN2(n18), .QN(n15) );
  NAND2X0 U27 ( .IN1(n15), .IN2(n16), .QN(n191) );
  OR2X1 U28 ( .IN1(n17), .IN2(n35), .Q(n16) );
  INVX0 U29 ( .INP(n33), .ZN(n17) );
  AND2X1 U30 ( .IN1(n204), .IN2(n33), .Q(n18) );
  NAND2X1 U31 ( .IN1(n227), .IN2(n22), .QN(n19) );
  NAND2X0 U32 ( .IN1(n19), .IN2(n20), .QN(n52) );
  OR2X1 U33 ( .IN1(n21), .IN2(n38), .Q(n20) );
  INVX0 U34 ( .INP(n36), .ZN(n21) );
  AND2X1 U35 ( .IN1(n226), .IN2(n36), .Q(n22) );
  NAND2X1 U36 ( .IN1(n204), .IN2(n205), .QN(n198) );
  AND2X1 U37 ( .IN1(n76), .IN2(n5), .Q(n23) );
  AND2X1 U38 ( .IN1(n24), .IN2(n25), .Q(n178) );
  AND2X1 U39 ( .IN1(n26), .IN2(n76), .Q(n25) );
  INVX0 U40 ( .INP(n28), .ZN(n26) );
  INVX0 U41 ( .INP(n177), .ZN(n27) );
  NOR2X0 U42 ( .IN1(n89), .IN2(n183), .QN(n28) );
  NAND2X0 U43 ( .IN1(n178), .IN2(n32), .QN(n29) );
  AND2X1 U44 ( .IN1(n29), .IN2(n30), .Q(n155) );
  OR2X1 U45 ( .IN1(n31), .IN2(n43), .Q(n30) );
  INVX0 U46 ( .INP(n156), .ZN(n31) );
  AND2X1 U47 ( .IN1(n45), .IN2(n156), .Q(n32) );
  OR2X1 U48 ( .IN1(n34), .IN2(n196), .Q(n33) );
  INVX0 U49 ( .INP(n192), .ZN(n34) );
  OR2X1 U50 ( .IN1(n37), .IN2(n218), .Q(n36) );
  INVX0 U51 ( .INP(n55), .ZN(n37) );
  AND2X1 U52 ( .IN1(n221), .IN2(n55), .Q(n38) );
  NAND2X0 U53 ( .IN1(n66), .IN2(n42), .QN(n39) );
  AND2X1 U54 ( .IN1(n39), .IN2(n40), .Q(n162) );
  OR2X1 U55 ( .IN1(n41), .IN2(n172), .Q(n40) );
  INVX0 U56 ( .INP(n163), .ZN(n41) );
  AND2X1 U57 ( .IN1(n174), .IN2(n163), .Q(n42) );
  OR2X1 U58 ( .IN1(n44), .IN2(n49), .Q(n43) );
  INVX0 U59 ( .INP(n73), .ZN(n44) );
  AND2X1 U60 ( .IN1(n51), .IN2(n73), .Q(n45) );
  NAND2X0 U61 ( .IN1(n65), .IN2(n48), .QN(n47) );
  OR2X1 U62 ( .IN1(n50), .IN2(n72), .Q(n49) );
  INVX0 U63 ( .INP(n70), .ZN(n50) );
  AND2X1 U64 ( .IN1(n177), .IN2(n70), .Q(n51) );
  NAND2X0 U65 ( .IN1(B[27]), .IN2(n181), .QN(n179) );
  AND4X4 U66 ( .IN1(n280), .IN2(n277), .IN3(n279), .IN4(n278), .Q(n91) );
  AND2X1 U67 ( .IN1(n52), .IN2(n53), .Q(n205) );
  OR2X1 U68 ( .IN1(n54), .IN2(n210), .Q(n53) );
  INVX0 U69 ( .INP(n206), .ZN(n54) );
  OR2X1 U70 ( .IN1(n47), .IN2(n226), .Q(n56) );
  AND2X1 U71 ( .IN1(n63), .IN2(n46), .Q(n57) );
  OR2X1 U72 ( .IN1(n59), .IN2(n218), .Q(n58) );
  INVX0 U73 ( .INP(n63), .ZN(n59) );
  OR2X1 U74 ( .IN1(n62), .IN2(n210), .Q(n61) );
  INVX0 U75 ( .INP(n65), .ZN(n62) );
  AND2X1 U76 ( .IN1(n213), .IN2(n65), .Q(n63) );
  INVX0 U77 ( .INP(n69), .ZN(n64) );
  AND2X1 U78 ( .IN1(n206), .IN2(n69), .Q(n65) );
  OR2X1 U79 ( .IN1(n68), .IN2(n196), .Q(n67) );
  INVX0 U80 ( .INP(n78), .ZN(n68) );
  AND2X1 U81 ( .IN1(n199), .IN2(n78), .Q(n69) );
  OR2X1 U82 ( .IN1(n71), .IN2(n172), .Q(n70) );
  INVX0 U83 ( .INP(n75), .ZN(n71) );
  AND2X1 U84 ( .IN1(n174), .IN2(n75), .Q(n72) );
  NAND2X0 U85 ( .IN1(n255), .IN2(n254), .QN(n237) );
  NAND2X0 U86 ( .IN1(n254), .IN2(n252), .QN(n259) );
  NAND2X0 U87 ( .IN1(n238), .IN2(n241), .QN(n248) );
  NAND2X0 U88 ( .IN1(n229), .IN2(n226), .QN(n230) );
  NAND2X0 U89 ( .IN1(n218), .IN2(n221), .QN(n223) );
  NAND2X0 U90 ( .IN1(B[18]), .IN2(n268), .QN(n254) );
  NAND2X0 U91 ( .IN1(A[14]), .IN2(n327), .QN(n287) );
  NAND2X0 U92 ( .IN1(B[19]), .IN2(n258), .QN(n238) );
  NAND2X0 U93 ( .IN1(B[21]), .IN2(n224), .QN(n221) );
  NAND2X0 U94 ( .IN1(B[22]), .IN2(n216), .QN(n213) );
  NAND2X0 U95 ( .IN1(B[20]), .IN2(n243), .QN(n229) );
  OR2X1 U96 ( .IN1(n74), .IN2(n161), .Q(n73) );
  INVX0 U97 ( .INP(n157), .ZN(n74) );
  AND2X1 U98 ( .IN1(n163), .IN2(n157), .Q(n75) );
  OR2X1 U99 ( .IN1(n77), .IN2(n190), .Q(n76) );
  INVX0 U100 ( .INP(n90), .ZN(n77) );
  AND2X1 U101 ( .IN1(n192), .IN2(n90), .Q(n78) );
  INVX0 U102 ( .INP(n123), .ZN(n122) );
  NOR2X0 U103 ( .IN1(n313), .IN2(n314), .QN(n312) );
  NOR2X0 U104 ( .IN1(n306), .IN2(n307), .QN(n304) );
  INVX0 U105 ( .INP(n297), .ZN(n307) );
  NAND2X0 U106 ( .IN1(n360), .IN2(n361), .QN(n123) );
  NOR2X0 U107 ( .IN1(n91), .IN2(n256), .QN(n261) );
  NOR2X0 U108 ( .IN1(n91), .IN2(n237), .QN(n250) );
  INVX0 U109 ( .INP(n131), .ZN(n133) );
  INVX0 U110 ( .INP(n355), .ZN(n357) );
  INVX0 U111 ( .INP(n323), .ZN(n324) );
  INVX0 U112 ( .INP(n118), .ZN(n117) );
  INVX0 U113 ( .INP(n329), .ZN(n330) );
  INVX0 U114 ( .INP(n137), .ZN(n140) );
  INVX0 U115 ( .INP(n335), .ZN(n338) );
  INVX0 U116 ( .INP(n170), .ZN(n244) );
  INVX0 U117 ( .INP(n144), .ZN(n146) );
  NOR2X0 U118 ( .IN1(n168), .IN2(n374), .QN(n371) );
  AND2X1 U119 ( .IN1(n99), .IN2(B[10]), .Q(n102) );
  INVX0 U120 ( .INP(n241), .ZN(n239) );
  NAND2X0 U121 ( .IN1(n266), .IN2(n265), .QN(n256) );
  NOR2X0 U122 ( .IN1(n289), .IN2(n290), .QN(n285) );
  NOR2X0 U123 ( .IN1(n111), .IN2(n287), .QN(n286) );
  INVX0 U124 ( .INP(n256), .ZN(n255) );
  NOR2X0 U125 ( .IN1(n371), .IN2(n372), .QN(n364) );
  INVX0 U126 ( .INP(n149), .ZN(n366) );
  AND2X1 U127 ( .IN1(n240), .IN2(n238), .Q(n79) );
  NOR2X0 U128 ( .IN1(n236), .IN2(n237), .QN(n234) );
  INVX0 U129 ( .INP(n238), .ZN(n236) );
  INVX0 U130 ( .INP(n293), .ZN(n292) );
  NAND2X0 U131 ( .IN1(n119), .IN2(n118), .QN(n358) );
  AND2X1 U132 ( .IN1(n183), .IN2(n184), .Q(n80) );
  NOR2X0 U133 ( .IN1(n91), .IN2(n272), .QN(n271) );
  INVX0 U134 ( .INP(n266), .ZN(n272) );
  NAND2X0 U135 ( .IN1(n293), .IN2(n334), .QN(n329) );
  NAND2X1 U136 ( .IN1(n335), .IN2(n336), .QN(n334) );
  OR2X1 U137 ( .IN1(n311), .IN2(n81), .Q(n144) );
  AND2X1 U138 ( .IN1(n106), .IN2(n110), .Q(n81) );
  NAND2X0 U139 ( .IN1(n289), .IN2(n328), .QN(n323) );
  NAND2X0 U140 ( .IN1(n329), .IN2(n316), .QN(n328) );
  NAND2X0 U141 ( .IN1(n339), .IN2(n340), .QN(n335) );
  NAND2X0 U142 ( .IN1(n168), .IN2(n169), .QN(n152) );
  NAND2X1 U143 ( .IN1(n152), .IN2(n153), .QN(n151) );
  NAND2X1 U144 ( .IN1(n125), .IN2(n359), .QN(n118) );
  NAND2X0 U145 ( .IN1(n93), .IN2(n123), .QN(n359) );
  NAND2X1 U146 ( .IN1(n141), .IN2(n142), .QN(n137) );
  NAND2X0 U147 ( .IN1(n143), .IN2(n144), .QN(n142) );
  NAND2X0 U148 ( .IN1(n129), .IN2(n130), .QN(n126) );
  NAND2X0 U149 ( .IN1(n287), .IN2(n322), .QN(n319) );
  NAND2X1 U150 ( .IN1(n246), .IN2(n104), .QN(n170) );
  AND2X1 U151 ( .IN1(n296), .IN2(n348), .Q(n82) );
  AND2X1 U152 ( .IN1(n150), .IN2(n153), .Q(n167) );
  NAND2X0 U153 ( .IN1(n289), .IN2(n316), .QN(n331) );
  NAND2X0 U154 ( .IN1(n143), .IN2(n141), .QN(n145) );
  NAND2X1 U155 ( .IN1(n93), .IN2(n125), .QN(n121) );
  NAND2X0 U156 ( .IN1(n336), .IN2(n293), .QN(n337) );
  AND2X1 U157 ( .IN1(n127), .IN2(n128), .Q(n83) );
  NAND2X0 U158 ( .IN1(n265), .IN2(n263), .QN(n269) );
  NAND2X1 U159 ( .IN1(n177), .IN2(n179), .QN(n180) );
  NAND2X1 U160 ( .IN1(n183), .IN2(n186), .QN(n187) );
  AND2X1 U161 ( .IN1(n106), .IN2(n149), .Q(n84) );
  NAND2X1 U162 ( .IN1(n210), .IN2(n213), .QN(n215) );
  NAND2X1 U163 ( .IN1(n204), .IN2(n206), .QN(n207) );
  NAND2X1 U164 ( .IN1(n196), .IN2(n199), .QN(n201) );
  NAND2X1 U165 ( .IN1(n190), .IN2(n192), .QN(n193) );
  AND2X1 U166 ( .IN1(n288), .IN2(n278), .Q(n85) );
  INVX0 U167 ( .INP(A[16]), .ZN(n318) );
  INVX0 U168 ( .INP(B[7]), .ZN(n386) );
  INVX0 U169 ( .INP(A[17]), .ZN(n275) );
  INVX0 U170 ( .INP(A[7]), .ZN(n381) );
  NAND2X1 U171 ( .IN1(A[30]), .IN2(n160), .QN(n156) );
  INVX0 U172 ( .INP(B[30]), .ZN(n160) );
  NAND2X1 U173 ( .IN1(A[29]), .IN2(n166), .QN(n161) );
  INVX0 U174 ( .INP(B[29]), .ZN(n166) );
  NAND2X1 U175 ( .IN1(A[28]), .IN2(n176), .QN(n172) );
  INVX0 U176 ( .INP(B[28]), .ZN(n176) );
  AND2X1 U177 ( .IN1(B[3]), .IN2(n375), .Q(n86) );
  INVX0 U178 ( .INP(A[18]), .ZN(n268) );
  XOR3X1 U179 ( .IN1(n165), .IN2(B[29]), .IN3(n164), .Q(DIFF[29]) );
  INVX0 U180 ( .INP(A[19]), .ZN(n258) );
  NAND2X0 U181 ( .IN1(A[18]), .IN2(n267), .QN(n252) );
  INVX0 U182 ( .INP(B[18]), .ZN(n267) );
  XOR3X1 U183 ( .IN1(n159), .IN2(B[30]), .IN3(n158), .Q(DIFF[30]) );
  NAND2X0 U184 ( .IN1(A[17]), .IN2(n274), .QN(n263) );
  INVX0 U185 ( .INP(B[17]), .ZN(n274) );
  NOR2X0 U186 ( .IN1(n87), .IN2(n88), .QN(n367) );
  NAND3X0 U187 ( .IN1(A[0]), .IN2(n171), .IN3(n153), .QN(n87) );
  NAND2X0 U188 ( .IN1(n106), .IN2(n368), .QN(n88) );
  INVX0 U189 ( .INP(B[8]), .ZN(n346) );
  INVX0 U190 ( .INP(B[0]), .ZN(n368) );
  NAND2X0 U191 ( .IN1(A[15]), .IN2(n320), .QN(n278) );
  NAND2X1 U192 ( .IN1(A[26]), .IN2(n189), .QN(n183) );
  INVX0 U193 ( .INP(B[26]), .ZN(n189) );
  INVX0 U194 ( .INP(A[27]), .ZN(n181) );
  NAND2X0 U195 ( .IN1(A[19]), .IN2(n257), .QN(n241) );
  INVX0 U196 ( .INP(B[19]), .ZN(n257) );
  NAND2X1 U197 ( .IN1(B[26]), .IN2(n188), .QN(n186) );
  INVX0 U198 ( .INP(A[26]), .ZN(n188) );
  NAND2X1 U199 ( .IN1(n96), .IN2(n246), .QN(DIFF[0]) );
  NAND2X0 U200 ( .IN1(A[20]), .IN2(n242), .QN(n226) );
  INVX0 U201 ( .INP(B[20]), .ZN(n242) );
  NAND2X1 U202 ( .IN1(A[23]), .IN2(n209), .QN(n204) );
  INVX0 U203 ( .INP(B[23]), .ZN(n209) );
  NAND2X0 U204 ( .IN1(A[21]), .IN2(n225), .QN(n218) );
  INVX0 U205 ( .INP(B[21]), .ZN(n225) );
  NAND2X0 U206 ( .IN1(A[22]), .IN2(n217), .QN(n210) );
  INVX0 U207 ( .INP(B[22]), .ZN(n217) );
  NAND2X1 U208 ( .IN1(A[24]), .IN2(n203), .QN(n196) );
  INVX0 U209 ( .INP(B[24]), .ZN(n203) );
  NAND2X1 U210 ( .IN1(A[25]), .IN2(n195), .QN(n190) );
  INVX0 U211 ( .INP(B[25]), .ZN(n195) );
  NAND2X1 U212 ( .IN1(A[27]), .IN2(n182), .QN(n177) );
  INVX0 U213 ( .INP(B[27]), .ZN(n182) );
  NAND2X1 U214 ( .IN1(B[23]), .IN2(n208), .QN(n206) );
  INVX0 U215 ( .INP(A[23]), .ZN(n208) );
  INVX0 U216 ( .INP(A[21]), .ZN(n224) );
  INVX0 U217 ( .INP(A[22]), .ZN(n216) );
  NAND2X1 U218 ( .IN1(B[24]), .IN2(n202), .QN(n199) );
  INVX0 U219 ( .INP(A[24]), .ZN(n202) );
  NAND2X1 U220 ( .IN1(B[25]), .IN2(n194), .QN(n192) );
  INVX0 U221 ( .INP(A[25]), .ZN(n194) );
  INVX0 U222 ( .INP(A[20]), .ZN(n243) );
  INVX0 U223 ( .INP(A[28]), .ZN(n175) );
  INVX0 U224 ( .INP(A[29]), .ZN(n165) );
  INVX0 U225 ( .INP(A[30]), .ZN(n159) );
  NAND2X1 U226 ( .IN1(B[28]), .IN2(n175), .QN(n174) );
  NAND2X1 U227 ( .IN1(B[29]), .IN2(n165), .QN(n163) );
  NAND2X1 U228 ( .IN1(B[30]), .IN2(n159), .QN(n157) );
  INVX0 U229 ( .INP(n220), .ZN(n222) );
  INVX0 U230 ( .INP(n212), .ZN(n214) );
  INVX0 U231 ( .INP(n179), .ZN(n89) );
  AND2X1 U232 ( .IN1(n186), .IN2(n179), .Q(n90) );
  NAND2X0 U233 ( .IN1(n311), .IN2(n312), .QN(n277) );
  INVX0 U234 ( .INP(A[31]), .ZN(n154) );
  INVX0 U235 ( .INP(A[6]), .ZN(n92) );
  NAND2X0 U236 ( .IN1(B[8]), .IN2(n387), .QN(n93) );
  NAND2X0 U237 ( .IN1(B[8]), .IN2(n387), .QN(n124) );
  INVX0 U238 ( .INP(A[8]), .ZN(n387) );
  AND3X1 U239 ( .IN1(n291), .IN2(n288), .IN3(n316), .Q(n94) );
  AND2X1 U240 ( .IN1(B[2]), .IN2(n376), .Q(n95) );
  NAND2X0 U241 ( .IN1(n385), .IN2(A[6]), .QN(n129) );
  NAND2X0 U242 ( .IN1(n135), .IN2(n136), .QN(n131) );
  NAND2X0 U243 ( .IN1(B[0]), .IN2(n391), .QN(n96) );
  NOR2X0 U244 ( .IN1(n97), .IN2(n98), .QN(n343) );
  NAND2X0 U245 ( .IN1(n348), .IN2(n349), .QN(n97) );
  NOR2X0 U246 ( .IN1(n102), .IN2(n120), .QN(n98) );
  INVX0 U247 ( .INP(A[14]), .ZN(n326) );
  INVX0 U248 ( .INP(A[10]), .ZN(n99) );
  NAND2X0 U249 ( .IN1(n253), .IN2(n254), .QN(n251) );
  NOR2X0 U250 ( .IN1(n261), .IN2(n253), .QN(n260) );
  NAND2X0 U251 ( .IN1(n262), .IN2(n263), .QN(n253) );
  INVX0 U252 ( .INP(B[4]), .ZN(n147) );
  NAND2X0 U253 ( .IN1(A[11]), .IN2(n352), .QN(n348) );
  NOR2X0 U254 ( .IN1(A[6]), .IN2(n385), .QN(n100) );
  NAND2X0 U255 ( .IN1(n170), .IN2(n171), .QN(n169) );
  NAND2X0 U256 ( .IN1(n168), .IN2(n171), .QN(n245) );
  NAND2X1 U257 ( .IN1(n150), .IN2(n151), .QN(n148) );
  NOR2X0 U258 ( .IN1(n86), .IN2(n150), .QN(n372) );
  NAND2X0 U259 ( .IN1(A[2]), .IN2(n373), .QN(n150) );
  NAND2X0 U260 ( .IN1(n92), .IN2(B[6]), .QN(n101) );
  INVX0 U261 ( .INP(B[1]), .ZN(n377) );
  INVX0 U262 ( .INP(B[10]), .ZN(n390) );
  NAND2X0 U263 ( .IN1(n124), .IN2(n119), .QN(n103) );
  NAND2X0 U264 ( .IN1(n349), .IN2(n354), .QN(n351) );
  NAND2X0 U265 ( .IN1(n390), .IN2(A[10]), .QN(n349) );
  NAND2X0 U266 ( .IN1(A[7]), .IN2(n386), .QN(n128) );
  NAND2X0 U267 ( .IN1(A[5]), .IN2(n384), .QN(n135) );
  INVX0 U268 ( .INP(n96), .ZN(n104) );
  NAND2X0 U269 ( .IN1(B[0]), .IN2(n391), .QN(n247) );
  AND4X1 U270 ( .IN1(n101), .IN2(n138), .IN3(A[4]), .IN4(n147), .Q(n105) );
  NAND2X0 U271 ( .IN1(B[3]), .IN2(n375), .QN(n106) );
  INVX0 U272 ( .INP(B[3]), .ZN(n370) );
  INVX0 U273 ( .INP(A[9]), .ZN(n388) );
  NAND2X0 U274 ( .IN1(n283), .IN2(n284), .QN(n282) );
  NOR2X0 U275 ( .IN1(n285), .IN2(n286), .QN(n284) );
  INVX0 U276 ( .INP(B[13]), .ZN(n333) );
  NAND2X1 U277 ( .IN1(B[13]), .IN2(n332), .QN(n316) );
  NAND2X0 U278 ( .IN1(n297), .IN2(n310), .QN(n314) );
  NAND2X0 U279 ( .IN1(n310), .IN2(n144), .QN(n361) );
  NOR2X0 U280 ( .IN1(n378), .IN2(n379), .QN(n310) );
  INVX0 U281 ( .INP(B[2]), .ZN(n373) );
  INVX0 U282 ( .INP(A[12]), .ZN(n315) );
  NAND2X1 U283 ( .IN1(A[12]), .IN2(n350), .QN(n293) );
  NAND2X0 U284 ( .IN1(n96), .IN2(n171), .QN(n107) );
  NAND2X0 U285 ( .IN1(n119), .IN2(n120), .QN(n116) );
  NAND2X0 U286 ( .IN1(n120), .IN2(n358), .QN(n355) );
  NAND2X0 U287 ( .IN1(A[9]), .IN2(n389), .QN(n120) );
  NOR2X0 U288 ( .IN1(n341), .IN2(n342), .QN(n108) );
  NOR2X0 U289 ( .IN1(n103), .IN2(n342), .QN(n303) );
  NAND2X0 U290 ( .IN1(n124), .IN2(n119), .QN(n341) );
  NAND2X1 U291 ( .IN1(n364), .IN2(n365), .QN(n311) );
  NOR2X0 U292 ( .IN1(n366), .IN2(n367), .QN(n365) );
  INVX0 U293 ( .INP(A[2]), .ZN(n376) );
  NAND2X0 U294 ( .IN1(B[5]), .IN2(n382), .QN(n109) );
  INVX0 U295 ( .INP(A[5]), .ZN(n382) );
  NAND2X1 U296 ( .IN1(B[4]), .IN2(n380), .QN(n143) );
  INVX0 U297 ( .INP(B[12]), .ZN(n350) );
  NAND2X1 U298 ( .IN1(B[12]), .IN2(n315), .QN(n297) );
  NAND2X0 U299 ( .IN1(n292), .IN2(n94), .QN(n283) );
  NAND2X0 U300 ( .IN1(n94), .IN2(n296), .QN(n295) );
  NOR2X0 U301 ( .IN1(n95), .IN2(n107), .QN(n110) );
  NAND2X0 U302 ( .IN1(n247), .IN2(n171), .QN(n363) );
  NOR2X0 U303 ( .IN1(n264), .IN2(n271), .QN(n270) );
  NAND2X0 U304 ( .IN1(n264), .IN2(n265), .QN(n262) );
  INVX0 U305 ( .INP(n273), .ZN(n264) );
  NAND2X0 U306 ( .IN1(n266), .IN2(n273), .QN(n276) );
  AND2X1 U307 ( .IN1(B[15]), .IN2(n321), .Q(n111) );
  INVX0 U308 ( .INP(A[15]), .ZN(n321) );
  NOR2X0 U309 ( .IN1(n100), .IN2(n135), .QN(n383) );
  NAND2X0 U310 ( .IN1(n377), .IN2(A[1]), .QN(n168) );
  INVX0 U311 ( .INP(A[1]), .ZN(n369) );
  INVX0 U312 ( .INP(n127), .ZN(n306) );
  NAND2X0 U313 ( .IN1(n153), .IN2(n106), .QN(n374) );
  NAND2X0 U314 ( .IN1(n137), .IN2(n109), .QN(n136) );
  NAND2X0 U315 ( .IN1(n109), .IN2(n135), .QN(n139) );
  NAND2X0 U316 ( .IN1(n143), .IN2(n109), .QN(n378) );
  NAND2X0 U317 ( .IN1(B[5]), .IN2(n382), .QN(n138) );
  NAND2X0 U318 ( .IN1(n291), .IN2(n288), .QN(n290) );
  NAND2X0 U319 ( .IN1(n323), .IN2(n291), .QN(n322) );
  NAND2X0 U320 ( .IN1(n287), .IN2(n291), .QN(n325) );
  NAND2X0 U321 ( .IN1(B[14]), .IN2(n326), .QN(n291) );
  NAND2X0 U322 ( .IN1(A[13]), .IN2(n333), .QN(n289) );
  INVX0 U323 ( .INP(A[13]), .ZN(n332) );
  NAND2X0 U324 ( .IN1(A[16]), .IN2(n317), .QN(n273) );
  NAND2X0 U325 ( .IN1(B[16]), .IN2(n318), .QN(n266) );
  INVX0 U326 ( .INP(A[4]), .ZN(n380) );
  NAND2X0 U327 ( .IN1(A[4]), .IN2(n147), .QN(n141) );
  NAND2X0 U328 ( .IN1(n112), .IN2(n113), .QN(n305) );
  AND2X1 U329 ( .IN1(n128), .IN2(n129), .Q(n112) );
  NOR2X0 U330 ( .IN1(n383), .IN2(n105), .QN(n113) );
  INVX0 U331 ( .INP(B[16]), .ZN(n317) );
  NAND2X0 U332 ( .IN1(n343), .IN2(n344), .QN(n114) );
  AND2X1 U333 ( .IN1(n106), .IN2(n362), .Q(n115) );
  NOR2X0 U334 ( .IN1(n363), .IN2(n95), .QN(n362) );
  INVX0 U335 ( .INP(B[9]), .ZN(n389) );
  NAND2X1 U336 ( .IN1(B[9]), .IN2(n388), .QN(n119) );
  NAND2X1 U337 ( .IN1(B[17]), .IN2(n275), .QN(n265) );
  INVX0 U338 ( .INP(B[11]), .ZN(n352) );
  NAND2X1 U339 ( .IN1(B[11]), .IN2(n353), .QN(n296) );
  NOR2X0 U340 ( .IN1(n301), .IN2(n302), .QN(n300) );
  NAND2X0 U341 ( .IN1(n303), .IN2(n94), .QN(n302) );
  NAND2X0 U342 ( .IN1(n94), .IN2(n108), .QN(n313) );
  NAND2X0 U343 ( .IN1(n108), .IN2(n123), .QN(n340) );
  NAND2X0 U344 ( .IN1(n343), .IN2(n344), .QN(n298) );
  INVX0 U345 ( .INP(A[3]), .ZN(n375) );
  NAND2X0 U346 ( .IN1(A[3]), .IN2(n370), .QN(n149) );
  NAND2X0 U347 ( .IN1(A[0]), .IN2(n368), .QN(n246) );
  NAND2X1 U348 ( .IN1(B[15]), .IN2(n321), .QN(n288) );
  INVX0 U349 ( .INP(B[15]), .ZN(n320) );
  NAND2X0 U350 ( .IN1(B[7]), .IN2(n381), .QN(n127) );
  INVX0 U351 ( .INP(B[14]), .ZN(n327) );
  NOR2X0 U352 ( .IN1(n250), .IN2(n240), .QN(n249) );
  NAND2X1 U353 ( .IN1(n251), .IN2(n252), .QN(n240) );
  INVX0 U354 ( .INP(n228), .ZN(n231) );
  INVX0 U355 ( .INP(A[0]), .ZN(n391) );
  NAND2X0 U356 ( .IN1(n232), .IN2(n233), .QN(n228) );
  NOR2X0 U357 ( .IN1(n239), .IN2(n79), .QN(n232) );
  NAND2X0 U358 ( .IN1(n305), .IN2(n127), .QN(n360) );
  NAND2X0 U359 ( .IN1(n304), .IN2(n305), .QN(n301) );
  NAND2X1 U360 ( .IN1(n369), .IN2(B[1]), .QN(n171) );
  NAND2X0 U361 ( .IN1(n115), .IN2(n108), .QN(n309) );
  NOR2X0 U362 ( .IN1(n281), .IN2(n282), .QN(n280) );
  INVX0 U363 ( .INP(A[10]), .ZN(n347) );
  NOR2X0 U364 ( .IN1(n294), .IN2(n295), .QN(n281) );
  INVX0 U365 ( .INP(n198), .ZN(n200) );
  NAND2X0 U366 ( .IN1(B[6]), .IN2(n92), .QN(n132) );
  INVX0 U367 ( .INP(B[6]), .ZN(n385) );
  INVX0 U368 ( .INP(A[11]), .ZN(n353) );
  NOR2X0 U369 ( .IN1(n300), .IN2(n299), .QN(n279) );
  NOR2X0 U370 ( .IN1(n309), .IN2(n308), .QN(n299) );
  INVX0 U371 ( .INP(B[5]), .ZN(n384) );
  NAND2X0 U372 ( .IN1(B[10]), .IN2(n347), .QN(n345) );
  NAND2X0 U373 ( .IN1(B[12]), .IN2(n315), .QN(n336) );
  NAND2X0 U374 ( .IN1(n129), .IN2(n132), .QN(n134) );
  NAND2X0 U375 ( .IN1(n131), .IN2(n132), .QN(n130) );
  NAND2X0 U376 ( .IN1(n172), .IN2(n173), .QN(n164) );
  NAND2X0 U377 ( .IN1(n174), .IN2(n66), .QN(n173) );
  NAND2X0 U378 ( .IN1(n127), .IN2(n132), .QN(n379) );
  NAND2X0 U379 ( .IN1(A[8]), .IN2(n346), .QN(n125) );
  NAND2X0 U380 ( .IN1(n218), .IN2(n219), .QN(n212) );
  NAND2X0 U381 ( .IN1(n212), .IN2(n213), .QN(n211) );
  NAND2X0 U382 ( .IN1(n345), .IN2(n349), .QN(n356) );
  NAND2X0 U383 ( .IN1(n355), .IN2(n345), .QN(n354) );
  NAND2X0 U384 ( .IN1(n114), .IN2(n296), .QN(n339) );
  NAND2X0 U385 ( .IN1(n221), .IN2(n220), .QN(n219) );
  NAND2X0 U386 ( .IN1(n297), .IN2(n298), .QN(n294) );
  NAND2X0 U387 ( .IN1(n296), .IN2(n345), .QN(n342) );
  NAND2X0 U388 ( .IN1(n226), .IN2(n227), .QN(n220) );
  NAND2X0 U389 ( .IN1(n228), .IN2(n229), .QN(n227) );
  NAND2X0 U390 ( .IN1(n185), .IN2(n186), .QN(n184) );
  NAND2X0 U391 ( .IN1(n161), .IN2(n162), .QN(n158) );
  NAND2X0 U392 ( .IN1(n190), .IN2(n191), .QN(n185) );
  NAND2X0 U393 ( .IN1(n198), .IN2(n199), .QN(n197) );
  NAND2X0 U394 ( .IN1(n234), .IN2(n235), .QN(n233) );
  XOR2X1 U395 ( .IN1(n116), .IN2(n117), .Q(DIFF[9]) );
  XOR2X1 U396 ( .IN1(n121), .IN2(n122), .Q(DIFF[8]) );
  XOR2X1 U397 ( .IN1(n126), .IN2(n83), .Q(DIFF[7]) );
  XOR2X1 U398 ( .IN1(n133), .IN2(n134), .Q(DIFF[6]) );
  XOR2X1 U399 ( .IN1(n139), .IN2(n140), .Q(DIFF[5]) );
  XOR2X1 U400 ( .IN1(n145), .IN2(n146), .Q(DIFF[4]) );
  XOR2X1 U401 ( .IN1(n148), .IN2(n84), .Q(DIFF[3]) );
  XOR3X1 U402 ( .IN1(n154), .IN2(B[31]), .IN3(n155), .Q(DIFF[31]) );
  XOR2X1 U403 ( .IN1(n152), .IN2(n167), .Q(DIFF[2]) );
  XOR2X1 U404 ( .IN1(n80), .IN2(n180), .Q(DIFF[27]) );
  XOR2X1 U405 ( .IN1(n3), .IN2(n187), .Q(DIFF[26]) );
  XOR2X1 U406 ( .IN1(n2), .IN2(n193), .Q(DIFF[25]) );
  XOR2X1 U407 ( .IN1(n200), .IN2(n201), .Q(DIFF[24]) );
  XOR2X1 U408 ( .IN1(n1), .IN2(n207), .Q(DIFF[23]) );
  XOR2X1 U409 ( .IN1(n214), .IN2(n215), .Q(DIFF[22]) );
  XOR2X1 U410 ( .IN1(n222), .IN2(n223), .Q(DIFF[21]) );
  XOR2X1 U411 ( .IN1(n230), .IN2(n231), .Q(DIFF[20]) );
  XOR2X1 U412 ( .IN1(n244), .IN2(n245), .Q(DIFF[1]) );
  XOR2X1 U413 ( .IN1(n248), .IN2(n249), .Q(DIFF[19]) );
  XOR2X1 U414 ( .IN1(n259), .IN2(n260), .Q(DIFF[18]) );
  XOR2X1 U415 ( .IN1(n269), .IN2(n270), .Q(DIFF[17]) );
  XOR2X1 U416 ( .IN1(n276), .IN2(n91), .Q(DIFF[16]) );
  NAND4X0 U417 ( .IN1(n279), .IN2(n277), .IN3(n280), .IN4(n278), .QN(n235) );
  NAND3X0 U418 ( .IN1(n94), .IN2(n297), .IN3(n310), .QN(n308) );
  XOR2X1 U419 ( .IN1(n319), .IN2(n85), .Q(DIFF[15]) );
  XOR2X1 U420 ( .IN1(n324), .IN2(n325), .Q(DIFF[14]) );
  XOR2X1 U421 ( .IN1(n330), .IN2(n331), .Q(DIFF[13]) );
  XOR2X1 U422 ( .IN1(n337), .IN2(n338), .Q(DIFF[12]) );
  NAND4X0 U423 ( .IN1(A[8]), .IN2(n345), .IN3(n119), .IN4(n346), .QN(n344) );
  XOR2X1 U424 ( .IN1(n351), .IN2(n82), .Q(DIFF[11]) );
  XOR2X1 U425 ( .IN1(n356), .IN2(n357), .Q(DIFF[10]) );
endmodule


module BoothMultiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342;

  OR2X1 U2 ( .IN1(n30), .IN2(n223), .Q(n29) );
  AND2X1 U3 ( .IN1(n65), .IN2(n338), .Q(n119) );
  XOR3X1 U4 ( .IN1(B[28]), .IN2(A[28]), .IN3(n188), .Q(SUM[28]) );
  DELLN1X2 U5 ( .INP(n266), .Z(n114) );
  NAND2X1 U6 ( .IN1(n247), .IN2(n248), .QN(n1) );
  AND2X1 U7 ( .IN1(n274), .IN2(n275), .Q(n2) );
  AND2X1 U8 ( .IN1(n104), .IN2(n232), .Q(n3) );
  AND2X1 U9 ( .IN1(n229), .IN2(n228), .Q(SUM[0]) );
  AND2X1 U10 ( .IN1(n3), .IN2(n225), .Q(n5) );
  AND2X1 U11 ( .IN1(n214), .IN2(n215), .Q(n6) );
  AND2X1 U12 ( .IN1(n210), .IN2(n211), .Q(n7) );
  AND2X1 U13 ( .IN1(n219), .IN2(n220), .Q(n8) );
  AND2X1 U14 ( .IN1(n223), .IN2(n224), .Q(n9) );
  OR2X1 U15 ( .IN1(n105), .IN2(n106), .Q(n10) );
  NAND2X1 U16 ( .IN1(n57), .IN2(n177), .QN(n11) );
  OR2X1 U17 ( .IN1(n122), .IN2(n126), .Q(n12) );
  AND2X1 U18 ( .IN1(B[10]), .IN2(n54), .Q(n109) );
  AND2X1 U19 ( .IN1(n87), .IN2(n88), .Q(n19) );
  AND2X1 U20 ( .IN1(n193), .IN2(n194), .Q(n13) );
  AND2X1 U21 ( .IN1(n197), .IN2(n198), .Q(n14) );
  NAND2X1 U22 ( .IN1(n211), .IN2(n18), .QN(n15) );
  NAND2X1 U23 ( .IN1(n15), .IN2(n16), .QN(n22) );
  OR2X1 U24 ( .IN1(n17), .IN2(n208), .Q(n16) );
  INVX0 U25 ( .INP(n207), .ZN(n17) );
  AND2X1 U26 ( .IN1(n210), .IN2(n207), .Q(n18) );
  AND2X1 U27 ( .IN1(n19), .IN2(n20), .Q(n204) );
  AND2X1 U28 ( .IN1(n97), .IN2(n91), .Q(n20) );
  AND2X1 U29 ( .IN1(n96), .IN2(n97), .Q(n21) );
  AND2X1 U30 ( .IN1(n87), .IN2(n23), .Q(n36) );
  AND2X1 U31 ( .IN1(n91), .IN2(n88), .Q(n23) );
  NAND2X0 U32 ( .IN1(n204), .IN2(n27), .QN(n24) );
  NAND2X0 U33 ( .IN1(n24), .IN2(n25), .QN(n175) );
  OR2X1 U34 ( .IN1(n26), .IN2(n41), .Q(n25) );
  INVX0 U35 ( .INP(n39), .ZN(n26) );
  AND2X1 U36 ( .IN1(n64), .IN2(n39), .Q(n27) );
  NAND2X0 U37 ( .IN1(n1), .IN2(n31), .QN(n28) );
  AND2X1 U38 ( .IN1(n28), .IN2(n29), .Q(n220) );
  INVX0 U39 ( .INP(n221), .ZN(n30) );
  AND2X1 U40 ( .IN1(n5), .IN2(n221), .Q(n31) );
  NAND2X0 U41 ( .IN1(n216), .IN2(n35), .QN(n32) );
  AND2X1 U42 ( .IN1(n32), .IN2(n33), .Q(n211) );
  OR2X1 U43 ( .IN1(n34), .IN2(n214), .Q(n33) );
  INVX0 U44 ( .INP(n212), .ZN(n34) );
  AND2X1 U45 ( .IN1(n217), .IN2(n212), .Q(n35) );
  NAND2X0 U46 ( .IN1(n36), .IN2(n37), .QN(n199) );
  AND2X1 U47 ( .IN1(n203), .IN2(n97), .Q(n37) );
  XNOR3X1 U48 ( .IN1(B[29]), .IN2(A[29]), .IN3(n38), .Q(SUM[29]) );
  NAND2X0 U49 ( .IN1(n50), .IN2(n51), .QN(n38) );
  OR2X1 U50 ( .IN1(n40), .IN2(n60), .Q(n39) );
  INVX0 U51 ( .INP(n58), .ZN(n40) );
  AND2X1 U52 ( .IN1(n62), .IN2(n58), .Q(n41) );
  NAND2X0 U53 ( .IN1(n66), .IN2(n67), .QN(n42) );
  OR2X1 U54 ( .IN1(n42), .IN2(n43), .Q(n47) );
  OR2X1 U55 ( .IN1(n11), .IN2(n45), .Q(n43) );
  NOR2X0 U56 ( .IN1(n44), .IN2(n45), .QN(n190) );
  NAND2X0 U57 ( .IN1(n66), .IN2(n67), .QN(n44) );
  NOR2X0 U58 ( .IN1(n100), .IN2(n193), .QN(n45) );
  NAND3X1 U59 ( .IN1(n172), .IN2(n333), .IN3(n334), .QN(n326) );
  XNOR3X1 U60 ( .IN1(B[30]), .IN2(A[30]), .IN3(n46), .Q(SUM[30]) );
  NAND2X0 U61 ( .IN1(n47), .IN2(n48), .QN(n46) );
  OR2X1 U62 ( .IN1(n49), .IN2(n55), .Q(n48) );
  INVX0 U63 ( .INP(n177), .ZN(n49) );
  NAND2X0 U64 ( .IN1(n190), .IN2(n53), .QN(n50) );
  OR2X1 U65 ( .IN1(n52), .IN2(n187), .Q(n51) );
  INVX0 U66 ( .INP(n186), .ZN(n52) );
  AND2X1 U67 ( .IN1(n189), .IN2(n186), .Q(n53) );
  NBUFFX2 U68 ( .INP(A[10]), .Z(n54) );
  OR2X1 U69 ( .IN1(n56), .IN2(n83), .Q(n55) );
  INVX0 U70 ( .INP(n81), .ZN(n56) );
  AND2X1 U71 ( .IN1(n189), .IN2(n81), .Q(n57) );
  OR2X1 U72 ( .IN1(n59), .IN2(n113), .Q(n58) );
  INVX0 U73 ( .INP(n70), .ZN(n59) );
  AND2X1 U74 ( .IN1(n193), .IN2(n70), .Q(n60) );
  NAND2X0 U75 ( .IN1(n21), .IN2(n64), .QN(n61) );
  NAND2X0 U76 ( .IN1(n61), .IN2(n62), .QN(n194) );
  OR2X1 U77 ( .IN1(n63), .IN2(n86), .Q(n62) );
  INVX0 U78 ( .INP(n84), .ZN(n63) );
  AND2X1 U79 ( .IN1(n203), .IN2(n84), .Q(n64) );
  NOR2X0 U80 ( .IN1(n75), .IN2(n142), .QN(n65) );
  NAND2X0 U81 ( .IN1(n199), .IN2(n69), .QN(n66) );
  OR2X1 U82 ( .IN1(n68), .IN2(n197), .Q(n67) );
  INVX0 U83 ( .INP(n101), .ZN(n68) );
  AND2X1 U84 ( .IN1(n200), .IN2(n101), .Q(n69) );
  AND2X1 U85 ( .IN1(n111), .IN2(n12), .Q(n70) );
  NAND2X1 U86 ( .IN1(n297), .IN2(n298), .QN(n292) );
  NAND2X0 U87 ( .IN1(n226), .IN2(n74), .QN(n71) );
  AND2X1 U88 ( .IN1(n71), .IN2(n72), .Q(n77) );
  OR2X1 U89 ( .IN1(n73), .IN2(n223), .Q(n72) );
  INVX0 U90 ( .INP(n80), .ZN(n73) );
  AND2X1 U91 ( .IN1(n5), .IN2(n80), .Q(n74) );
  AND2X1 U92 ( .IN1(n302), .IN2(n301), .Q(n300) );
  INVX0 U93 ( .INP(n148), .ZN(n75) );
  NAND2X0 U94 ( .IN1(n1), .IN2(n5), .QN(n224) );
  AND2X1 U95 ( .IN1(n333), .IN2(n172), .Q(n328) );
  NAND2X0 U96 ( .IN1(n203), .IN2(n21), .QN(n76) );
  AND2X1 U97 ( .IN1(n77), .IN2(n78), .Q(n87) );
  OR2X1 U98 ( .IN1(n79), .IN2(n219), .Q(n78) );
  INVX0 U99 ( .INP(n90), .ZN(n79) );
  AND2X1 U100 ( .IN1(n221), .IN2(n90), .Q(n80) );
  OR2X1 U101 ( .IN1(n82), .IN2(n186), .Q(n81) );
  INVX0 U102 ( .INP(n178), .ZN(n82) );
  AND2X1 U103 ( .IN1(n187), .IN2(n178), .Q(n83) );
  OR2X1 U104 ( .IN1(n85), .IN2(n197), .Q(n84) );
  INVX0 U105 ( .INP(n195), .ZN(n85) );
  AND2X1 U106 ( .IN1(n200), .IN2(n195), .Q(n86) );
  OR2X1 U107 ( .IN1(n89), .IN2(n214), .Q(n88) );
  INVX0 U108 ( .INP(n93), .ZN(n89) );
  AND2X1 U109 ( .IN1(n217), .IN2(n93), .Q(n90) );
  NAND2X0 U110 ( .IN1(n94), .IN2(n95), .QN(n230) );
  NAND2X0 U111 ( .IN1(n3), .IN2(n1), .QN(n95) );
  AND2X1 U112 ( .IN1(n19), .IN2(n91), .Q(n96) );
  OR2X1 U113 ( .IN1(n92), .IN2(n210), .Q(n91) );
  INVX0 U114 ( .INP(n99), .ZN(n92) );
  AND2X1 U115 ( .IN1(n212), .IN2(n99), .Q(n93) );
  NAND2X0 U116 ( .IN1(n153), .IN2(n154), .QN(n152) );
  NAND3X1 U117 ( .IN1(n310), .IN2(n301), .IN3(n311), .QN(n305) );
  NAND2X0 U118 ( .IN1(n317), .IN2(n318), .QN(n314) );
  NAND2X0 U119 ( .IN1(n323), .IN2(n324), .QN(n135) );
  NAND2X0 U120 ( .IN1(n158), .IN2(n159), .QN(n153) );
  NAND2X0 U121 ( .IN1(n239), .IN2(n240), .QN(n235) );
  NAND2X0 U122 ( .IN1(n139), .IN2(n322), .QN(n130) );
  AND2X1 U123 ( .IN1(n233), .IN2(n234), .Q(n94) );
  NAND2X0 U124 ( .IN1(n219), .IN2(n221), .QN(n222) );
  NAND2X0 U125 ( .IN1(B[21]), .IN2(A[21]), .QN(n214) );
  NAND2X0 U126 ( .IN1(B[22]), .IN2(A[22]), .QN(n210) );
  OR2X1 U127 ( .IN1(n98), .IN2(n207), .Q(n97) );
  INVX0 U128 ( .INP(n205), .ZN(n98) );
  AND2X1 U129 ( .IN1(n208), .IN2(n205), .Q(n99) );
  NAND2X0 U130 ( .IN1(n247), .IN2(n248), .QN(n226) );
  INVX0 U131 ( .INP(n191), .ZN(n100) );
  AND2X1 U132 ( .IN1(n195), .IN2(n191), .Q(n101) );
  INVX0 U133 ( .INP(n302), .ZN(n138) );
  INVX0 U134 ( .INP(n282), .ZN(n283) );
  NAND2X0 U135 ( .IN1(n151), .IN2(n152), .QN(n147) );
  OR2X1 U136 ( .IN1(n235), .IN2(n102), .Q(n236) );
  AND2X1 U137 ( .IN1(n104), .IN2(n1), .Q(n102) );
  NOR2X0 U138 ( .IN1(n156), .IN2(n157), .QN(n155) );
  INVX0 U139 ( .INP(n151), .ZN(n156) );
  NOR2X0 U140 ( .IN1(n264), .IN2(n118), .QN(n294) );
  NOR2X0 U141 ( .IN1(n180), .IN2(n181), .QN(n179) );
  OR2X1 U142 ( .IN1(B[5]), .IN2(A[5]), .Q(n154) );
  NOR2X0 U143 ( .IN1(n110), .IN2(n10), .QN(n223) );
  AND2X1 U144 ( .IN1(n256), .IN2(n257), .Q(n103) );
  INVX0 U145 ( .INP(n242), .ZN(n241) );
  NOR2X0 U146 ( .IN1(n277), .IN2(n118), .QN(n274) );
  INVX0 U147 ( .INP(n169), .ZN(n180) );
  NAND2X0 U148 ( .IN1(n302), .IN2(n135), .QN(n322) );
  NAND2X0 U149 ( .IN1(n290), .IN2(n291), .QN(n286) );
  NAND2X0 U150 ( .IN1(n292), .IN2(n293), .QN(n290) );
  NAND2X0 U151 ( .IN1(n258), .IN2(n285), .QN(n282) );
  INVX0 U152 ( .INP(n172), .ZN(n181) );
  NAND2X0 U153 ( .IN1(n271), .IN2(n281), .QN(n278) );
  AND2X1 U154 ( .IN1(n232), .IN2(n225), .Q(n117) );
  INVX0 U155 ( .INP(n182), .ZN(n334) );
  AND2X1 U156 ( .IN1(n237), .IN2(n238), .Q(n104) );
  INVX0 U157 ( .INP(n301), .ZN(n133) );
  NAND2X0 U158 ( .IN1(n134), .IN2(n321), .QN(n319) );
  NAND2X0 U159 ( .IN1(n301), .IN2(n130), .QN(n321) );
  NAND2X0 U160 ( .IN1(n119), .IN2(n114), .QN(n324) );
  NAND2X0 U161 ( .IN1(n250), .IN2(n251), .QN(n249) );
  INVX0 U162 ( .INP(n272), .ZN(n303) );
  INVX0 U163 ( .INP(n253), .ZN(n142) );
  NAND2X0 U164 ( .IN1(n269), .IN2(n270), .QN(n268) );
  INVX0 U165 ( .INP(n271), .ZN(n269) );
  AND2X1 U166 ( .IN1(n235), .IN2(n117), .Q(n105) );
  NOR2X0 U167 ( .IN1(n116), .IN2(n234), .QN(n106) );
  NAND2X0 U168 ( .IN1(n145), .IN2(n146), .QN(n140) );
  NAND2X0 U169 ( .IN1(n160), .IN2(n114), .QN(n159) );
  INVX0 U170 ( .INP(n291), .ZN(n264) );
  NAND2X0 U171 ( .IN1(n244), .IN2(n242), .QN(n243) );
  NAND2X0 U172 ( .IN1(n235), .IN2(n232), .QN(n233) );
  INVX0 U173 ( .INP(n146), .ZN(n150) );
  INVX0 U174 ( .INP(n250), .ZN(n280) );
  INVX0 U175 ( .INP(n228), .ZN(n184) );
  NAND2X0 U176 ( .IN1(n185), .IN2(n182), .QN(n227) );
  NAND2X0 U177 ( .IN1(n182), .IN2(n183), .QN(n171) );
  NAND2X1 U178 ( .IN1(n184), .IN2(n185), .QN(n183) );
  NOR2X0 U179 ( .IN1(n303), .IN2(n316), .QN(n315) );
  INVX0 U180 ( .INP(n306), .ZN(n316) );
  NOR2X0 U181 ( .IN1(n142), .IN2(n143), .QN(n141) );
  INVX0 U182 ( .INP(n144), .ZN(n143) );
  NOR2X0 U183 ( .IN1(n132), .IN2(n133), .QN(n131) );
  INVX0 U184 ( .INP(n134), .ZN(n132) );
  NOR2X0 U185 ( .IN1(n289), .IN2(n277), .QN(n288) );
  INVX0 U186 ( .INP(n258), .ZN(n289) );
  NOR2X0 U187 ( .IN1(n162), .IN2(n163), .QN(n161) );
  INVX0 U188 ( .INP(n158), .ZN(n162) );
  NOR2X0 U189 ( .IN1(n137), .IN2(n138), .QN(n136) );
  INVX0 U190 ( .INP(n139), .ZN(n137) );
  NAND2X0 U191 ( .IN1(n237), .IN2(n242), .QN(n246) );
  NAND2X0 U192 ( .IN1(n169), .IN2(n170), .QN(n164) );
  NOR2X0 U193 ( .IN1(n166), .IN2(n167), .QN(n165) );
  INVX0 U194 ( .INP(n168), .ZN(n166) );
  AND2X1 U195 ( .IN1(n234), .IN2(n232), .Q(n107) );
  AND2X1 U196 ( .IN1(n240), .IN2(n238), .Q(n108) );
  NOR2X0 U197 ( .IN1(n110), .IN2(n116), .QN(n231) );
  NAND2X1 U198 ( .IN1(n189), .IN2(n191), .QN(n192) );
  NAND2X1 U199 ( .IN1(n214), .IN2(n217), .QN(n218) );
  NAND2X1 U200 ( .IN1(n210), .IN2(n212), .QN(n213) );
  NAND2X1 U201 ( .IN1(n207), .IN2(n208), .QN(n209) );
  NAND2X1 U202 ( .IN1(n203), .IN2(n205), .QN(n206) );
  NAND2X1 U203 ( .IN1(n197), .IN2(n200), .QN(n202) );
  NAND2X1 U204 ( .IN1(n193), .IN2(n195), .QN(n196) );
  NAND2X0 U205 ( .IN1(n144), .IN2(n146), .QN(n341) );
  OR2X1 U206 ( .IN1(B[13]), .IN2(A[13]), .Q(n287) );
  OR2X1 U207 ( .IN1(B[18]), .IN2(A[18]), .Q(n232) );
  OR2X1 U208 ( .IN1(B[11]), .IN2(A[11]), .Q(n272) );
  OR2X1 U209 ( .IN1(B[7]), .IN2(A[7]), .Q(n253) );
  OR2X1 U210 ( .IN1(B[14]), .IN2(A[14]), .Q(n257) );
  OR2X1 U211 ( .IN1(B[6]), .IN2(A[6]), .Q(n148) );
  OR2X1 U212 ( .IN1(B[10]), .IN2(A[10]), .Q(n310) );
  OR2X1 U213 ( .IN1(B[3]), .IN2(A[3]), .Q(n333) );
  OR2X1 U214 ( .IN1(B[9]), .IN2(A[9]), .Q(n301) );
  OR2X1 U215 ( .IN1(B[19]), .IN2(A[19]), .Q(n225) );
  NOR2X0 U216 ( .IN1(n115), .IN2(n330), .QN(n329) );
  OR2X1 U217 ( .IN1(B[4]), .IN2(A[4]), .Q(n160) );
  OR2X1 U218 ( .IN1(B[16]), .IN2(A[16]), .Q(n237) );
  INVX0 U219 ( .INP(A[8]), .ZN(n312) );
  OR2X1 U220 ( .IN1(B[17]), .IN2(A[17]), .Q(n238) );
  OR2X1 U221 ( .IN1(B[15]), .IN2(A[15]), .Q(n270) );
  NAND2X0 U222 ( .IN1(B[18]), .IN2(A[18]), .QN(n234) );
  AND2X1 U223 ( .IN1(B[19]), .IN2(A[19]), .Q(n110) );
  NAND2X0 U224 ( .IN1(B[20]), .IN2(A[20]), .QN(n219) );
  NAND2X1 U225 ( .IN1(B[23]), .IN2(A[23]), .QN(n207) );
  NAND2X1 U226 ( .IN1(B[24]), .IN2(A[24]), .QN(n203) );
  NAND2X1 U227 ( .IN1(B[25]), .IN2(A[25]), .QN(n197) );
  OR2X1 U228 ( .IN1(B[29]), .IN2(A[29]), .Q(n178) );
  OR2X1 U229 ( .IN1(B[28]), .IN2(A[28]), .Q(n187) );
  OR2X1 U230 ( .IN1(B[30]), .IN2(A[30]), .Q(n176) );
  NAND2X1 U231 ( .IN1(B[29]), .IN2(A[29]), .QN(n177) );
  OR2X1 U232 ( .IN1(B[20]), .IN2(A[20]), .Q(n221) );
  OR2X1 U233 ( .IN1(B[21]), .IN2(A[21]), .Q(n217) );
  OR2X1 U234 ( .IN1(B[24]), .IN2(A[24]), .Q(n205) );
  OR2X1 U235 ( .IN1(B[25]), .IN2(A[25]), .Q(n200) );
  OR2X1 U236 ( .IN1(B[26]), .IN2(A[26]), .Q(n195) );
  OR2X1 U237 ( .IN1(B[22]), .IN2(A[22]), .Q(n212) );
  OR2X1 U238 ( .IN1(B[23]), .IN2(A[23]), .Q(n208) );
  NAND2X1 U239 ( .IN1(B[27]), .IN2(A[27]), .QN(n189) );
  OR2X1 U240 ( .IN1(B[0]), .IN2(A[0]), .Q(n229) );
  NAND2X1 U241 ( .IN1(B[26]), .IN2(A[26]), .QN(n193) );
  OR2X1 U242 ( .IN1(B[27]), .IN2(A[27]), .Q(n191) );
  NAND2X1 U243 ( .IN1(B[28]), .IN2(A[28]), .QN(n186) );
  NAND2X1 U244 ( .IN1(B[30]), .IN2(A[30]), .QN(n174) );
  INVX0 U245 ( .INP(n1), .ZN(n245) );
  INVX0 U246 ( .INP(n76), .ZN(n201) );
  OR2X1 U247 ( .IN1(n112), .IN2(n189), .Q(n111) );
  INVX0 U248 ( .INP(n123), .ZN(n112) );
  AND2X1 U249 ( .IN1(n191), .IN2(n123), .Q(n113) );
  INVX0 U250 ( .INP(n333), .ZN(n167) );
  NAND2X0 U251 ( .IN1(n180), .IN2(n333), .QN(n325) );
  NOR2X0 U252 ( .IN1(n150), .IN2(n75), .QN(n149) );
  NAND2X0 U253 ( .IN1(n286), .IN2(n287), .QN(n285) );
  INVX0 U254 ( .INP(n287), .ZN(n277) );
  AND2X1 U255 ( .IN1(n331), .IN2(n332), .Q(n115) );
  INVX0 U256 ( .INP(n225), .ZN(n116) );
  AND2X1 U257 ( .IN1(n295), .IN2(n296), .Q(n118) );
  NAND4X0 U258 ( .IN1(B[4]), .IN2(A[4]), .IN3(n154), .IN4(n148), .QN(n340) );
  INVX0 U259 ( .INP(n154), .ZN(n157) );
  NOR2X0 U260 ( .IN1(n75), .IN2(n142), .QN(n337) );
  NAND2X0 U261 ( .IN1(n337), .IN2(n338), .QN(n254) );
  AND2X1 U262 ( .IN1(n299), .IN2(n300), .Q(n120) );
  NOR2X0 U263 ( .IN1(n303), .IN2(n304), .QN(n299) );
  INVX0 U264 ( .INP(n270), .ZN(n121) );
  NAND2X1 U265 ( .IN1(n295), .IN2(n296), .QN(n293) );
  NOR2X0 U266 ( .IN1(n109), .IN2(n309), .QN(n320) );
  NAND2X0 U267 ( .IN1(n319), .IN2(n310), .QN(n318) );
  NAND2X0 U268 ( .IN1(n273), .IN2(n272), .QN(n297) );
  NOR2X0 U269 ( .IN1(n309), .IN2(n134), .QN(n308) );
  INVX0 U270 ( .INP(A[2]), .ZN(n336) );
  NAND2X1 U271 ( .IN1(n335), .IN2(n336), .QN(n172) );
  NAND2X0 U272 ( .IN1(n299), .IN2(n300), .QN(n255) );
  NAND2X0 U273 ( .IN1(n147), .IN2(n148), .QN(n145) );
  NAND2X0 U274 ( .IN1(n339), .IN2(n340), .QN(n252) );
  INVX0 U275 ( .INP(B[2]), .ZN(n335) );
  INVX0 U276 ( .INP(A[12]), .ZN(n296) );
  NOR2X0 U277 ( .IN1(n280), .IN2(n259), .QN(n279) );
  NOR2X0 U278 ( .IN1(n121), .IN2(n276), .QN(n275) );
  NOR2X0 U279 ( .IN1(n258), .IN2(n259), .QN(n256) );
  INVX0 U280 ( .INP(n270), .ZN(n259) );
  INVX0 U281 ( .INP(n124), .ZN(n122) );
  AND2X1 U282 ( .IN1(n187), .IN2(n124), .Q(n123) );
  INVX0 U283 ( .INP(B[12]), .ZN(n295) );
  NAND2X1 U284 ( .IN1(n313), .IN2(n312), .QN(n302) );
  NOR2X0 U285 ( .IN1(n312), .IN2(n313), .QN(n311) );
  INVX0 U286 ( .INP(B[8]), .ZN(n313) );
  NAND2X0 U287 ( .IN1(n257), .IN2(n271), .QN(n284) );
  NAND2X0 U288 ( .IN1(n282), .IN2(n257), .QN(n281) );
  INVX0 U289 ( .INP(n257), .ZN(n276) );
  INVX0 U290 ( .INP(A[1]), .ZN(n332) );
  NAND2X0 U291 ( .IN1(B[13]), .IN2(A[13]), .QN(n258) );
  NAND2X0 U292 ( .IN1(B[4]), .IN2(A[4]), .QN(n158) );
  OR2X1 U293 ( .IN1(n125), .IN2(n129), .Q(n124) );
  INVX0 U294 ( .INP(n127), .ZN(n125) );
  AND2X1 U295 ( .IN1(n186), .IN2(n127), .Q(n126) );
  NAND2X0 U296 ( .IN1(B[9]), .IN2(A[9]), .QN(n134) );
  NAND2X0 U297 ( .IN1(n241), .IN2(n238), .QN(n239) );
  NAND2X0 U298 ( .IN1(B[17]), .IN2(A[17]), .QN(n240) );
  NAND2X0 U299 ( .IN1(B[3]), .IN2(A[3]), .QN(n168) );
  OR2X1 U300 ( .IN1(n128), .IN2(n177), .Q(n127) );
  INVX0 U301 ( .INP(n176), .ZN(n128) );
  AND2X1 U302 ( .IN1(n178), .IN2(n176), .Q(n129) );
  NAND2X0 U303 ( .IN1(B[0]), .IN2(A[0]), .QN(n228) );
  NAND2X1 U304 ( .IN1(B[16]), .IN2(A[16]), .QN(n242) );
  NAND2X0 U305 ( .IN1(B[15]), .IN2(A[15]), .QN(n250) );
  NAND2X0 U306 ( .IN1(n252), .IN2(n253), .QN(n323) );
  NAND2X0 U307 ( .IN1(B[7]), .IN2(A[7]), .QN(n144) );
  NAND2X0 U308 ( .IN1(B[14]), .IN2(A[14]), .QN(n271) );
  NAND2X0 U309 ( .IN1(n120), .IN2(n135), .QN(n298) );
  NAND2X0 U310 ( .IN1(n264), .IN2(n2), .QN(n263) );
  NAND2X0 U311 ( .IN1(B[0]), .IN2(A[0]), .QN(n330) );
  NAND2X0 U312 ( .IN1(n171), .IN2(n172), .QN(n170) );
  NAND2X0 U313 ( .IN1(n328), .IN2(n329), .QN(n327) );
  NAND2X0 U314 ( .IN1(B[2]), .IN2(A[2]), .QN(n169) );
  INVX0 U315 ( .INP(n310), .ZN(n309) );
  NOR2X0 U316 ( .IN1(n308), .IN2(n109), .QN(n307) );
  NOR2X0 U317 ( .IN1(n342), .IN2(n341), .QN(n339) );
  NOR2X0 U318 ( .IN1(n254), .IN2(n255), .QN(n265) );
  INVX0 U319 ( .INP(B[1]), .ZN(n331) );
  NAND2X1 U320 ( .IN1(n331), .IN2(n332), .QN(n185) );
  NAND2X0 U321 ( .IN1(B[1]), .IN2(A[1]), .QN(n182) );
  NAND2X0 U322 ( .IN1(n262), .IN2(n263), .QN(n261) );
  NOR2X0 U323 ( .IN1(n163), .IN2(n157), .QN(n338) );
  INVX0 U324 ( .INP(n160), .ZN(n163) );
  NOR2X0 U325 ( .IN1(n75), .IN2(n151), .QN(n342) );
  NOR2X0 U326 ( .IN1(n260), .IN2(n261), .QN(n247) );
  NAND2X0 U327 ( .IN1(n174), .IN2(n175), .QN(n173) );
  NAND2X0 U328 ( .IN1(B[5]), .IN2(A[5]), .QN(n151) );
  NAND2X0 U329 ( .IN1(n267), .IN2(n268), .QN(n260) );
  NAND2X0 U330 ( .IN1(n237), .IN2(n1), .QN(n244) );
  NAND2X0 U331 ( .IN1(B[12]), .IN2(A[12]), .QN(n291) );
  NAND2X0 U332 ( .IN1(n189), .IN2(n190), .QN(n188) );
  NAND2X0 U333 ( .IN1(B[11]), .IN2(A[11]), .QN(n306) );
  NAND2X0 U334 ( .IN1(B[8]), .IN2(A[8]), .QN(n139) );
  NAND2X0 U335 ( .IN1(n216), .IN2(n217), .QN(n215) );
  NOR2X0 U336 ( .IN1(n103), .IN2(n249), .QN(n248) );
  NAND2X0 U337 ( .IN1(n219), .IN2(n220), .QN(n216) );
  NAND2X0 U338 ( .IN1(n200), .IN2(n76), .QN(n198) );
  NAND2X0 U339 ( .IN1(B[6]), .IN2(A[6]), .QN(n146) );
  NAND2X0 U340 ( .IN1(B[10]), .IN2(n54), .QN(n317) );
  NOR2X0 U341 ( .IN1(n54), .IN2(B[10]), .QN(n304) );
  XOR2X1 U342 ( .IN1(n130), .IN2(n131), .Q(SUM[9]) );
  XOR2X1 U343 ( .IN1(n135), .IN2(n136), .Q(SUM[8]) );
  XOR2X1 U344 ( .IN1(n140), .IN2(n141), .Q(SUM[7]) );
  XOR2X1 U345 ( .IN1(n147), .IN2(n149), .Q(SUM[6]) );
  XOR2X1 U346 ( .IN1(n153), .IN2(n155), .Q(SUM[5]) );
  XOR2X1 U347 ( .IN1(n114), .IN2(n161), .Q(SUM[4]) );
  XOR2X1 U348 ( .IN1(n164), .IN2(n165), .Q(SUM[3]) );
  XOR3X1 U349 ( .IN1(B[31]), .IN2(A[31]), .IN3(n173), .Q(SUM[31]) );
  XOR2X1 U350 ( .IN1(n171), .IN2(n179), .Q(SUM[2]) );
  XOR2X1 U351 ( .IN1(n13), .IN2(n192), .Q(SUM[27]) );
  XOR2X1 U352 ( .IN1(n14), .IN2(n196), .Q(SUM[26]) );
  XOR2X1 U353 ( .IN1(n201), .IN2(n202), .Q(SUM[25]) );
  XOR2X1 U354 ( .IN1(n22), .IN2(n206), .Q(SUM[24]) );
  XOR2X1 U355 ( .IN1(n7), .IN2(n209), .Q(SUM[23]) );
  XOR2X1 U356 ( .IN1(n6), .IN2(n213), .Q(SUM[22]) );
  XOR2X1 U357 ( .IN1(n8), .IN2(n218), .Q(SUM[21]) );
  XOR2X1 U358 ( .IN1(n9), .IN2(n222), .Q(SUM[20]) );
  XOR2X1 U359 ( .IN1(n227), .IN2(n228), .Q(SUM[1]) );
  XOR2X1 U360 ( .IN1(n230), .IN2(n231), .Q(SUM[19]) );
  XOR2X1 U361 ( .IN1(n236), .IN2(n107), .Q(SUM[18]) );
  XOR2X1 U362 ( .IN1(n243), .IN2(n108), .Q(SUM[17]) );
  XOR2X1 U363 ( .IN1(n245), .IN2(n246), .Q(SUM[16]) );
  NAND4X0 U364 ( .IN1(n252), .IN2(n2), .IN3(n120), .IN4(n253), .QN(n251) );
  NAND3X0 U365 ( .IN1(n265), .IN2(n2), .IN3(n266), .QN(n262) );
  NAND3X0 U366 ( .IN1(n2), .IN2(n272), .IN3(n273), .QN(n267) );
  XOR2X1 U367 ( .IN1(n278), .IN2(n279), .Q(SUM[15]) );
  XOR2X1 U368 ( .IN1(n283), .IN2(n284), .Q(SUM[14]) );
  XOR2X1 U369 ( .IN1(n286), .IN2(n288), .Q(SUM[13]) );
  XOR2X1 U370 ( .IN1(n292), .IN2(n294), .Q(SUM[12]) );
  NAND3X0 U371 ( .IN1(n307), .IN2(n306), .IN3(n305), .QN(n273) );
  XOR2X1 U372 ( .IN1(n314), .IN2(n315), .Q(SUM[11]) );
  XOR2X1 U373 ( .IN1(n319), .IN2(n320), .Q(SUM[10]) );
  NAND4X0 U374 ( .IN1(n325), .IN2(n326), .IN3(n327), .IN4(n168), .QN(n266) );
endmodule


module BoothMultiplier ( clk, oClk, rst, oRst, M, Q, P );
  input [31:0] M;
  input [31:0] Q;
  output [63:0] P;
  input clk, oClk, rst, oRst;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N110, N111, N112, N113, N114, n8, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411;
  wire   [31:0] Acc;
  wire   [5:0] count;
  wire   [31:0] M_reg;
  wire   [64:33] case_add;
  wire   [64:33] case_sub;

  DFFX1 \P_reg[6]  ( .D(N12), .CLK(oClk), .Q(P[6]) );
  DFFX1 \P_reg[5]  ( .D(N11), .CLK(oClk), .Q(P[5]) );
  DFFX1 \P_reg[4]  ( .D(N10), .CLK(oClk), .Q(P[4]) );
  DFFX1 \P_reg[32]  ( .D(N38), .CLK(oClk), .Q(P[32]) );
  DFFX1 \P_reg[33]  ( .D(N39), .CLK(oClk), .Q(P[33]) );
  DFFX1 \P_reg[34]  ( .D(N40), .CLK(oClk), .Q(P[34]) );
  DFFX1 \P_reg[35]  ( .D(N41), .CLK(oClk), .Q(P[35]) );
  DFFX1 \P_reg[36]  ( .D(N42), .CLK(oClk), .Q(P[36]) );
  DFFX1 \P_reg[37]  ( .D(N43), .CLK(oClk), .Q(P[37]) );
  DFFX1 \P_reg[38]  ( .D(N44), .CLK(oClk), .Q(P[38]) );
  DFFX1 \P_reg[39]  ( .D(N45), .CLK(oClk), .Q(P[39]) );
  DFFX1 \P_reg[40]  ( .D(N46), .CLK(oClk), .Q(P[40]) );
  DFFX1 \P_reg[41]  ( .D(N47), .CLK(oClk), .Q(P[41]) );
  DFFX1 \P_reg[42]  ( .D(N48), .CLK(oClk), .Q(P[42]) );
  DFFX1 \P_reg[43]  ( .D(N49), .CLK(oClk), .Q(P[43]) );
  DFFX1 \P_reg[44]  ( .D(N50), .CLK(oClk), .Q(P[44]) );
  DFFX1 \P_reg[45]  ( .D(N51), .CLK(oClk), .Q(P[45]) );
  DFFX1 \P_reg[46]  ( .D(N52), .CLK(oClk), .Q(P[46]) );
  DFFX1 \P_reg[47]  ( .D(N53), .CLK(oClk), .Q(P[47]) );
  DFFX1 \P_reg[48]  ( .D(N54), .CLK(oClk), .Q(P[48]) );
  DFFX1 \P_reg[49]  ( .D(N55), .CLK(oClk), .Q(P[49]) );
  DFFX1 \P_reg[50]  ( .D(N56), .CLK(oClk), .Q(P[50]) );
  DFFX1 \P_reg[51]  ( .D(N57), .CLK(oClk), .Q(P[51]) );
  DFFX1 \P_reg[52]  ( .D(N58), .CLK(oClk), .Q(P[52]) );
  DFFX1 \P_reg[53]  ( .D(N59), .CLK(oClk), .Q(P[53]) );
  DFFX1 \P_reg[54]  ( .D(N60), .CLK(oClk), .Q(P[54]) );
  DFFX1 \P_reg[55]  ( .D(N61), .CLK(oClk), .Q(P[55]) );
  DFFX1 \P_reg[56]  ( .D(N62), .CLK(oClk), .Q(P[56]) );
  DFFX1 \P_reg[57]  ( .D(N63), .CLK(oClk), .Q(P[57]) );
  DFFX1 \P_reg[58]  ( .D(N64), .CLK(oClk), .Q(P[58]) );
  DFFX1 \P_reg[59]  ( .D(N65), .CLK(oClk), .Q(P[59]) );
  DFFX1 \P_reg[60]  ( .D(N66), .CLK(oClk), .Q(P[60]) );
  DFFX1 \P_reg[61]  ( .D(N67), .CLK(oClk), .Q(P[61]) );
  DFFX1 \P_reg[63]  ( .D(n325), .CLK(oClk), .Q(P[63]) );
  DFFX1 \P_reg[62]  ( .D(n325), .CLK(oClk), .Q(P[62]) );
  DFFX1 \P_reg[0]  ( .D(N6), .CLK(oClk), .Q(P[0]) );
  DFFX1 \P_reg[1]  ( .D(N7), .CLK(oClk), .Q(P[1]) );
  DFFX1 \P_reg[2]  ( .D(N8), .CLK(oClk), .Q(P[2]) );
  DFFX1 \P_reg[3]  ( .D(N9), .CLK(oClk), .Q(P[3]) );
  DFFX1 \P_reg[7]  ( .D(N13), .CLK(oClk), .Q(P[7]) );
  DFFX1 \P_reg[8]  ( .D(N14), .CLK(oClk), .Q(P[8]) );
  DFFX1 \P_reg[9]  ( .D(N15), .CLK(oClk), .Q(P[9]) );
  DFFX1 \P_reg[10]  ( .D(N16), .CLK(oClk), .Q(P[10]) );
  DFFX1 \P_reg[11]  ( .D(N17), .CLK(oClk), .Q(P[11]) );
  DFFX1 \P_reg[12]  ( .D(N18), .CLK(oClk), .Q(P[12]) );
  DFFX1 \P_reg[13]  ( .D(N19), .CLK(oClk), .Q(P[13]) );
  DFFX1 \P_reg[14]  ( .D(N20), .CLK(oClk), .Q(P[14]) );
  DFFX1 \P_reg[15]  ( .D(N21), .CLK(oClk), .Q(P[15]) );
  DFFX1 \P_reg[16]  ( .D(N22), .CLK(oClk), .Q(P[16]) );
  DFFX1 \P_reg[17]  ( .D(N23), .CLK(oClk), .Q(P[17]) );
  DFFX1 \P_reg[18]  ( .D(N24), .CLK(oClk), .Q(P[18]) );
  DFFX1 \P_reg[19]  ( .D(N25), .CLK(oClk), .Q(P[19]) );
  DFFX1 \P_reg[20]  ( .D(N26), .CLK(oClk), .Q(P[20]) );
  DFFX1 \P_reg[21]  ( .D(N27), .CLK(oClk), .Q(P[21]) );
  DFFX1 \P_reg[22]  ( .D(N28), .CLK(oClk), .Q(P[22]) );
  DFFX1 \P_reg[23]  ( .D(N29), .CLK(oClk), .Q(P[23]) );
  DFFX1 \P_reg[24]  ( .D(N30), .CLK(oClk), .Q(P[24]) );
  DFFX1 \P_reg[25]  ( .D(N31), .CLK(oClk), .Q(P[25]) );
  DFFX1 \P_reg[26]  ( .D(N32), .CLK(oClk), .Q(P[26]) );
  DFFX1 \P_reg[27]  ( .D(N33), .CLK(oClk), .Q(P[27]) );
  DFFX1 \P_reg[28]  ( .D(N34), .CLK(oClk), .Q(P[28]) );
  DFFX1 \P_reg[29]  ( .D(N35), .CLK(oClk), .Q(P[29]) );
  DFFX1 \P_reg[30]  ( .D(N36), .CLK(oClk), .Q(P[30]) );
  DFFX1 \P_reg[31]  ( .D(N37), .CLK(oClk), .Q(P[31]) );
  DFFX1 \M_reg_reg[31]  ( .D(n280), .CLK(clk), .Q(M_reg[31]) );
  DFFX1 \M_reg_reg[30]  ( .D(n279), .CLK(clk), .Q(M_reg[30]) );
  DFFX1 \M_reg_reg[29]  ( .D(n278), .CLK(clk), .Q(M_reg[29]) );
  DFFX1 \M_reg_reg[28]  ( .D(n277), .CLK(clk), .Q(M_reg[28]) );
  DFFX1 \M_reg_reg[27]  ( .D(n276), .CLK(clk), .Q(M_reg[27]) );
  DFFX1 \M_reg_reg[26]  ( .D(n275), .CLK(clk), .Q(M_reg[26]) );
  DFFX1 \M_reg_reg[25]  ( .D(n274), .CLK(clk), .Q(M_reg[25]) );
  DFFX1 \M_reg_reg[24]  ( .D(n273), .CLK(clk), .Q(M_reg[24]) );
  DFFX1 \M_reg_reg[23]  ( .D(n272), .CLK(clk), .Q(M_reg[23]) );
  DFFX1 \M_reg_reg[22]  ( .D(n271), .CLK(clk), .Q(M_reg[22]) );
  DFFX1 \M_reg_reg[21]  ( .D(n270), .CLK(clk), .Q(M_reg[21]) );
  DFFX1 \M_reg_reg[20]  ( .D(n269), .CLK(clk), .Q(M_reg[20]) );
  DFFX1 \M_reg_reg[19]  ( .D(n268), .CLK(clk), .Q(M_reg[19]) );
  DFFX1 \M_reg_reg[18]  ( .D(n267), .CLK(clk), .Q(M_reg[18]) );
  DFFX1 \M_reg_reg[17]  ( .D(n266), .CLK(clk), .Q(M_reg[17]) );
  DFFX1 \M_reg_reg[16]  ( .D(n265), .CLK(clk), .Q(M_reg[16]) );
  DFFX1 \M_reg_reg[15]  ( .D(n264), .CLK(clk), .Q(M_reg[15]) );
  DFFX1 \M_reg_reg[14]  ( .D(n263), .CLK(clk), .Q(M_reg[14]) );
  DFFX1 \M_reg_reg[13]  ( .D(n262), .CLK(clk), .Q(M_reg[13]) );
  DFFX1 \M_reg_reg[12]  ( .D(n261), .CLK(clk), .Q(M_reg[12]) );
  DFFX1 \M_reg_reg[11]  ( .D(n260), .CLK(clk), .Q(M_reg[11]) );
  DFFX1 \M_reg_reg[10]  ( .D(n259), .CLK(clk), .Q(M_reg[10]), .QN(n338) );
  DFFX1 \M_reg_reg[9]  ( .D(n258), .CLK(clk), .Q(M_reg[9]), .QN(n333) );
  DFFX1 \M_reg_reg[8]  ( .D(n257), .CLK(clk), .Q(M_reg[8]) );
  DFFX1 \M_reg_reg[7]  ( .D(n256), .CLK(clk), .Q(M_reg[7]) );
  DFFX1 \M_reg_reg[6]  ( .D(n255), .CLK(clk), .Q(M_reg[6]), .QN(n331) );
  DFFX1 \M_reg_reg[5]  ( .D(n254), .CLK(clk), .Q(M_reg[5]), .QN(n336) );
  DFFX1 \M_reg_reg[4]  ( .D(n253), .CLK(clk), .Q(M_reg[4]) );
  DFFX1 \M_reg_reg[3]  ( .D(n252), .CLK(clk), .Q(M_reg[3]) );
  DFFX1 \M_reg_reg[2]  ( .D(n251), .CLK(clk), .Q(M_reg[2]) );
  DFFX1 \M_reg_reg[1]  ( .D(n250), .CLK(clk), .Q(M_reg[1]) );
  DFFX1 \M_reg_reg[0]  ( .D(n249), .CLK(clk), .Q(M_reg[0]) );
  DFFX1 \count_reg[0]  ( .D(n248), .CLK(clk), .Q(count[0]), .QN(n316) );
  DFFX1 \count_reg[5]  ( .D(n247), .CLK(clk), .Q(count[5]) );
  DFFX1 \count_reg[4]  ( .D(n246), .CLK(clk), .Q(count[4]) );
  DFFX1 \count_reg[3]  ( .D(n245), .CLK(clk), .Q(count[3]) );
  DFFX1 \count_reg[2]  ( .D(n244), .CLK(clk), .Q(count[2]), .QN(n298) );
  DFFX1 \count_reg[1]  ( .D(n243), .CLK(clk), .Q(count[1]) );
  DFFX1 \Acc_reg[0]  ( .D(n242), .CLK(clk), .Q(Acc[0]), .QN(n177) );
  DFFX1 \Q_reg_reg[31]  ( .D(n241), .CLK(clk), .Q(n315), .QN(n173) );
  DFFX1 \Q_reg_reg[30]  ( .D(n240), .CLK(clk), .Q(n293), .QN(n172) );
  DFFX1 \Q_reg_reg[29]  ( .D(n239), .CLK(clk), .Q(n309), .QN(n171) );
  DFFX1 \Q_reg_reg[28]  ( .D(n238), .CLK(clk), .Q(n292), .QN(n170) );
  DFFX1 \Q_reg_reg[27]  ( .D(n237), .CLK(clk), .Q(n308), .QN(n169) );
  DFFX1 \Q_reg_reg[26]  ( .D(n236), .CLK(clk), .Q(n291), .QN(n168) );
  DFFX1 \Q_reg_reg[25]  ( .D(n235), .CLK(clk), .Q(n307), .QN(n167) );
  DFFX1 \Q_reg_reg[24]  ( .D(n234), .CLK(clk), .Q(n290), .QN(n166) );
  DFFX1 \Q_reg_reg[23]  ( .D(n233), .CLK(clk), .Q(n306), .QN(n165) );
  DFFX1 \Q_reg_reg[22]  ( .D(n232), .CLK(clk), .Q(n289), .QN(n164) );
  DFFX1 \Q_reg_reg[21]  ( .D(n231), .CLK(clk), .Q(n305), .QN(n163) );
  DFFX1 \Q_reg_reg[20]  ( .D(n230), .CLK(clk), .Q(n288), .QN(n162) );
  DFFX1 \Q_reg_reg[19]  ( .D(n229), .CLK(clk), .Q(n304), .QN(n161) );
  DFFX1 \Q_reg_reg[18]  ( .D(n228), .CLK(clk), .Q(n287), .QN(n160) );
  DFFX1 \Q_reg_reg[17]  ( .D(n227), .CLK(clk), .Q(n303), .QN(n159) );
  DFFX1 \Q_reg_reg[16]  ( .D(n226), .CLK(clk), .Q(n286), .QN(n158) );
  DFFX1 \Q_reg_reg[15]  ( .D(n225), .CLK(clk), .Q(n302), .QN(n157) );
  DFFX1 \Q_reg_reg[14]  ( .D(n224), .CLK(clk), .Q(n285), .QN(n156) );
  DFFX1 \Q_reg_reg[13]  ( .D(n223), .CLK(clk), .Q(n301), .QN(n155) );
  DFFX1 \Q_reg_reg[12]  ( .D(n222), .CLK(clk), .Q(n284), .QN(n154) );
  DFFX1 \Q_reg_reg[11]  ( .D(n221), .CLK(clk), .Q(n282), .QN(n153) );
  DFFX1 \Q_reg_reg[10]  ( .D(n220), .CLK(clk), .Q(n314), .QN(n152) );
  DFFX1 \Q_reg_reg[9]  ( .D(n219), .CLK(clk), .Q(n297), .QN(n151) );
  DFFX1 \Q_reg_reg[8]  ( .D(n218), .CLK(clk), .Q(n313), .QN(n150) );
  DFFX1 \Q_reg_reg[7]  ( .D(n217), .CLK(clk), .Q(n296), .QN(n149) );
  DFFX1 \Q_reg_reg[6]  ( .D(n216), .CLK(clk), .Q(n312), .QN(n148) );
  DFFX1 \Q_reg_reg[5]  ( .D(n215), .CLK(clk), .Q(n295), .QN(n147) );
  DFFX1 \Q_reg_reg[4]  ( .D(n214), .CLK(clk), .Q(n311), .QN(n146) );
  DFFX1 \Q_reg_reg[3]  ( .D(n213), .CLK(clk), .Q(n294), .QN(n145) );
  DFFX1 \Q_reg_reg[2]  ( .D(n212), .CLK(clk), .Q(n310), .QN(n144) );
  DFFX1 \Q_reg_reg[1]  ( .D(n211), .CLK(clk), .Q(n283), .QN(n143) );
  DFFX1 \Q_reg_reg[0]  ( .D(n210), .CLK(clk), .Q(n281), .QN(n175) );
  DFFX1 Q_prev_reg ( .D(n209), .CLK(clk), .Q(n174), .QN(n300) );
  DFFX1 \Acc_reg[31]  ( .D(n208), .CLK(clk), .Q(n299) );
  DFFX1 \Acc_reg[30]  ( .D(n207), .CLK(clk), .Q(Acc[30]), .QN(n141) );
  DFFX1 \Acc_reg[29]  ( .D(n206), .CLK(clk), .Q(Acc[29]), .QN(n140) );
  DFFX1 \Acc_reg[28]  ( .D(n205), .CLK(clk), .Q(Acc[28]), .QN(n139) );
  DFFX1 \Acc_reg[27]  ( .D(n204), .CLK(clk), .Q(Acc[27]), .QN(n138) );
  DFFX1 \Acc_reg[26]  ( .D(n203), .CLK(clk), .Q(Acc[26]), .QN(n137) );
  DFFX1 \Acc_reg[25]  ( .D(n202), .CLK(clk), .Q(Acc[25]), .QN(n136) );
  DFFX1 \Acc_reg[24]  ( .D(n201), .CLK(clk), .Q(Acc[24]), .QN(n135) );
  DFFX1 \Acc_reg[23]  ( .D(n200), .CLK(clk), .Q(Acc[23]), .QN(n134) );
  DFFX1 \Acc_reg[22]  ( .D(n199), .CLK(clk), .Q(Acc[22]), .QN(n133) );
  DFFX1 \Acc_reg[21]  ( .D(n198), .CLK(clk), .Q(Acc[21]), .QN(n132) );
  DFFX1 \Acc_reg[20]  ( .D(n197), .CLK(clk), .Q(Acc[20]), .QN(n131) );
  DFFX1 \Acc_reg[19]  ( .D(n196), .CLK(clk), .Q(Acc[19]), .QN(n130) );
  DFFX1 \Acc_reg[18]  ( .D(n195), .CLK(clk), .Q(Acc[18]), .QN(n129) );
  DFFX1 \Acc_reg[17]  ( .D(n194), .CLK(clk), .Q(Acc[17]), .QN(n128) );
  DFFX1 \Acc_reg[16]  ( .D(n193), .CLK(clk), .Q(Acc[16]), .QN(n127) );
  DFFX1 \Acc_reg[15]  ( .D(n192), .CLK(clk), .Q(Acc[15]), .QN(n126) );
  DFFX1 \Acc_reg[14]  ( .D(n191), .CLK(clk), .Q(Acc[14]), .QN(n125) );
  DFFX1 \Acc_reg[13]  ( .D(n190), .CLK(clk), .Q(Acc[13]), .QN(n124) );
  DFFX1 \Acc_reg[12]  ( .D(n189), .CLK(clk), .Q(Acc[12]), .QN(n123) );
  DFFX1 \Acc_reg[11]  ( .D(n188), .CLK(clk), .Q(Acc[11]), .QN(n122) );
  DFFX1 \Acc_reg[10]  ( .D(n187), .CLK(clk), .Q(Acc[10]), .QN(n121) );
  DFFX1 \Acc_reg[9]  ( .D(n186), .CLK(clk), .Q(Acc[9]), .QN(n120) );
  DFFX1 \Acc_reg[8]  ( .D(n185), .CLK(clk), .Q(Acc[8]), .QN(n119) );
  DFFX1 \Acc_reg[7]  ( .D(n184), .CLK(clk), .Q(Acc[7]), .QN(n118) );
  DFFX1 \Acc_reg[6]  ( .D(n183), .CLK(clk), .Q(Acc[6]), .QN(n117) );
  DFFX1 \Acc_reg[5]  ( .D(n182), .CLK(clk), .Q(Acc[5]), .QN(n116) );
  DFFX1 \Acc_reg[4]  ( .D(n181), .CLK(clk), .Q(Acc[4]), .QN(n115) );
  DFFX1 \Acc_reg[3]  ( .D(n180), .CLK(clk), .Q(Acc[3]), .QN(n114) );
  DFFX1 \Acc_reg[2]  ( .D(n179), .CLK(clk), .Q(Acc[2]), .QN(n113) );
  DFFX1 \Acc_reg[1]  ( .D(n178), .CLK(clk), .Q(Acc[1]), .QN(n176) );
  AO22X1 U3 ( .IN1(n352), .IN2(count[5]), .IN3(N114), .IN4(n355), .Q(n247) );
  AO221X1 U4 ( .IN1(N113), .IN2(n411), .IN3(n352), .IN4(count[4]), .IN5(n362), 
        .Q(n246) );
  AO221X1 U5 ( .IN1(N112), .IN2(n411), .IN3(n352), .IN4(count[3]), .IN5(n362), 
        .Q(n245) );
  AO221X1 U6 ( .IN1(N111), .IN2(n411), .IN3(n352), .IN4(count[2]), .IN5(n362), 
        .Q(n244) );
  AO221X1 U10 ( .IN1(N110), .IN2(n411), .IN3(n352), .IN4(count[1]), .IN5(n362), 
        .Q(n243) );
  AO221X1 U11 ( .IN1(n316), .IN2(n411), .IN3(n352), .IN4(count[0]), .IN5(n362), 
        .Q(n248) );
  AO222X1 U12 ( .IN1(n355), .IN2(n314), .IN3(Q[9]), .IN4(n362), .IN5(n352), 
        .IN6(n297), .Q(n219) );
  AO222X1 U13 ( .IN1(n355), .IN2(n297), .IN3(Q[8]), .IN4(n362), .IN5(n351), 
        .IN6(n313), .Q(n218) );
  AO222X1 U15 ( .IN1(n355), .IN2(n313), .IN3(Q[7]), .IN4(n363), .IN5(n351), 
        .IN6(n296), .Q(n217) );
  AO222X1 U17 ( .IN1(n355), .IN2(n296), .IN3(Q[6]), .IN4(n363), .IN5(n351), 
        .IN6(n312), .Q(n216) );
  AO222X1 U19 ( .IN1(n355), .IN2(n312), .IN3(Q[5]), .IN4(n363), .IN5(n351), 
        .IN6(n295), .Q(n215) );
  AO222X1 U21 ( .IN1(n355), .IN2(n295), .IN3(Q[4]), .IN4(n363), .IN5(n351), 
        .IN6(n311), .Q(n214) );
  AO222X1 U23 ( .IN1(n355), .IN2(n311), .IN3(Q[3]), .IN4(n363), .IN5(n351), 
        .IN6(n294), .Q(n213) );
  AO222X1 U27 ( .IN1(n355), .IN2(n315), .IN3(Q[30]), .IN4(n363), .IN5(n351), 
        .IN6(n293), .Q(n240) );
  AO222X1 U29 ( .IN1(n355), .IN2(n294), .IN3(Q[2]), .IN4(n363), .IN5(n351), 
        .IN6(n310), .Q(n212) );
  AO222X1 U31 ( .IN1(n355), .IN2(n293), .IN3(Q[29]), .IN4(n363), .IN5(n351), 
        .IN6(n309), .Q(n239) );
  AO222X1 U33 ( .IN1(n355), .IN2(n309), .IN3(Q[28]), .IN4(n363), .IN5(n352), 
        .IN6(n292), .Q(n238) );
  AO222X1 U35 ( .IN1(n355), .IN2(n292), .IN3(Q[27]), .IN4(n363), .IN5(n351), 
        .IN6(n308), .Q(n237) );
  AO222X1 U37 ( .IN1(n356), .IN2(n308), .IN3(Q[26]), .IN4(n363), .IN5(n351), 
        .IN6(n291), .Q(n236) );
  AO222X1 U39 ( .IN1(n356), .IN2(n291), .IN3(Q[25]), .IN4(n363), .IN5(n351), 
        .IN6(n307), .Q(n235) );
  AO222X1 U41 ( .IN1(n356), .IN2(n307), .IN3(Q[24]), .IN4(n363), .IN5(n351), 
        .IN6(n290), .Q(n234) );
  AO222X1 U43 ( .IN1(n356), .IN2(n290), .IN3(Q[23]), .IN4(n363), .IN5(n351), 
        .IN6(n306), .Q(n233) );
  AO222X1 U45 ( .IN1(n356), .IN2(n306), .IN3(Q[22]), .IN4(n363), .IN5(n351), 
        .IN6(n289), .Q(n232) );
  AO222X1 U47 ( .IN1(n356), .IN2(n289), .IN3(Q[21]), .IN4(n363), .IN5(n350), 
        .IN6(n305), .Q(n231) );
  AO222X1 U49 ( .IN1(n356), .IN2(n305), .IN3(Q[20]), .IN4(n363), .IN5(n350), 
        .IN6(n288), .Q(n230) );
  AO222X1 U51 ( .IN1(n356), .IN2(n310), .IN3(Q[1]), .IN4(n363), .IN5(n350), 
        .IN6(n283), .Q(n211) );
  AO222X1 U53 ( .IN1(n356), .IN2(n288), .IN3(Q[19]), .IN4(n363), .IN5(n350), 
        .IN6(n304), .Q(n229) );
  AO222X1 U55 ( .IN1(n356), .IN2(n304), .IN3(Q[18]), .IN4(n363), .IN5(n350), 
        .IN6(n287), .Q(n228) );
  AO222X1 U57 ( .IN1(n356), .IN2(n287), .IN3(Q[17]), .IN4(n363), .IN5(n350), 
        .IN6(n303), .Q(n227) );
  AO222X1 U59 ( .IN1(n356), .IN2(n303), .IN3(Q[16]), .IN4(n363), .IN5(n350), 
        .IN6(n286), .Q(n226) );
  AO222X1 U61 ( .IN1(n356), .IN2(n286), .IN3(Q[15]), .IN4(n363), .IN5(n350), 
        .IN6(n302), .Q(n225) );
  AO222X1 U63 ( .IN1(n357), .IN2(n302), .IN3(Q[14]), .IN4(n363), .IN5(n351), 
        .IN6(n285), .Q(n224) );
  AO222X1 U65 ( .IN1(n357), .IN2(n285), .IN3(Q[13]), .IN4(n363), .IN5(n350), 
        .IN6(n301), .Q(n223) );
  AO222X1 U67 ( .IN1(n357), .IN2(n301), .IN3(Q[12]), .IN4(n363), .IN5(n350), 
        .IN6(n284), .Q(n222) );
  AO222X1 U69 ( .IN1(n357), .IN2(n284), .IN3(Q[11]), .IN4(n363), .IN5(n350), 
        .IN6(n282), .Q(n221) );
  AO222X1 U71 ( .IN1(n357), .IN2(n282), .IN3(Q[10]), .IN4(n362), .IN5(n350), 
        .IN6(n314), .Q(n220) );
  BoothMultiplier_DW01_sub_1 sub_61 ( .A({n299, Acc[30:0]}), .B({M_reg[31:11], 
        n339, n334, M_reg[8:7], n332, M_reg[5:0]}), .CI(1'b0), .DIFF(case_sub)
         );
  BoothMultiplier_DW01_add_1 add_57 ( .A({n299, Acc[30:11], n340, Acc[9:7], 
        n335, n330, Acc[4:2], n398, n320}), .B({M_reg[31:6], n337, M_reg[4:0]}), .CI(1'b0), .SUM(case_add) );
  NBUFFX2 U278 ( .INP(n117), .Z(n321) );
  MUX21X1 U279 ( .IN1(M_reg[2]), .IN2(M[2]), .S(n363), .Q(n251) );
  AND2X1 U280 ( .IN1(n317), .IN2(n318), .Q(n319) );
  NAND2X0 U281 ( .IN1(case_sub[62]), .IN2(n347), .QN(n317) );
  AOI22X1 U282 ( .IN1(n354), .IN2(Acc[28]), .IN3(n341), .IN4(Acc[29]), .QN(
        n318) );
  INVX0 U283 ( .INP(n177), .ZN(n320) );
  MUX21X1 U284 ( .IN1(M_reg[10]), .IN2(M[10]), .S(n363), .Q(n259) );
  NAND2X0 U285 ( .IN1(n322), .IN2(n319), .QN(n205) );
  NAND2X0 U286 ( .IN1(n344), .IN2(case_add[62]), .QN(n322) );
  INVX0 U287 ( .INP(Acc[10]), .ZN(n323) );
  NBUFFX2 U288 ( .INP(n8), .Z(n357) );
  NBUFFX2 U289 ( .INP(n402), .Z(n354) );
  NOR2X0 U290 ( .IN1(n350), .IN2(n363), .QN(n8) );
  INVX0 U291 ( .INP(n411), .ZN(n402) );
  NBUFFX2 U292 ( .INP(n328), .Z(n349) );
  NBUFFX2 U293 ( .INP(n326), .Z(n343) );
  NBUFFX2 U294 ( .INP(n327), .Z(n346) );
  AND2X1 U295 ( .IN1(n411), .IN2(n364), .Q(n324) );
  INVX0 U296 ( .INP(n364), .ZN(n362) );
  INVX0 U297 ( .INP(n364), .ZN(n363) );
  INVX0 U298 ( .INP(n405), .ZN(n409) );
  INVX0 U299 ( .INP(n403), .ZN(n407) );
  INVX0 U300 ( .INP(n404), .ZN(n408) );
  AND2X1 U301 ( .IN1(n299), .IN2(n361), .Q(n325) );
  INVX0 U302 ( .INP(n361), .ZN(n360) );
  INVX0 U303 ( .INP(n361), .ZN(n359) );
  INVX0 U304 ( .INP(n361), .ZN(n358) );
  AND3X1 U305 ( .IN1(n366), .IN2(n364), .IN3(n365), .Q(n326) );
  AND3X1 U306 ( .IN1(n174), .IN2(n175), .IN3(n324), .Q(n327) );
  AND3X1 U307 ( .IN1(n281), .IN2(n300), .IN3(n324), .Q(n328) );
  INVX0 U308 ( .INP(rst), .ZN(n364) );
  NOR2X0 U309 ( .IN1(count[1]), .IN2(n410), .QN(n329) );
  MUX21X1 U310 ( .IN1(M_reg[3]), .IN2(M[3]), .S(rst), .Q(n252) );
  MUX21X1 U311 ( .IN1(M_reg[4]), .IN2(M[4]), .S(rst), .Q(n253) );
  MUX21X1 U312 ( .IN1(M_reg[6]), .IN2(M[6]), .S(rst), .Q(n255) );
  MUX21X1 U313 ( .IN1(M_reg[7]), .IN2(M[7]), .S(rst), .Q(n256) );
  MUX21X1 U314 ( .IN1(M_reg[9]), .IN2(M[9]), .S(rst), .Q(n258) );
  MUX21X1 U315 ( .IN1(M_reg[11]), .IN2(M[11]), .S(rst), .Q(n260) );
  MUX21X1 U316 ( .IN1(M_reg[12]), .IN2(M[12]), .S(rst), .Q(n261) );
  MUX21X1 U317 ( .IN1(M_reg[13]), .IN2(M[13]), .S(rst), .Q(n262) );
  MUX21X1 U318 ( .IN1(M_reg[14]), .IN2(M[14]), .S(rst), .Q(n263) );
  MUX21X1 U319 ( .IN1(M_reg[15]), .IN2(M[15]), .S(rst), .Q(n264) );
  MUX21X1 U320 ( .IN1(M_reg[16]), .IN2(M[16]), .S(rst), .Q(n265) );
  MUX21X1 U321 ( .IN1(M_reg[17]), .IN2(M[17]), .S(rst), .Q(n266) );
  NOR2X0 U322 ( .IN1(n360), .IN2(n129), .QN(N55) );
  NOR2X0 U323 ( .IN1(n360), .IN2(n128), .QN(N54) );
  NOR2X0 U324 ( .IN1(n360), .IN2(n127), .QN(N53) );
  NOR2X0 U325 ( .IN1(n360), .IN2(n126), .QN(N52) );
  NOR2X0 U326 ( .IN1(n360), .IN2(n125), .QN(N51) );
  NOR2X0 U327 ( .IN1(n360), .IN2(n124), .QN(N50) );
  NOR2X0 U328 ( .IN1(n360), .IN2(n123), .QN(N49) );
  NOR2X0 U329 ( .IN1(n360), .IN2(n122), .QN(N48) );
  NOR2X0 U330 ( .IN1(n360), .IN2(n323), .QN(N47) );
  NOR2X0 U331 ( .IN1(n360), .IN2(n120), .QN(N46) );
  NOR2X0 U332 ( .IN1(n359), .IN2(n177), .QN(N37) );
  NOR2X0 U333 ( .IN1(n358), .IN2(n141), .QN(N67) );
  NOR2X0 U334 ( .IN1(n359), .IN2(n140), .QN(N66) );
  NOR2X0 U335 ( .IN1(n358), .IN2(n139), .QN(N65) );
  NOR2X0 U336 ( .IN1(n359), .IN2(n138), .QN(N64) );
  NOR2X0 U337 ( .IN1(n358), .IN2(n137), .QN(N63) );
  NOR2X0 U338 ( .IN1(n359), .IN2(n136), .QN(N62) );
  NOR2X0 U339 ( .IN1(n358), .IN2(n135), .QN(N61) );
  NOR2X0 U340 ( .IN1(oRst), .IN2(n134), .QN(N60) );
  NOR2X0 U341 ( .IN1(oRst), .IN2(n133), .QN(N59) );
  NOR2X0 U342 ( .IN1(oRst), .IN2(n132), .QN(N58) );
  NOR2X0 U343 ( .IN1(oRst), .IN2(n131), .QN(N57) );
  NOR2X0 U344 ( .IN1(oRst), .IN2(n130), .QN(N56) );
  NOR2X0 U345 ( .IN1(oRst), .IN2(n119), .QN(N45) );
  NOR2X0 U346 ( .IN1(oRst), .IN2(n118), .QN(N44) );
  NOR2X0 U347 ( .IN1(oRst), .IN2(n321), .QN(N43) );
  NOR2X0 U348 ( .IN1(oRst), .IN2(n116), .QN(N42) );
  NOR2X0 U349 ( .IN1(oRst), .IN2(n115), .QN(N41) );
  NOR2X0 U350 ( .IN1(oRst), .IN2(n114), .QN(N40) );
  NOR2X0 U351 ( .IN1(oRst), .IN2(n113), .QN(N39) );
  NOR2X0 U352 ( .IN1(oRst), .IN2(n176), .QN(N38) );
  NOR2X0 U353 ( .IN1(n360), .IN2(n173), .QN(N36) );
  NOR2X0 U354 ( .IN1(n360), .IN2(n172), .QN(N35) );
  NOR2X0 U355 ( .IN1(n360), .IN2(n171), .QN(N34) );
  NOR2X0 U356 ( .IN1(n360), .IN2(n146), .QN(N9) );
  NOR2X0 U357 ( .IN1(n360), .IN2(n145), .QN(N8) );
  NOR2X0 U358 ( .IN1(n360), .IN2(n144), .QN(N7) );
  NOR2X0 U359 ( .IN1(n360), .IN2(n143), .QN(N6) );
  NOR2X0 U360 ( .IN1(n359), .IN2(n170), .QN(N33) );
  NOR2X0 U361 ( .IN1(n359), .IN2(n169), .QN(N32) );
  NOR2X0 U362 ( .IN1(n359), .IN2(n168), .QN(N31) );
  NOR2X0 U363 ( .IN1(n359), .IN2(n167), .QN(N30) );
  NOR2X0 U364 ( .IN1(n359), .IN2(n166), .QN(N29) );
  NOR2X0 U365 ( .IN1(n359), .IN2(n165), .QN(N28) );
  NOR2X0 U366 ( .IN1(n359), .IN2(n164), .QN(N27) );
  NOR2X0 U367 ( .IN1(n359), .IN2(n163), .QN(N26) );
  NOR2X0 U368 ( .IN1(n359), .IN2(n162), .QN(N25) );
  NOR2X0 U369 ( .IN1(n359), .IN2(n161), .QN(N24) );
  NOR2X0 U370 ( .IN1(n359), .IN2(n160), .QN(N23) );
  NOR2X0 U371 ( .IN1(n359), .IN2(n159), .QN(N22) );
  NOR2X0 U372 ( .IN1(n358), .IN2(n158), .QN(N21) );
  NOR2X0 U373 ( .IN1(n358), .IN2(n157), .QN(N20) );
  NOR2X0 U374 ( .IN1(n358), .IN2(n156), .QN(N19) );
  NOR2X0 U375 ( .IN1(n358), .IN2(n155), .QN(N18) );
  NOR2X0 U376 ( .IN1(n358), .IN2(n154), .QN(N17) );
  NOR2X0 U377 ( .IN1(n358), .IN2(n153), .QN(N16) );
  NOR2X0 U378 ( .IN1(n358), .IN2(n152), .QN(N15) );
  NOR2X0 U379 ( .IN1(n358), .IN2(n151), .QN(N14) );
  NOR2X0 U380 ( .IN1(n358), .IN2(n150), .QN(N13) );
  NOR2X0 U381 ( .IN1(n358), .IN2(n147), .QN(N10) );
  NOR2X0 U382 ( .IN1(n358), .IN2(n148), .QN(N11) );
  NOR2X0 U383 ( .IN1(n358), .IN2(n149), .QN(N12) );
  INVX0 U384 ( .INP(n321), .ZN(n392) );
  INVX0 U385 ( .INP(n141), .ZN(n367) );
  INVX0 U386 ( .INP(n125), .ZN(n383) );
  INVX0 U387 ( .INP(n176), .ZN(n398) );
  INVX0 U388 ( .INP(oRst), .ZN(n361) );
  INVX0 U389 ( .INP(n116), .ZN(n330) );
  INVX0 U390 ( .INP(n331), .ZN(n332) );
  INVX0 U391 ( .INP(n333), .ZN(n334) );
  INVX0 U392 ( .INP(n117), .ZN(n335) );
  INVX0 U393 ( .INP(n336), .ZN(n337) );
  INVX0 U394 ( .INP(n338), .ZN(n339) );
  INVX0 U395 ( .INP(n121), .ZN(n340) );
  NBUFFX2 U396 ( .INP(n326), .Z(n341) );
  NBUFFX2 U397 ( .INP(n326), .Z(n342) );
  NBUFFX2 U398 ( .INP(n327), .Z(n344) );
  NBUFFX2 U399 ( .INP(n327), .Z(n345) );
  NBUFFX2 U400 ( .INP(n328), .Z(n347) );
  NBUFFX2 U401 ( .INP(n328), .Z(n348) );
  NBUFFX2 U402 ( .INP(n402), .Z(n350) );
  NBUFFX2 U403 ( .INP(n402), .Z(n351) );
  NBUFFX2 U404 ( .INP(n402), .Z(n352) );
  NBUFFX2 U405 ( .INP(n402), .Z(n353) );
  NBUFFX2 U406 ( .INP(n8), .Z(n355) );
  NBUFFX2 U407 ( .INP(n8), .Z(n356) );
  NAND4X0 U408 ( .IN1(n329), .IN2(n298), .IN3(n316), .IN4(n364), .QN(n411) );
  AO222X1 U409 ( .IN1(n283), .IN2(n357), .IN3(n350), .IN4(n281), .IN5(Q[0]), 
        .IN6(n363), .Q(n210) );
  AO22X1 U410 ( .IN1(n174), .IN2(n352), .IN3(n357), .IN4(n281), .Q(n209) );
  XOR2X1 U411 ( .IN1(n174), .IN2(n175), .Q(n366) );
  NAND3X0 U412 ( .IN1(n298), .IN2(n316), .IN3(n329), .QN(n365) );
  AO222X1 U413 ( .IN1(case_sub[64]), .IN2(n349), .IN3(n344), .IN4(case_add[64]), .IN5(n341), .IN6(n299), .Q(n400) );
  AO21X1 U414 ( .IN1(n352), .IN2(n367), .IN3(n400), .Q(n207) );
  AO22X1 U415 ( .IN1(n354), .IN2(Acc[29]), .IN3(n341), .IN4(n367), .Q(n368) );
  AO221X1 U416 ( .IN1(n344), .IN2(case_add[63]), .IN3(case_sub[63]), .IN4(n347), .IN5(n368), .Q(n206) );
  AO22X1 U417 ( .IN1(n354), .IN2(Acc[27]), .IN3(n341), .IN4(Acc[28]), .Q(n369)
         );
  AO221X1 U418 ( .IN1(case_add[61]), .IN2(n344), .IN3(case_sub[61]), .IN4(n347), .IN5(n369), .Q(n204) );
  AO22X1 U419 ( .IN1(n354), .IN2(Acc[26]), .IN3(n341), .IN4(Acc[27]), .Q(n370)
         );
  AO221X1 U420 ( .IN1(case_add[60]), .IN2(n344), .IN3(case_sub[60]), .IN4(n347), .IN5(n370), .Q(n203) );
  AO22X1 U421 ( .IN1(n353), .IN2(Acc[25]), .IN3(n341), .IN4(Acc[26]), .Q(n371)
         );
  AO221X1 U422 ( .IN1(case_add[59]), .IN2(n344), .IN3(case_sub[59]), .IN4(n347), .IN5(n371), .Q(n202) );
  AO22X1 U423 ( .IN1(n353), .IN2(Acc[24]), .IN3(n341), .IN4(Acc[25]), .Q(n372)
         );
  AO221X1 U424 ( .IN1(case_add[58]), .IN2(n344), .IN3(case_sub[58]), .IN4(n347), .IN5(n372), .Q(n201) );
  AO22X1 U425 ( .IN1(n353), .IN2(Acc[23]), .IN3(n341), .IN4(Acc[24]), .Q(n373)
         );
  AO221X1 U426 ( .IN1(case_add[57]), .IN2(n344), .IN3(case_sub[57]), .IN4(n347), .IN5(n373), .Q(n200) );
  AO22X1 U427 ( .IN1(n353), .IN2(Acc[22]), .IN3(n342), .IN4(Acc[23]), .Q(n374)
         );
  AO221X1 U428 ( .IN1(case_add[56]), .IN2(n345), .IN3(case_sub[56]), .IN4(n348), .IN5(n374), .Q(n199) );
  AO22X1 U429 ( .IN1(n353), .IN2(Acc[21]), .IN3(n341), .IN4(Acc[22]), .Q(n375)
         );
  AO221X1 U430 ( .IN1(case_add[55]), .IN2(n344), .IN3(case_sub[55]), .IN4(n347), .IN5(n375), .Q(n198) );
  AO22X1 U431 ( .IN1(n353), .IN2(Acc[20]), .IN3(n341), .IN4(Acc[21]), .Q(n376)
         );
  AO221X1 U432 ( .IN1(case_add[54]), .IN2(n344), .IN3(case_sub[54]), .IN4(n347), .IN5(n376), .Q(n197) );
  AO22X1 U433 ( .IN1(n353), .IN2(Acc[19]), .IN3(n341), .IN4(Acc[20]), .Q(n377)
         );
  AO221X1 U434 ( .IN1(case_add[53]), .IN2(n344), .IN3(case_sub[53]), .IN4(n347), .IN5(n377), .Q(n196) );
  AO22X1 U435 ( .IN1(n353), .IN2(Acc[18]), .IN3(n341), .IN4(Acc[19]), .Q(n378)
         );
  AO221X1 U436 ( .IN1(case_add[52]), .IN2(n344), .IN3(case_sub[52]), .IN4(n347), .IN5(n378), .Q(n195) );
  AO22X1 U437 ( .IN1(n354), .IN2(Acc[17]), .IN3(n342), .IN4(Acc[18]), .Q(n379)
         );
  AO221X1 U438 ( .IN1(case_add[51]), .IN2(n345), .IN3(case_sub[51]), .IN4(n347), .IN5(n379), .Q(n194) );
  AO22X1 U439 ( .IN1(n353), .IN2(Acc[16]), .IN3(n342), .IN4(Acc[17]), .Q(n380)
         );
  AO221X1 U440 ( .IN1(case_add[50]), .IN2(n345), .IN3(case_sub[50]), .IN4(n348), .IN5(n380), .Q(n193) );
  AO22X1 U441 ( .IN1(n353), .IN2(Acc[15]), .IN3(n342), .IN4(Acc[16]), .Q(n381)
         );
  AO221X1 U442 ( .IN1(case_add[49]), .IN2(n345), .IN3(case_sub[49]), .IN4(n348), .IN5(n381), .Q(n192) );
  AO22X1 U443 ( .IN1(n353), .IN2(n383), .IN3(n342), .IN4(Acc[15]), .Q(n382) );
  AO221X1 U444 ( .IN1(case_add[48]), .IN2(n345), .IN3(case_sub[48]), .IN4(n348), .IN5(n382), .Q(n191) );
  AO22X1 U445 ( .IN1(n353), .IN2(Acc[13]), .IN3(n342), .IN4(n383), .Q(n384) );
  AO221X1 U446 ( .IN1(case_add[47]), .IN2(n345), .IN3(case_sub[47]), .IN4(n348), .IN5(n384), .Q(n190) );
  AO22X1 U447 ( .IN1(n353), .IN2(Acc[12]), .IN3(n342), .IN4(Acc[13]), .Q(n385)
         );
  AO221X1 U448 ( .IN1(case_add[46]), .IN2(n345), .IN3(case_sub[46]), .IN4(n348), .IN5(n385), .Q(n189) );
  AO22X1 U449 ( .IN1(n353), .IN2(Acc[11]), .IN3(n342), .IN4(Acc[12]), .Q(n386)
         );
  AO221X1 U450 ( .IN1(case_add[45]), .IN2(n345), .IN3(case_sub[45]), .IN4(n348), .IN5(n386), .Q(n188) );
  AO22X1 U451 ( .IN1(n353), .IN2(n340), .IN3(n342), .IN4(Acc[11]), .Q(n387) );
  AO221X1 U452 ( .IN1(case_add[44]), .IN2(n345), .IN3(case_sub[44]), .IN4(n348), .IN5(n387), .Q(n187) );
  AO22X1 U453 ( .IN1(n353), .IN2(Acc[9]), .IN3(n342), .IN4(Acc[10]), .Q(n388)
         );
  AO221X1 U454 ( .IN1(case_add[43]), .IN2(n345), .IN3(case_sub[43]), .IN4(n348), .IN5(n388), .Q(n186) );
  AO22X1 U455 ( .IN1(n353), .IN2(Acc[8]), .IN3(n342), .IN4(Acc[9]), .Q(n389)
         );
  AO221X1 U456 ( .IN1(case_add[42]), .IN2(n345), .IN3(case_sub[42]), .IN4(n348), .IN5(n389), .Q(n185) );
  AO22X1 U457 ( .IN1(n352), .IN2(Acc[7]), .IN3(n342), .IN4(Acc[8]), .Q(n390)
         );
  AO221X1 U458 ( .IN1(case_add[41]), .IN2(n345), .IN3(case_sub[41]), .IN4(n348), .IN5(n390), .Q(n184) );
  AO22X1 U459 ( .IN1(n353), .IN2(n392), .IN3(n342), .IN4(Acc[7]), .Q(n391) );
  AO221X1 U460 ( .IN1(case_add[40]), .IN2(n345), .IN3(case_sub[40]), .IN4(n348), .IN5(n391), .Q(n183) );
  AO22X1 U461 ( .IN1(n352), .IN2(n330), .IN3(n342), .IN4(n392), .Q(n393) );
  AO221X1 U462 ( .IN1(case_add[39]), .IN2(n345), .IN3(case_sub[39]), .IN4(n349), .IN5(n393), .Q(n182) );
  AO22X1 U463 ( .IN1(n352), .IN2(Acc[4]), .IN3(n343), .IN4(Acc[5]), .Q(n394)
         );
  AO221X1 U464 ( .IN1(case_add[38]), .IN2(n346), .IN3(case_sub[38]), .IN4(n349), .IN5(n394), .Q(n181) );
  AO22X1 U465 ( .IN1(n352), .IN2(Acc[3]), .IN3(n343), .IN4(Acc[4]), .Q(n395)
         );
  AO221X1 U466 ( .IN1(case_add[37]), .IN2(n346), .IN3(case_sub[37]), .IN4(n349), .IN5(n395), .Q(n180) );
  AO22X1 U467 ( .IN1(n353), .IN2(Acc[2]), .IN3(n343), .IN4(Acc[3]), .Q(n396)
         );
  AO221X1 U468 ( .IN1(case_add[36]), .IN2(n346), .IN3(case_sub[36]), .IN4(n349), .IN5(n396), .Q(n179) );
  AO22X1 U469 ( .IN1(n352), .IN2(n398), .IN3(n343), .IN4(Acc[2]), .Q(n397) );
  AO221X1 U470 ( .IN1(case_add[35]), .IN2(n346), .IN3(case_sub[35]), .IN4(n349), .IN5(n397), .Q(n178) );
  AO22X1 U471 ( .IN1(n352), .IN2(n320), .IN3(n341), .IN4(n398), .Q(n399) );
  AO221X1 U472 ( .IN1(case_add[34]), .IN2(n344), .IN3(case_sub[34]), .IN4(n349), .IN5(n399), .Q(n242) );
  MUX21X1 U473 ( .IN1(M_reg[31]), .IN2(M[31]), .S(n362), .Q(n280) );
  MUX21X1 U474 ( .IN1(M_reg[30]), .IN2(M[30]), .S(n362), .Q(n279) );
  MUX21X1 U475 ( .IN1(M_reg[29]), .IN2(M[29]), .S(n362), .Q(n278) );
  MUX21X1 U476 ( .IN1(M_reg[28]), .IN2(M[28]), .S(n362), .Q(n277) );
  MUX21X1 U477 ( .IN1(M_reg[27]), .IN2(M[27]), .S(n362), .Q(n276) );
  MUX21X1 U478 ( .IN1(M_reg[26]), .IN2(M[26]), .S(n362), .Q(n275) );
  MUX21X1 U479 ( .IN1(M_reg[25]), .IN2(M[25]), .S(n362), .Q(n274) );
  MUX21X1 U480 ( .IN1(M_reg[24]), .IN2(M[24]), .S(n362), .Q(n273) );
  MUX21X1 U481 ( .IN1(M_reg[23]), .IN2(M[23]), .S(n362), .Q(n272) );
  MUX21X1 U482 ( .IN1(M_reg[22]), .IN2(M[22]), .S(n362), .Q(n271) );
  MUX21X1 U483 ( .IN1(M_reg[21]), .IN2(M[21]), .S(n362), .Q(n270) );
  MUX21X1 U484 ( .IN1(M_reg[20]), .IN2(M[20]), .S(n362), .Q(n269) );
  MUX21X1 U485 ( .IN1(M_reg[19]), .IN2(M[19]), .S(n362), .Q(n268) );
  MUX21X1 U486 ( .IN1(M_reg[18]), .IN2(M[18]), .S(n362), .Q(n267) );
  MUX21X1 U487 ( .IN1(M_reg[8]), .IN2(M[8]), .S(rst), .Q(n257) );
  MUX21X1 U488 ( .IN1(n337), .IN2(M[5]), .S(rst), .Q(n254) );
  MUX21X1 U489 ( .IN1(M_reg[1]), .IN2(M[1]), .S(rst), .Q(n250) );
  MUX21X1 U490 ( .IN1(M_reg[0]), .IN2(M[0]), .S(rst), .Q(n249) );
  AO21X1 U491 ( .IN1(n352), .IN2(n299), .IN3(n400), .Q(n208) );
  AO222X1 U492 ( .IN1(case_sub[33]), .IN2(n349), .IN3(case_add[33]), .IN4(n344), .IN5(n341), .IN6(n320), .Q(n401) );
  AO221X1 U493 ( .IN1(n352), .IN2(n315), .IN3(Q[31]), .IN4(n362), .IN5(n401), 
        .Q(n241) );
  NOR2X0 U494 ( .IN1(count[1]), .IN2(count[0]), .QN(n403) );
  AO21X1 U495 ( .IN1(count[1]), .IN2(count[0]), .IN3(n403), .Q(N110) );
  NOR2X0 U496 ( .IN1(n407), .IN2(count[2]), .QN(n404) );
  AO21X1 U497 ( .IN1(count[2]), .IN2(n407), .IN3(n404), .Q(N111) );
  NOR2X0 U498 ( .IN1(n408), .IN2(count[3]), .QN(n405) );
  AO21X1 U499 ( .IN1(count[3]), .IN2(n408), .IN3(n405), .Q(N112) );
  XNOR2X1 U500 ( .IN1(count[4]), .IN2(n409), .Q(N113) );
  NOR2X0 U501 ( .IN1(count[4]), .IN2(n409), .QN(n406) );
  XOR2X1 U502 ( .IN1(count[5]), .IN2(n406), .Q(N114) );
  OR3X1 U503 ( .IN1(count[5]), .IN2(count[4]), .IN3(count[3]), .Q(n410) );
endmodule

