
module BoothMultiplier_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387;

  OR2X1 U3 ( .IN1(n58), .IN2(n325), .Q(n57) );
  AND2X1 U4 ( .IN1(n365), .IN2(n366), .Q(n39) );
  AND2X1 U5 ( .IN1(n214), .IN2(n213), .Q(n33) );
  NAND4X0 U6 ( .IN1(A[4]), .IN2(n150), .IN3(n157), .IN4(n166), .QN(n100) );
  OR2X1 U7 ( .IN1(A[1]), .IN2(n377), .Q(n192) );
  OR2X1 U8 ( .IN1(A[5]), .IN2(n384), .Q(n157) );
  NBUFFX2 U9 ( .INP(n150), .Z(n63) );
  AND2X1 U10 ( .IN1(n138), .IN2(n358), .Q(n14) );
  NBUFFX2 U11 ( .INP(n24), .Z(n30) );
  AND2X1 U12 ( .IN1(n324), .IN2(n57), .Q(n49) );
  AND2X1 U13 ( .IN1(n31), .IN2(n231), .Q(n22) );
  AND2X1 U14 ( .IN1(n168), .IN2(n169), .Q(n114) );
  OR2X1 U15 ( .IN1(n28), .IN2(n325), .Q(n27) );
  AND2X1 U16 ( .IN1(n33), .IN2(n208), .Q(n106) );
  OR2X1 U17 ( .IN1(n249), .IN2(n250), .Q(n1) );
  AND4X1 U18 ( .IN1(n324), .IN2(n325), .IN3(n302), .IN4(n303), .Q(n2) );
  AND2X1 U19 ( .IN1(A[11]), .IN2(n357), .Q(n3) );
  AND2X1 U20 ( .IN1(n314), .IN2(n338), .Q(n4) );
  AND2X1 U21 ( .IN1(n138), .IN2(n360), .Q(n5) );
  NOR2X0 U22 ( .IN1(n51), .IN2(n112), .QN(n6) );
  AO221X1 U23 ( .IN1(n56), .IN2(n41), .IN3(n101), .IN4(n130), .IN5(n112), .Q(
        n35) );
  AND2X1 U24 ( .IN1(n33), .IN2(n204), .Q(n130) );
  AO22X1 U25 ( .IN1(n306), .IN2(n65), .IN3(n163), .IN4(n8), .Q(n141) );
  AO21X1 U26 ( .IN1(n348), .IN2(n67), .IN3(n323), .Q(n341) );
  AO22X1 U27 ( .IN1(n341), .IN2(n342), .IN3(B[12]), .IN4(n354), .Q(n338) );
  AND4X1 U28 ( .IN1(n311), .IN2(n318), .IN3(n319), .IN4(n312), .Q(n295) );
  AO21X1 U29 ( .IN1(n295), .IN2(n296), .IN3(n1), .Q(n41) );
  AO21X1 U30 ( .IN1(n88), .IN2(n89), .IN3(n7), .Q(n214) );
  INVX0 U31 ( .INP(n209), .ZN(n7) );
  AO21X1 U32 ( .IN1(n295), .IN2(n296), .IN3(n1), .Q(n248) );
  NOR2X0 U33 ( .IN1(n379), .IN2(n378), .QN(n8) );
  AND2X1 U34 ( .IN1(n274), .IN2(n275), .Q(n9) );
  NAND2X0 U35 ( .IN1(n90), .IN2(n230), .QN(n10) );
  NAND2X0 U36 ( .IN1(n360), .IN2(n14), .QN(n11) );
  AND2X1 U37 ( .IN1(n11), .IN2(n12), .Q(n355) );
  OR2X1 U38 ( .IN1(n13), .IN2(n30), .Q(n12) );
  INVX0 U39 ( .INP(n358), .ZN(n13) );
  OR2X1 U40 ( .IN1(A[1]), .IN2(n377), .Q(n15) );
  OR2X2 U41 ( .IN1(A[2]), .IN2(n375), .Q(n173) );
  INVX0 U42 ( .INP(n173), .ZN(n16) );
  NAND2X0 U43 ( .IN1(n10), .IN2(n20), .QN(n17) );
  NAND2X0 U44 ( .IN1(n17), .IN2(n18), .QN(n207) );
  OR2X1 U45 ( .IN1(n19), .IN2(n209), .Q(n18) );
  INVX0 U46 ( .INP(n213), .ZN(n19) );
  AND2X1 U47 ( .IN1(n89), .IN2(n213), .Q(n20) );
  NAND2X0 U48 ( .IN1(n93), .IN2(n248), .QN(n21) );
  NAND2X0 U49 ( .IN1(n302), .IN2(n303), .QN(n301) );
  OR2X1 U50 ( .IN1(n320), .IN2(n302), .Q(n71) );
  NAND2X1 U51 ( .IN1(B[14]), .IN2(n333), .QN(n302) );
  NAND2X0 U52 ( .IN1(n31), .IN2(n23), .QN(n89) );
  NAND2X1 U53 ( .IN1(n229), .IN2(n84), .QN(n23) );
  NAND2X0 U54 ( .IN1(B[10]), .IN2(n347), .QN(n24) );
  NAND2X1 U55 ( .IN1(n238), .IN2(n239), .QN(n230) );
  AND2X1 U56 ( .IN1(A[24]), .IN2(n234), .Q(n32) );
  AND2X1 U57 ( .IN1(B[10]), .IN2(n347), .Q(n25) );
  OR2X1 U58 ( .IN1(A[24]), .IN2(n234), .Q(n221) );
  AND2X1 U59 ( .IN1(n387), .IN2(n73), .Q(n350) );
  NAND2X0 U60 ( .IN1(n338), .IN2(n29), .QN(n26) );
  AND2X1 U61 ( .IN1(n26), .IN2(n27), .Q(n330) );
  INVX0 U62 ( .INP(n300), .ZN(n28) );
  AND2X1 U63 ( .IN1(n314), .IN2(n300), .Q(n29) );
  NAND2X1 U64 ( .IN1(n39), .IN2(n310), .QN(n163) );
  OR2X1 U65 ( .IN1(n221), .IN2(n32), .Q(n31) );
  OR2X1 U66 ( .IN1(n166), .IN2(A[4]), .Q(n162) );
  NAND2X0 U67 ( .IN1(B[10]), .IN2(n347), .QN(n351) );
  NAND2X0 U68 ( .IN1(n146), .IN2(n148), .QN(n382) );
  AND2X1 U69 ( .IN1(n247), .IN2(n41), .Q(n34) );
  NAND2X0 U70 ( .IN1(n64), .IN2(n101), .QN(n36) );
  NOR2X0 U71 ( .IN1(n122), .IN2(A[6]), .QN(n37) );
  XOR3X1 U72 ( .IN1(n185), .IN2(B[29]), .IN3(n184), .Q(DIFF[29]) );
  NAND2X0 U73 ( .IN1(n33), .IN2(n204), .QN(n38) );
  XOR2X1 U74 ( .IN1(n331), .IN2(n330), .Q(DIFF[14]) );
  NAND2X0 U75 ( .IN1(n40), .IN2(n54), .QN(n199) );
  AND2X1 U76 ( .IN1(n55), .IN2(n6), .Q(n40) );
  NAND2X0 U77 ( .IN1(n125), .IN2(n45), .QN(n42) );
  NAND2X0 U78 ( .IN1(n42), .IN2(n43), .QN(n179) );
  OR2X1 U79 ( .IN1(n44), .IN2(n83), .Q(n43) );
  INVX0 U80 ( .INP(n81), .ZN(n44) );
  AND2X1 U81 ( .IN1(n126), .IN2(n81), .Q(n45) );
  NAND2X0 U82 ( .IN1(n50), .IN2(n49), .QN(n46) );
  NAND2X0 U83 ( .IN1(n46), .IN2(n47), .QN(n70) );
  OR2X1 U84 ( .IN1(n48), .IN2(n59), .Q(n47) );
  INVX0 U85 ( .INP(n57), .ZN(n48) );
  NAND2X0 U86 ( .IN1(n341), .IN2(n342), .QN(n50) );
  INVX0 U87 ( .INP(n200), .ZN(n51) );
  NAND2X0 U88 ( .IN1(n22), .IN2(n230), .QN(n52) );
  XOR3X1 U89 ( .IN1(A[28]), .IN2(n197), .IN3(n195), .Q(DIFF[28]) );
  AND2X1 U90 ( .IN1(n21), .IN2(n36), .Q(n125) );
  AND2X1 U91 ( .IN1(n61), .IN2(n177), .Q(n53) );
  NAND2X0 U92 ( .IN1(n41), .IN2(n56), .QN(n54) );
  OR2X1 U93 ( .IN1(n38), .IN2(n102), .Q(n55) );
  AND2X1 U94 ( .IN1(n247), .IN2(n130), .Q(n56) );
  INVX0 U95 ( .INP(n72), .ZN(n58) );
  AND2X1 U96 ( .IN1(n314), .IN2(n72), .Q(n59) );
  NAND2X0 U97 ( .IN1(n125), .IN2(n126), .QN(n60) );
  AND2X1 U98 ( .IN1(n95), .IN2(n103), .Q(n61) );
  NAND4X0 U99 ( .IN1(n324), .IN2(n325), .IN3(n302), .IN4(n303), .QN(n62) );
  NAND2X1 U100 ( .IN1(B[15]), .IN2(n328), .QN(n303) );
  NAND2X0 U101 ( .IN1(n172), .IN2(n173), .QN(n171) );
  OR2X1 U102 ( .IN1(n385), .IN2(A[7]), .Q(n145) );
  NAND2X0 U103 ( .IN1(n191), .IN2(n192), .QN(n190) );
  OR2X1 U104 ( .IN1(A[9]), .IN2(n386), .Q(n137) );
  NAND2X0 U105 ( .IN1(n64), .IN2(n101), .QN(n92) );
  AND2X1 U106 ( .IN1(n207), .IN2(n128), .Q(n64) );
  OR2X1 U107 ( .IN1(n357), .IN2(A[11]), .Q(n346) );
  OR2X1 U108 ( .IN1(A[8]), .IN2(n352), .Q(n142) );
  NAND2X0 U109 ( .IN1(B[7]), .IN2(n381), .QN(n65) );
  NAND2X0 U110 ( .IN1(B[4]), .IN2(n380), .QN(n66) );
  NOR2X0 U111 ( .IN1(n68), .IN2(n3), .QN(n67) );
  AND4X1 U112 ( .IN1(A[8]), .IN2(n345), .IN3(n137), .IN4(n352), .Q(n68) );
  NAND2X0 U113 ( .IN1(n346), .IN2(n24), .QN(n69) );
  AND2X1 U114 ( .IN1(n70), .IN2(n71), .Q(n326) );
  AND2X1 U115 ( .IN1(n300), .IN2(n329), .Q(n72) );
  NAND2X0 U116 ( .IN1(n66), .IN2(n160), .QN(n164) );
  NAND2X0 U117 ( .IN1(n377), .IN2(A[1]), .QN(n189) );
  NAND2X0 U118 ( .IN1(n156), .IN2(n157), .QN(n155) );
  INVX0 U119 ( .INP(n347), .ZN(n73) );
  AND2X1 U120 ( .IN1(n168), .IN2(n362), .Q(n74) );
  NAND2X0 U121 ( .IN1(n142), .IN2(n137), .QN(n75) );
  OR2X1 U122 ( .IN1(A[3]), .IN2(n372), .Q(n168) );
  NAND2X0 U123 ( .IN1(n65), .IN2(n306), .QN(n76) );
  NAND2X0 U124 ( .IN1(n348), .IN2(n67), .QN(n322) );
  NAND2X0 U125 ( .IN1(n162), .IN2(n157), .QN(n378) );
  OR2X1 U126 ( .IN1(A[0]), .IN2(n371), .Q(n269) );
  NOR2X0 U127 ( .IN1(n75), .IN2(n69), .QN(n77) );
  NOR2X0 U128 ( .IN1(n344), .IN2(n343), .QN(n305) );
  NAND2X0 U129 ( .IN1(n9), .IN2(n80), .QN(n78) );
  AND2X1 U130 ( .IN1(n78), .IN2(n79), .Q(n107) );
  OR2X1 U131 ( .IN1(n249), .IN2(n260), .Q(n79) );
  AND2X1 U132 ( .IN1(n261), .IN2(n252), .Q(n80) );
  OR2X1 U133 ( .IN1(n82), .IN2(n183), .Q(n81) );
  INVX0 U134 ( .INP(n182), .ZN(n82) );
  AND2X1 U135 ( .IN1(n193), .IN2(n182), .Q(n83) );
  NAND2X0 U136 ( .IN1(n234), .IN2(A[24]), .QN(n84) );
  NAND2X0 U137 ( .IN1(n52), .IN2(n89), .QN(n85) );
  NAND2X0 U138 ( .IN1(n91), .IN2(n86), .QN(n94) );
  AND2X1 U139 ( .IN1(n92), .IN2(n97), .Q(n86) );
  NAND2X0 U140 ( .IN1(n269), .IN2(n267), .QN(DIFF[0]) );
  NAND2X0 U141 ( .IN1(n269), .IN2(n15), .QN(n363) );
  NAND2X0 U142 ( .IN1(A[16]), .IN2(n294), .QN(n87) );
  XOR2X2 U143 ( .IN1(n174), .IN2(n175), .Q(DIFF[31]) );
  NAND2X0 U144 ( .IN1(n274), .IN2(n275), .QN(n262) );
  NAND2X0 U145 ( .IN1(n90), .IN2(n230), .QN(n88) );
  AND2X1 U146 ( .IN1(n31), .IN2(n231), .Q(n90) );
  NAND3X0 U147 ( .IN1(n192), .IN2(n173), .IN3(A[0]), .QN(n369) );
  NAND2X0 U148 ( .IN1(n366), .IN2(n365), .QN(n315) );
  NAND2X0 U149 ( .IN1(A[21]), .IN2(n254), .QN(n242) );
  NAND2X0 U150 ( .IN1(n282), .IN2(n283), .QN(n276) );
  NAND2X0 U151 ( .IN1(n93), .IN2(n248), .QN(n91) );
  AND2X1 U152 ( .IN1(n247), .IN2(n127), .Q(n93) );
  OR2X1 U153 ( .IN1(n96), .IN2(n193), .Q(n95) );
  INVX0 U154 ( .INP(n105), .ZN(n96) );
  AND2X1 U155 ( .IN1(n126), .IN2(n105), .Q(n97) );
  NAND2X0 U156 ( .IN1(A[28]), .IN2(n197), .QN(n193) );
  NAND2X0 U157 ( .IN1(n295), .IN2(n296), .QN(n98) );
  NAND2X0 U158 ( .IN1(n259), .IN2(n260), .QN(n251) );
  NAND2X0 U159 ( .IN1(n240), .IN2(n241), .QN(n238) );
  NAND2X0 U160 ( .IN1(n160), .IN2(n161), .QN(n156) );
  NAND2X0 U161 ( .IN1(n111), .IN2(n261), .QN(n250) );
  NAND2X0 U162 ( .IN1(n232), .IN2(n231), .QN(n222) );
  NAND2X0 U163 ( .IN1(n243), .IN2(n241), .QN(n233) );
  NAND2X0 U164 ( .IN1(n132), .IN2(n115), .QN(n131) );
  NAND2X0 U165 ( .IN1(n200), .IN2(n194), .QN(n115) );
  NAND2X0 U166 ( .IN1(n231), .IN2(n229), .QN(n235) );
  NAND2X0 U167 ( .IN1(A[23]), .IN2(n124), .QN(n229) );
  NAND2X0 U168 ( .IN1(B[27]), .IN2(n202), .QN(n200) );
  NAND2X0 U169 ( .IN1(A[27]), .IN2(n203), .QN(n198) );
  NAND2X0 U170 ( .IN1(B[18]), .IN2(n280), .QN(n275) );
  NAND2X0 U171 ( .IN1(B[21]), .IN2(n255), .QN(n243) );
  NAND2X0 U172 ( .IN1(A[18]), .IN2(n279), .QN(n277) );
  INVX0 U173 ( .INP(B[22]), .ZN(n123) );
  INVX0 U174 ( .INP(B[23]), .ZN(n124) );
  NAND2X0 U175 ( .IN1(B[20]), .IN2(n264), .QN(n252) );
  NAND2X0 U176 ( .IN1(B[19]), .IN2(n272), .QN(n261) );
  INVX0 U177 ( .INP(B[6]), .ZN(n122) );
  NAND2X0 U178 ( .IN1(n100), .IN2(n99), .QN(n306) );
  NOR2X0 U179 ( .IN1(n383), .IN2(n382), .QN(n99) );
  NAND2X0 U180 ( .IN1(n210), .IN2(n209), .QN(n101) );
  NAND2X0 U181 ( .IN1(n211), .IN2(n102), .QN(n208) );
  INVX0 U182 ( .INP(n101), .ZN(n102) );
  NAND2X0 U183 ( .IN1(B[25]), .IN2(n224), .QN(n209) );
  OR2X1 U184 ( .IN1(n104), .IN2(n182), .Q(n103) );
  INVX0 U185 ( .INP(n178), .ZN(n104) );
  AND2X1 U186 ( .IN1(n183), .IN2(n178), .Q(n105) );
  NAND2X0 U187 ( .IN1(n221), .IN2(n84), .QN(n225) );
  INVX0 U188 ( .INP(n221), .ZN(n108) );
  INVX0 U189 ( .INP(n163), .ZN(n165) );
  NOR2X0 U190 ( .IN1(n258), .IN2(n251), .QN(n257) );
  NOR2X0 U191 ( .IN1(n291), .IN2(n250), .QN(n258) );
  NOR2X0 U192 ( .IN1(n237), .IN2(n230), .QN(n236) );
  NOR2X0 U193 ( .IN1(n34), .IN2(n233), .QN(n237) );
  NOR2X0 U194 ( .IN1(n219), .IN2(n85), .QN(n218) );
  NOR2X0 U195 ( .IN1(n34), .IN2(n212), .QN(n219) );
  NAND2X0 U196 ( .IN1(n273), .IN2(n262), .QN(n270) );
  INVX0 U197 ( .INP(n191), .ZN(n265) );
  INVX0 U198 ( .INP(n136), .ZN(n135) );
  INVX0 U199 ( .INP(n141), .ZN(n140) );
  INVX0 U200 ( .INP(n50), .ZN(n340) );
  INVX0 U201 ( .INP(n156), .ZN(n159) );
  NOR2X0 U202 ( .IN1(n37), .IN2(n154), .QN(n383) );
  INVX0 U203 ( .INP(n212), .ZN(n210) );
  NOR2X0 U204 ( .IN1(n25), .IN2(n138), .QN(n349) );
  NOR2X0 U205 ( .IN1(n376), .IN2(n189), .QN(n373) );
  AND2X1 U206 ( .IN1(n253), .IN2(n107), .Q(n247) );
  NOR2X0 U207 ( .IN1(n323), .IN2(n62), .QN(n321) );
  INVX0 U208 ( .INP(n63), .ZN(n153) );
  INVX0 U209 ( .INP(n242), .ZN(n240) );
  NAND2X0 U210 ( .IN1(n9), .IN2(n261), .QN(n259) );
  NOR2X0 U211 ( .IN1(n374), .IN2(n373), .QN(n365) );
  INVX0 U212 ( .INP(n169), .ZN(n367) );
  NAND2X0 U213 ( .IN1(n230), .IN2(n231), .QN(n228) );
  INVX0 U214 ( .INP(A[10]), .ZN(n347) );
  NAND2X0 U215 ( .IN1(n168), .IN2(n362), .QN(n310) );
  NOR2X0 U216 ( .IN1(n363), .IN2(n16), .QN(n362) );
  NAND2X0 U217 ( .IN1(n313), .IN2(n2), .QN(n312) );
  INVX0 U218 ( .INP(n314), .ZN(n313) );
  NAND2X0 U219 ( .IN1(n154), .IN2(n155), .QN(n149) );
  NOR2X0 U220 ( .IN1(n300), .IN2(n301), .QN(n299) );
  NAND2X0 U221 ( .IN1(n228), .IN2(n229), .QN(n220) );
  NOR2X0 U222 ( .IN1(n34), .IN2(n222), .QN(n227) );
  NOR2X0 U223 ( .IN1(n320), .IN2(n332), .QN(n331) );
  INVX0 U224 ( .INP(n302), .ZN(n332) );
  NOR2X0 U225 ( .IN1(n152), .IN2(n153), .QN(n151) );
  INVX0 U226 ( .INP(n148), .ZN(n152) );
  INVX0 U227 ( .INP(n329), .ZN(n320) );
  NOR2X0 U228 ( .IN1(n188), .IN2(n16), .QN(n187) );
  INVX0 U229 ( .INP(n170), .ZN(n188) );
  NAND2X0 U230 ( .IN1(n143), .IN2(n361), .QN(n136) );
  NAND2X0 U231 ( .IN1(n142), .IN2(n141), .QN(n361) );
  INVX0 U232 ( .INP(n252), .ZN(n249) );
  NOR2X0 U233 ( .IN1(n323), .IN2(n3), .QN(n356) );
  INVX0 U234 ( .INP(n233), .ZN(n232) );
  OR2X1 U235 ( .IN1(n222), .IN2(n108), .Q(n212) );
  NAND2X0 U236 ( .IN1(n189), .IN2(n190), .QN(n172) );
  NAND2X0 U237 ( .IN1(n147), .IN2(n148), .QN(n144) );
  NAND2X0 U238 ( .IN1(n149), .IN2(n63), .QN(n147) );
  NAND2X0 U239 ( .IN1(n170), .IN2(n171), .QN(n167) );
  NAND2X0 U240 ( .IN1(n136), .IN2(n137), .QN(n360) );
  AND2X1 U241 ( .IN1(n303), .IN2(n308), .Q(n109) );
  NAND2X0 U242 ( .IN1(n66), .IN2(n163), .QN(n161) );
  AND2X1 U243 ( .IN1(n286), .IN2(n283), .Q(n110) );
  INVX0 U244 ( .INP(n346), .ZN(n323) );
  NAND2X1 U245 ( .IN1(n267), .IN2(n268), .QN(n191) );
  INVX0 U246 ( .INP(n269), .ZN(n268) );
  AND2X1 U247 ( .IN1(n110), .IN2(n275), .Q(n111) );
  NOR2X0 U248 ( .IN1(n129), .IN2(n205), .QN(n112) );
  NAND2X1 U249 ( .IN1(n205), .IN2(n204), .QN(n206) );
  AND2X1 U250 ( .IN1(n261), .IN2(n260), .Q(n113) );
  NAND2X1 U251 ( .IN1(n209), .IN2(n213), .QN(n217) );
  NAND2X1 U252 ( .IN1(n198), .IN2(n200), .QN(n201) );
  NAND2X0 U253 ( .IN1(n320), .IN2(n303), .QN(n319) );
  NAND2X0 U254 ( .IN1(n131), .IN2(n116), .QN(n128) );
  NAND2X0 U255 ( .IN1(n204), .IN2(n132), .QN(n116) );
  AND2X1 U256 ( .IN1(n241), .IN2(n239), .Q(n117) );
  AND2X1 U257 ( .IN1(n275), .IN2(n277), .Q(n118) );
  NAND2X0 U258 ( .IN1(n128), .IN2(n119), .QN(n126) );
  NAND2X0 U259 ( .IN1(n205), .IN2(n131), .QN(n119) );
  AND2X1 U260 ( .IN1(n283), .IN2(n284), .Q(n120) );
  NAND2X0 U261 ( .IN1(n157), .IN2(n154), .QN(n158) );
  NAND2X0 U262 ( .IN1(n137), .IN2(n138), .QN(n134) );
  NAND2X1 U263 ( .IN1(n142), .IN2(n143), .QN(n139) );
  NAND2X0 U264 ( .IN1(n324), .IN2(n314), .QN(n339) );
  NAND2X0 U265 ( .IN1(n300), .IN2(n325), .QN(n335) );
  NAND2X0 U266 ( .IN1(n189), .IN2(n15), .QN(n266) );
  NAND2X1 U267 ( .IN1(n252), .IN2(n253), .QN(n256) );
  AND2X1 U268 ( .IN1(n65), .IN2(n146), .Q(n121) );
  INVX0 U269 ( .INP(B[5]), .ZN(n384) );
  OR2X1 U270 ( .IN1(A[6]), .IN2(n122), .Q(n150) );
  INVX0 U271 ( .INP(B[28]), .ZN(n197) );
  INVX0 U272 ( .INP(B[16]), .ZN(n294) );
  NAND2X0 U273 ( .IN1(n142), .IN2(n137), .QN(n343) );
  NAND2X0 U274 ( .IN1(B[10]), .IN2(n347), .QN(n345) );
  NOR2X0 U275 ( .IN1(n349), .IN2(n350), .QN(n348) );
  INVX0 U276 ( .INP(B[17]), .ZN(n288) );
  INVX0 U277 ( .INP(A[4]), .ZN(n380) );
  OR2X1 U278 ( .IN1(n123), .IN2(A[22]), .Q(n241) );
  NAND2X1 U279 ( .IN1(A[30]), .IN2(n181), .QN(n177) );
  INVX0 U280 ( .INP(B[30]), .ZN(n181) );
  NAND2X1 U281 ( .IN1(A[29]), .IN2(n186), .QN(n182) );
  INVX0 U282 ( .INP(B[29]), .ZN(n186) );
  NOR2X0 U283 ( .IN1(n369), .IN2(n370), .QN(n368) );
  NAND2X0 U284 ( .IN1(B[17]), .IN2(n289), .QN(n283) );
  INVX0 U285 ( .INP(A[7]), .ZN(n381) );
  INVX0 U286 ( .INP(B[9]), .ZN(n386) );
  INVX0 U287 ( .INP(B[2]), .ZN(n375) );
  INVX0 U288 ( .INP(B[12]), .ZN(n353) );
  INVX0 U289 ( .INP(B[13]), .ZN(n337) );
  INVX0 U290 ( .INP(B[14]), .ZN(n334) );
  INVX0 U291 ( .INP(B[15]), .ZN(n327) );
  INVX0 U292 ( .INP(B[7]), .ZN(n385) );
  INVX0 U293 ( .INP(B[21]), .ZN(n254) );
  INVX0 U294 ( .INP(B[11]), .ZN(n357) );
  INVX0 U295 ( .INP(B[1]), .ZN(n377) );
  INVX0 U296 ( .INP(B[3]), .ZN(n372) );
  OR2X1 U297 ( .IN1(n124), .IN2(A[23]), .Q(n231) );
  INVX0 U298 ( .INP(A[19]), .ZN(n272) );
  INVX0 U299 ( .INP(A[18]), .ZN(n280) );
  INVX0 U300 ( .INP(A[28]), .ZN(n196) );
  INVX0 U301 ( .INP(A[29]), .ZN(n185) );
  INVX0 U302 ( .INP(A[30]), .ZN(n180) );
  INVX0 U303 ( .INP(A[25]), .ZN(n224) );
  NAND2X0 U304 ( .IN1(A[19]), .IN2(n271), .QN(n260) );
  INVX0 U305 ( .INP(B[19]), .ZN(n271) );
  NAND2X0 U306 ( .IN1(A[4]), .IN2(n166), .QN(n160) );
  NAND2X1 U307 ( .IN1(A[26]), .IN2(n215), .QN(n204) );
  INVX0 U308 ( .INP(B[26]), .ZN(n215) );
  NAND2X0 U309 ( .IN1(A[22]), .IN2(n123), .QN(n239) );
  INVX0 U310 ( .INP(B[27]), .ZN(n203) );
  INVX0 U311 ( .INP(B[24]), .ZN(n234) );
  NAND2X1 U312 ( .IN1(B[26]), .IN2(n216), .QN(n205) );
  INVX0 U313 ( .INP(A[26]), .ZN(n216) );
  NAND2X0 U314 ( .IN1(A[20]), .IN2(n263), .QN(n253) );
  INVX0 U315 ( .INP(B[20]), .ZN(n263) );
  NAND2X0 U316 ( .IN1(A[25]), .IN2(n223), .QN(n213) );
  INVX0 U317 ( .INP(B[25]), .ZN(n223) );
  NAND2X0 U318 ( .IN1(B[12]), .IN2(n354), .QN(n324) );
  NAND2X0 U319 ( .IN1(B[13]), .IN2(n336), .QN(n325) );
  INVX0 U320 ( .INP(A[20]), .ZN(n264) );
  INVX0 U321 ( .INP(A[27]), .ZN(n202) );
  INVX0 U322 ( .INP(B[18]), .ZN(n279) );
  XOR3X1 U323 ( .IN1(n180), .IN2(B[30]), .IN3(n179), .Q(DIFF[30]) );
  NAND2X0 U324 ( .IN1(B[28]), .IN2(n196), .QN(n194) );
  INVX0 U325 ( .INP(A[21]), .ZN(n255) );
  NAND2X1 U326 ( .IN1(B[30]), .IN2(n180), .QN(n178) );
  NAND2X1 U327 ( .IN1(B[29]), .IN2(n185), .QN(n183) );
  NAND2X0 U328 ( .IN1(B[16]), .IN2(n293), .QN(n286) );
  INVX0 U329 ( .INP(A[16]), .ZN(n293) );
  INVX0 U330 ( .INP(B[10]), .ZN(n387) );
  INVX0 U331 ( .INP(A[31]), .ZN(n176) );
  INVX0 U332 ( .INP(B[4]), .ZN(n166) );
  INVX0 U333 ( .INP(B[8]), .ZN(n352) );
  INVX0 U334 ( .INP(B[0]), .ZN(n371) );
  NAND2X0 U335 ( .IN1(n308), .IN2(n307), .QN(n297) );
  INVX0 U336 ( .INP(n98), .ZN(n291) );
  NAND2X0 U337 ( .IN1(A[8]), .IN2(n352), .QN(n143) );
  NAND2X0 U338 ( .IN1(n77), .IN2(n141), .QN(n342) );
  NAND2X0 U339 ( .IN1(n77), .IN2(n2), .QN(n304) );
  NOR2X0 U340 ( .IN1(n379), .IN2(n378), .QN(n309) );
  NAND2X0 U341 ( .IN1(n245), .IN2(n242), .QN(n244) );
  NAND2X0 U342 ( .IN1(n243), .IN2(n242), .QN(n246) );
  NOR2X0 U343 ( .IN1(n227), .IN2(n220), .QN(n226) );
  NAND2X0 U344 ( .IN1(n281), .IN2(n276), .QN(n278) );
  NAND2X0 U345 ( .IN1(A[0]), .IN2(n371), .QN(n267) );
  NOR2X0 U346 ( .IN1(n364), .IN2(n170), .QN(n374) );
  INVX0 U347 ( .INP(n168), .ZN(n364) );
  AND2X1 U348 ( .IN1(n207), .IN2(n128), .Q(n127) );
  NOR2X0 U349 ( .IN1(n76), .IN2(n304), .QN(n298) );
  INVX0 U350 ( .INP(n204), .ZN(n129) );
  NAND2X0 U351 ( .IN1(A[13]), .IN2(n337), .QN(n300) );
  INVX0 U352 ( .INP(A[13]), .ZN(n336) );
  NAND2X0 U353 ( .IN1(A[14]), .IN2(n334), .QN(n329) );
  INVX0 U354 ( .INP(A[14]), .ZN(n333) );
  NAND2X0 U355 ( .IN1(n384), .IN2(A[5]), .QN(n154) );
  NAND2X0 U356 ( .IN1(A[9]), .IN2(n386), .QN(n138) );
  INVX0 U357 ( .INP(A[12]), .ZN(n354) );
  NAND2X0 U358 ( .IN1(A[12]), .IN2(n353), .QN(n314) );
  INVX0 U359 ( .INP(A[15]), .ZN(n328) );
  NAND2X0 U360 ( .IN1(A[15]), .IN2(n327), .QN(n308) );
  NAND2X0 U361 ( .IN1(n375), .IN2(A[2]), .QN(n170) );
  NAND2X0 U362 ( .IN1(n122), .IN2(A[6]), .QN(n148) );
  NAND2X0 U363 ( .IN1(n351), .IN2(n346), .QN(n344) );
  INVX0 U364 ( .INP(A[17]), .ZN(n289) );
  NAND2X0 U365 ( .IN1(n276), .IN2(n277), .QN(n274) );
  OR2X1 U366 ( .IN1(n133), .IN2(n198), .Q(n132) );
  INVX0 U367 ( .INP(n194), .ZN(n133) );
  NOR2X0 U368 ( .IN1(n368), .IN2(n367), .QN(n366) );
  NAND2X0 U369 ( .IN1(n173), .IN2(n168), .QN(n376) );
  NAND2X0 U370 ( .IN1(A[3]), .IN2(n372), .QN(n169) );
  NAND2X0 U371 ( .IN1(n168), .IN2(n371), .QN(n370) );
  NAND2X0 U372 ( .IN1(n30), .IN2(n358), .QN(n359) );
  NAND2X0 U373 ( .IN1(n321), .IN2(n322), .QN(n318) );
  NOR2X0 U374 ( .IN1(n317), .IN2(n62), .QN(n316) );
  NAND2X0 U375 ( .IN1(n198), .IN2(n199), .QN(n195) );
  NAND2X0 U376 ( .IN1(n315), .IN2(n316), .QN(n311) );
  NAND2X0 U377 ( .IN1(n305), .IN2(n309), .QN(n317) );
  NAND2X0 U378 ( .IN1(A[7]), .IN2(n385), .QN(n146) );
  NAND2X0 U379 ( .IN1(n145), .IN2(n150), .QN(n379) );
  NAND2X0 U380 ( .IN1(A[17]), .IN2(n288), .QN(n284) );
  NAND2X0 U381 ( .IN1(n193), .IN2(n60), .QN(n184) );
  NAND2X0 U382 ( .IN1(n243), .IN2(n211), .QN(n245) );
  NAND2X0 U383 ( .IN1(n247), .IN2(n41), .QN(n211) );
  NAND2X0 U384 ( .IN1(n87), .IN2(n286), .QN(n292) );
  NAND2X0 U385 ( .IN1(n290), .IN2(n87), .QN(n287) );
  NAND2X0 U386 ( .IN1(n284), .IN2(n285), .QN(n282) );
  NAND2X0 U387 ( .IN1(A[16]), .IN2(n294), .QN(n285) );
  NAND2X0 U388 ( .IN1(n53), .IN2(n94), .QN(n174) );
  NAND2X0 U389 ( .IN1(n111), .IN2(n98), .QN(n273) );
  NAND2X0 U390 ( .IN1(n110), .IN2(n98), .QN(n281) );
  NAND2X0 U391 ( .IN1(n286), .IN2(n98), .QN(n290) );
  NAND2X0 U392 ( .IN1(n73), .IN2(n387), .QN(n358) );
  XOR2X1 U393 ( .IN1(n134), .IN2(n135), .Q(DIFF[9]) );
  XOR2X1 U394 ( .IN1(n139), .IN2(n140), .Q(DIFF[8]) );
  XOR2X1 U395 ( .IN1(n144), .IN2(n121), .Q(DIFF[7]) );
  XOR2X1 U396 ( .IN1(n149), .IN2(n151), .Q(DIFF[6]) );
  XOR2X1 U397 ( .IN1(n158), .IN2(n159), .Q(DIFF[5]) );
  XOR2X1 U398 ( .IN1(n164), .IN2(n165), .Q(DIFF[4]) );
  XOR2X1 U399 ( .IN1(n167), .IN2(n114), .Q(DIFF[3]) );
  XOR2X1 U400 ( .IN1(n176), .IN2(B[31]), .Q(n175) );
  XOR2X1 U401 ( .IN1(n172), .IN2(n187), .Q(DIFF[2]) );
  XOR2X1 U402 ( .IN1(n201), .IN2(n35), .Q(DIFF[27]) );
  XOR2X1 U403 ( .IN1(n206), .IN2(n106), .Q(DIFF[26]) );
  XOR2X1 U404 ( .IN1(n217), .IN2(n218), .Q(DIFF[25]) );
  XOR2X1 U405 ( .IN1(n225), .IN2(n226), .Q(DIFF[24]) );
  XOR2X1 U406 ( .IN1(n235), .IN2(n236), .Q(DIFF[23]) );
  XOR2X1 U407 ( .IN1(n244), .IN2(n117), .Q(DIFF[22]) );
  XOR2X1 U408 ( .IN1(n246), .IN2(n34), .Q(DIFF[21]) );
  XOR2X1 U409 ( .IN1(n256), .IN2(n257), .Q(DIFF[20]) );
  XOR2X1 U410 ( .IN1(n265), .IN2(n266), .Q(DIFF[1]) );
  XOR2X1 U411 ( .IN1(n270), .IN2(n113), .Q(DIFF[19]) );
  XOR2X1 U412 ( .IN1(n278), .IN2(n118), .Q(DIFF[18]) );
  XOR2X1 U413 ( .IN1(n287), .IN2(n120), .Q(DIFF[17]) );
  XOR2X1 U414 ( .IN1(n291), .IN2(n292), .Q(DIFF[16]) );
  NOR3X0 U415 ( .IN1(n297), .IN2(n298), .IN3(n299), .QN(n296) );
  NAND4X0 U416 ( .IN1(n77), .IN2(n74), .IN3(n2), .IN4(n8), .QN(n307) );
  XOR2X1 U417 ( .IN1(n109), .IN2(n326), .Q(DIFF[15]) );
  XOR2X1 U418 ( .IN1(n4), .IN2(n335), .Q(DIFF[13]) );
  XOR2X1 U419 ( .IN1(n339), .IN2(n340), .Q(DIFF[12]) );
  XOR2X1 U420 ( .IN1(n356), .IN2(n355), .Q(DIFF[11]) );
  XOR2X1 U421 ( .IN1(n359), .IN2(n5), .Q(DIFF[10]) );
endmodule


module BoothMultiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335;

  OR2X1 U2 ( .IN1(B[24]), .IN2(A[24]), .Q(n192) );
  NAND3X0 U3 ( .IN1(n294), .IN2(n295), .IN3(n296), .QN(n267) );
  INVX0 U4 ( .INP(B[31]), .ZN(n64) );
  OR2X1 U5 ( .IN1(A[10]), .IN2(B[10]), .Q(n85) );
  OR2X1 U6 ( .IN1(A[9]), .IN2(B[9]), .Q(n15) );
  AND2X1 U7 ( .IN1(n45), .IN2(n290), .Q(n110) );
  AND2X1 U8 ( .IN1(n285), .IN2(n280), .Q(n52) );
  NBUFFX2 U9 ( .INP(n171), .Z(n17) );
  NBUFFX2 U10 ( .INP(n144), .Z(n21) );
  AND2X1 U11 ( .IN1(n326), .IN2(n327), .Q(n125) );
  AND2X1 U12 ( .IN1(A[9]), .IN2(B[9]), .Q(n120) );
  NBUFFX2 U13 ( .INP(n15), .Z(n115) );
  NAND3X0 U14 ( .IN1(n110), .IN2(n125), .IN3(n23), .QN(n59) );
  OR2X1 U15 ( .IN1(B[16]), .IN2(A[16]), .Q(n238) );
  OR2X1 U16 ( .IN1(B[21]), .IN2(A[21]), .Q(n201) );
  AND2X1 U17 ( .IN1(n76), .IN2(n166), .Q(n69) );
  OR2X1 U18 ( .IN1(B[0]), .IN2(A[0]), .Q(n224) );
  AND2X1 U19 ( .IN1(n140), .IN2(n16), .Q(n143) );
  AND2X1 U20 ( .IN1(n297), .IN2(n109), .Q(n309) );
  OR2X1 U21 ( .IN1(n194), .IN2(n96), .Q(n195) );
  OR2X1 U22 ( .IN1(n189), .IN2(n94), .Q(n190) );
  AO22X1 U23 ( .IN1(A[28]), .IN2(B[28]), .IN3(n76), .IN4(n75), .Q(n84) );
  XOR2X1 U24 ( .IN1(n23), .IN2(n152), .Q(SUM[4]) );
  XOR2X1 U25 ( .IN1(n131), .IN2(n132), .Q(SUM[8]) );
  XOR2X1 U26 ( .IN1(n284), .IN2(n286), .Q(SUM[12]) );
  NAND2X0 U27 ( .IN1(n244), .IN2(n243), .QN(n1) );
  OR2X1 U28 ( .IN1(n219), .IN2(n48), .Q(n2) );
  AND2X1 U29 ( .IN1(n6), .IN2(n211), .Q(n3) );
  AND2X1 U30 ( .IN1(B[19]), .IN2(A[19]), .Q(n4) );
  AND2X1 U31 ( .IN1(n100), .IN2(n192), .Q(n5) );
  AND2X1 U32 ( .IN1(n99), .IN2(n218), .Q(n6) );
  NAND2X1 U33 ( .IN1(n47), .IN2(n213), .QN(n7) );
  AND2X1 U34 ( .IN1(n254), .IN2(n278), .Q(n8) );
  AND2X1 U35 ( .IN1(n185), .IN2(n186), .Q(n9) );
  AND2X1 U36 ( .IN1(n5), .IN2(n187), .Q(n10) );
  NAND2X1 U37 ( .IN1(n183), .IN2(n93), .QN(n11) );
  AND2X1 U38 ( .IN1(n224), .IN2(n223), .Q(SUM[0]) );
  NAND2X0 U39 ( .IN1(n320), .IN2(n321), .QN(n174) );
  NAND3X1 U40 ( .IN1(n11), .IN2(n91), .IN3(n89), .QN(n76) );
  NAND4X0 U41 ( .IN1(n297), .IN2(n295), .IN3(n111), .IN4(n294), .QN(n83) );
  AO21X1 U42 ( .IN1(n202), .IN2(n205), .IN3(n13), .Q(n199) );
  INVX0 U43 ( .INP(n204), .ZN(n13) );
  AND3X1 U44 ( .IN1(n245), .IN2(n251), .IN3(n246), .Q(n244) );
  AO21X1 U45 ( .IN1(n330), .IN2(n331), .IN3(n14), .Q(n312) );
  INVX0 U46 ( .INP(n112), .ZN(n14) );
  NAND4X0 U47 ( .IN1(n247), .IN2(n126), .IN3(n112), .IN4(n110), .QN(n246) );
  OR2X1 U48 ( .IN1(B[28]), .IN2(A[28]), .Q(n176) );
  AND4X1 U49 ( .IN1(n257), .IN2(n262), .IN3(n261), .IN4(n256), .Q(n243) );
  OAI21X1 U50 ( .IN1(n19), .IN2(n37), .IN3(n18), .QN(n40) );
  AO22X1 U51 ( .IN1(n22), .IN2(n3), .IN3(n7), .IN4(n2), .Q(n108) );
  AO21X1 U52 ( .IN1(n118), .IN2(n274), .IN3(n263), .Q(n271) );
  AO22X1 U53 ( .IN1(n212), .IN2(n3), .IN3(n7), .IN4(n2), .Q(n188) );
  INVX0 U54 ( .INP(n122), .ZN(n16) );
  OR2X1 U55 ( .IN1(A[7]), .IN2(B[7]), .Q(n248) );
  NAND2X0 U56 ( .IN1(n297), .IN2(n307), .QN(n302) );
  NAND2X1 U57 ( .IN1(n39), .IN2(n20), .QN(n18) );
  INVX0 U58 ( .INP(n187), .ZN(n19) );
  AND2X1 U59 ( .IN1(n199), .IN2(n187), .Q(n20) );
  OR2X1 U60 ( .IN1(n43), .IN2(n95), .Q(n200) );
  OR2X1 U61 ( .IN1(A[6]), .IN2(B[6]), .Q(n142) );
  NAND2X0 U62 ( .IN1(n244), .IN2(n243), .QN(n22) );
  NAND4X0 U63 ( .IN1(n316), .IN2(n315), .IN3(n314), .IN4(n155), .QN(n23) );
  XOR3X1 U64 ( .IN1(B[29]), .IN2(A[29]), .IN3(n84), .Q(SUM[29]) );
  NOR2X0 U65 ( .IN1(A[6]), .IN2(B[6]), .QN(n122) );
  NAND2X0 U66 ( .IN1(n186), .IN2(n27), .QN(n24) );
  NAND2X0 U67 ( .IN1(n24), .IN2(n25), .QN(n29) );
  OR2X1 U68 ( .IN1(n26), .IN2(n183), .Q(n25) );
  INVX0 U69 ( .INP(n182), .ZN(n26) );
  AND2X1 U70 ( .IN1(n185), .IN2(n182), .Q(n27) );
  NAND2X1 U71 ( .IN1(n287), .IN2(n288), .QN(n284) );
  AND2X1 U72 ( .IN1(n228), .IN2(n28), .Q(n219) );
  AND2X1 U73 ( .IN1(n229), .IN2(n218), .Q(n28) );
  AND2X1 U74 ( .IN1(n165), .IN2(n67), .Q(n30) );
  NAND2X0 U75 ( .IN1(n34), .IN2(n186), .QN(n31) );
  NAND2X0 U76 ( .IN1(n32), .IN2(n31), .QN(n179) );
  OR2X1 U77 ( .IN1(n33), .IN2(n58), .Q(n32) );
  INVX0 U78 ( .INP(n56), .ZN(n33) );
  AND2X1 U79 ( .IN1(n185), .IN2(n56), .Q(n34) );
  AND2X1 U80 ( .IN1(n77), .IN2(n72), .Q(n35) );
  NAND2X0 U81 ( .IN1(n199), .IN2(n39), .QN(n36) );
  NAND2X0 U82 ( .IN1(n36), .IN2(n37), .QN(n189) );
  OR2X1 U83 ( .IN1(n38), .IN2(n55), .Q(n37) );
  INVX0 U84 ( .INP(n53), .ZN(n38) );
  AND2X1 U85 ( .IN1(n196), .IN2(n53), .Q(n39) );
  NOR2X0 U86 ( .IN1(n40), .IN2(n41), .QN(n79) );
  OR2X1 U87 ( .IN1(n42), .IN2(n107), .Q(n41) );
  INVX0 U88 ( .INP(n89), .ZN(n42) );
  NAND2X0 U89 ( .IN1(n203), .IN2(n204), .QN(n43) );
  INVX0 U90 ( .INP(n159), .ZN(n44) );
  NOR2X0 U91 ( .IN1(A[3]), .IN2(B[3]), .QN(n119) );
  NOR2X0 U92 ( .IN1(A[11]), .IN2(B[11]), .QN(n123) );
  NOR2X0 U93 ( .IN1(n123), .IN2(n293), .QN(n45) );
  OR2X1 U94 ( .IN1(B[14]), .IN2(A[14]), .Q(n253) );
  NAND2X0 U95 ( .IN1(n10), .IN2(n188), .QN(n46) );
  INVX0 U96 ( .INP(n106), .ZN(n47) );
  OR2X1 U97 ( .IN1(n4), .IN2(n106), .Q(n48) );
  NAND2X0 U98 ( .IN1(n284), .IN2(n52), .QN(n49) );
  AND2X1 U99 ( .IN1(n49), .IN2(n50), .Q(n278) );
  OR2X1 U100 ( .IN1(n51), .IN2(n283), .Q(n50) );
  INVX0 U101 ( .INP(n280), .ZN(n51) );
  OR2X1 U102 ( .IN1(n54), .IN2(n192), .Q(n53) );
  INVX0 U103 ( .INP(n193), .ZN(n54) );
  AND2X1 U104 ( .IN1(n198), .IN2(n193), .Q(n55) );
  OR2X1 U105 ( .IN1(n57), .IN2(n182), .Q(n56) );
  INVX0 U106 ( .INP(n180), .ZN(n57) );
  AND2X1 U107 ( .IN1(n183), .IN2(n180), .Q(n58) );
  AND2X1 U108 ( .IN1(n59), .IN2(n60), .Q(n288) );
  OR2X1 U109 ( .IN1(n61), .IN2(n312), .Q(n60) );
  INVX0 U110 ( .INP(n110), .ZN(n61) );
  NAND2X0 U111 ( .IN1(n312), .IN2(n313), .QN(n131) );
  NAND2X0 U112 ( .IN1(n35), .IN2(n46), .QN(n62) );
  NAND2X0 U113 ( .IN1(n62), .IN2(n63), .QN(n65) );
  AND2X1 U114 ( .IN1(n70), .IN2(n73), .Q(n63) );
  NOR2X0 U115 ( .IN1(B[1]), .IN2(A[1]), .QN(n124) );
  XOR3X1 U116 ( .IN1(n64), .IN2(A[31]), .IN3(n65), .Q(SUM[31]) );
  OR2X1 U117 ( .IN1(A[5]), .IN2(B[5]), .Q(n147) );
  NAND2X0 U118 ( .IN1(n69), .IN2(n75), .QN(n66) );
  OR2X1 U119 ( .IN1(n68), .IN2(n175), .Q(n67) );
  INVX0 U120 ( .INP(n166), .ZN(n68) );
  OR2X1 U121 ( .IN1(n71), .IN2(n80), .Q(n70) );
  INVX0 U122 ( .INP(n160), .ZN(n71) );
  AND2X1 U123 ( .IN1(n82), .IN2(n160), .Q(n72) );
  OR2X1 U124 ( .IN1(n74), .IN2(n76), .Q(n73) );
  INVX0 U125 ( .INP(n72), .ZN(n74) );
  NAND2X0 U126 ( .IN1(n77), .IN2(n46), .QN(n75) );
  AND2X1 U127 ( .IN1(n79), .IN2(n91), .Q(n77) );
  AND2X1 U128 ( .IN1(n189), .IN2(n187), .Q(n78) );
  NAND2X1 U129 ( .IN1(n282), .IN2(n283), .QN(n279) );
  NAND2X0 U130 ( .IN1(B[21]), .IN2(A[21]), .QN(n206) );
  OR2X1 U131 ( .IN1(n81), .IN2(n88), .Q(n80) );
  INVX0 U132 ( .INP(n86), .ZN(n81) );
  AND2X1 U133 ( .IN1(n175), .IN2(n86), .Q(n82) );
  OR2X1 U134 ( .IN1(A[8]), .IN2(B[8]), .Q(n292) );
  NAND2X0 U135 ( .IN1(n10), .IN2(n188), .QN(n186) );
  OR2X1 U136 ( .IN1(n87), .IN2(n165), .Q(n86) );
  INVX0 U137 ( .INP(n161), .ZN(n87) );
  AND2X1 U138 ( .IN1(n166), .IN2(n161), .Q(n88) );
  OR2X1 U139 ( .IN1(n90), .IN2(n182), .Q(n89) );
  INVX0 U140 ( .INP(n93), .ZN(n90) );
  NAND2X0 U141 ( .IN1(n244), .IN2(n243), .QN(n212) );
  OR2X1 U142 ( .IN1(n92), .IN2(n178), .Q(n91) );
  INVX0 U143 ( .INP(n176), .ZN(n92) );
  AND2X1 U144 ( .IN1(n180), .IN2(n176), .Q(n93) );
  NAND2X0 U145 ( .IN1(B[28]), .IN2(A[28]), .QN(n175) );
  NAND2X0 U146 ( .IN1(B[27]), .IN2(A[27]), .QN(n178) );
  INVX0 U147 ( .INP(n108), .ZN(n209) );
  AND2X1 U148 ( .IN1(n108), .IN2(n5), .Q(n94) );
  AND2X1 U149 ( .IN1(n98), .IN2(n108), .Q(n95) );
  AND2X1 U150 ( .IN1(n108), .IN2(n100), .Q(n96) );
  NAND2X0 U151 ( .IN1(n125), .IN2(n23), .QN(n313) );
  NAND3X0 U152 ( .IN1(n322), .IN2(n159), .IN3(n323), .QN(n315) );
  NOR2X0 U153 ( .IN1(n107), .IN2(n78), .QN(n185) );
  INVX0 U154 ( .INP(n265), .ZN(n263) );
  AND2X1 U155 ( .IN1(n238), .IN2(n235), .Q(n97) );
  INVX0 U156 ( .INP(n156), .ZN(n170) );
  INVX0 U157 ( .INP(n218), .ZN(n220) );
  AND2X1 U158 ( .IN1(n201), .IN2(n202), .Q(n98) );
  AND2X1 U159 ( .IN1(n97), .IN2(n229), .Q(n99) );
  AND2X1 U160 ( .IN1(n98), .IN2(n196), .Q(n100) );
  INVX0 U161 ( .INP(n206), .ZN(n205) );
  NAND3X0 U162 ( .IN1(n85), .IN2(n15), .IN3(n299), .QN(n294) );
  NOR2X0 U163 ( .IN1(n254), .IN2(n255), .QN(n252) );
  NBUFFX2 U164 ( .INP(n85), .Z(n109) );
  NAND2X1 U165 ( .IN1(n173), .IN2(n174), .QN(n172) );
  NAND2X0 U166 ( .IN1(n208), .IN2(n206), .QN(n207) );
  INVX0 U167 ( .INP(n223), .ZN(n173) );
  NAND2X0 U168 ( .IN1(n254), .IN2(n278), .QN(n274) );
  INVX0 U169 ( .INP(n283), .ZN(n258) );
  NAND2X0 U170 ( .IN1(n130), .IN2(n310), .QN(n308) );
  NAND2X0 U171 ( .IN1(n149), .IN2(n150), .QN(n146) );
  NOR2X0 U172 ( .IN1(n273), .IN2(n255), .QN(n272) );
  INVX0 U173 ( .INP(n245), .ZN(n273) );
  NAND2X0 U174 ( .IN1(n156), .IN2(n157), .QN(n153) );
  NAND2X0 U175 ( .IN1(n158), .IN2(n159), .QN(n157) );
  NAND2X0 U176 ( .IN1(n135), .IN2(n311), .QN(n127) );
  NAND2X0 U177 ( .IN1(n201), .IN2(n206), .QN(n210) );
  NOR2X0 U178 ( .IN1(n133), .IN2(n134), .QN(n132) );
  INVX0 U179 ( .INP(n135), .ZN(n133) );
  AND2X1 U180 ( .IN1(n149), .IN2(n151), .Q(n152) );
  INVX0 U181 ( .INP(n211), .ZN(n213) );
  NOR2X0 U182 ( .IN1(n106), .IN2(n213), .QN(n216) );
  NOR2X0 U183 ( .IN1(n4), .IN2(n220), .QN(n226) );
  NOR2X0 U184 ( .IN1(n107), .IN2(n19), .QN(n191) );
  NAND2X1 U185 ( .IN1(n182), .IN2(n183), .QN(n184) );
  NAND2X1 U186 ( .IN1(n178), .IN2(n180), .QN(n181) );
  AND2X1 U187 ( .IN1(n204), .IN2(n202), .Q(n101) );
  AND2X1 U188 ( .IN1(n231), .IN2(n229), .Q(n102) );
  AND2X1 U189 ( .IN1(n198), .IN2(n196), .Q(n103) );
  AND2X1 U190 ( .IN1(n193), .IN2(n192), .Q(n104) );
  AND2X1 U191 ( .IN1(n112), .IN2(n138), .Q(n137) );
  AND2X1 U192 ( .IN1(n254), .IN2(n280), .Q(n281) );
  AND2X1 U193 ( .IN1(n21), .IN2(n113), .Q(n148) );
  NOR2X0 U194 ( .IN1(n258), .IN2(n270), .QN(n286) );
  AND2X1 U195 ( .IN1(n155), .IN2(n322), .Q(n154) );
  INVX0 U196 ( .INP(n295), .ZN(n304) );
  AND2X1 U197 ( .IN1(n236), .IN2(n235), .Q(n105) );
  OR2X1 U198 ( .IN1(A[4]), .IN2(B[4]), .Q(n151) );
  NAND2X1 U199 ( .IN1(B[29]), .IN2(A[29]), .QN(n165) );
  NAND2X1 U200 ( .IN1(n167), .IN2(n168), .QN(n166) );
  NAND2X1 U201 ( .IN1(B[30]), .IN2(A[30]), .QN(n160) );
  NAND2X1 U202 ( .IN1(n163), .IN2(n164), .QN(n161) );
  OR2X1 U203 ( .IN1(B[2]), .IN2(A[2]), .Q(n159) );
  OR2X1 U204 ( .IN1(B[18]), .IN2(A[18]), .Q(n229) );
  OR2X1 U205 ( .IN1(B[12]), .IN2(A[12]), .Q(n285) );
  OR2X1 U206 ( .IN1(B[13]), .IN2(A[13]), .Q(n280) );
  OR2X1 U207 ( .IN1(B[15]), .IN2(A[15]), .Q(n264) );
  OR2X1 U208 ( .IN1(B[17]), .IN2(A[17]), .Q(n235) );
  OR2X1 U209 ( .IN1(B[22]), .IN2(A[22]), .Q(n202) );
  OR2X1 U210 ( .IN1(B[19]), .IN2(A[19]), .Q(n218) );
  OR2X1 U211 ( .IN1(B[23]), .IN2(A[23]), .Q(n196) );
  NAND2X0 U212 ( .IN1(B[22]), .IN2(A[22]), .QN(n204) );
  AND2X1 U213 ( .IN1(B[20]), .IN2(A[20]), .Q(n106) );
  NAND2X0 U214 ( .IN1(B[26]), .IN2(A[26]), .QN(n182) );
  NAND2X0 U215 ( .IN1(B[24]), .IN2(A[24]), .QN(n193) );
  NAND2X0 U216 ( .IN1(B[23]), .IN2(A[23]), .QN(n198) );
  NAND2X0 U217 ( .IN1(B[18]), .IN2(A[18]), .QN(n231) );
  NAND2X0 U218 ( .IN1(B[4]), .IN2(n117), .QN(n149) );
  INVX0 U219 ( .INP(A[30]), .ZN(n164) );
  INVX0 U220 ( .INP(A[29]), .ZN(n168) );
  OR2X1 U221 ( .IN1(B[25]), .IN2(A[25]), .Q(n187) );
  AND2X1 U222 ( .IN1(B[25]), .IN2(A[25]), .Q(n107) );
  XOR3X1 U223 ( .IN1(B[30]), .IN2(A[30]), .IN3(n162), .Q(SUM[30]) );
  XOR3X1 U224 ( .IN1(B[28]), .IN2(A[28]), .IN3(n177), .Q(SUM[28]) );
  OR2X1 U225 ( .IN1(B[26]), .IN2(A[26]), .Q(n183) );
  OR2X1 U226 ( .IN1(B[27]), .IN2(A[27]), .Q(n180) );
  OR2X1 U227 ( .IN1(B[20]), .IN2(A[20]), .Q(n211) );
  INVX0 U228 ( .INP(B[30]), .ZN(n163) );
  INVX0 U229 ( .INP(B[29]), .ZN(n167) );
  INVX0 U230 ( .INP(B[5]), .ZN(n332) );
  INVX0 U231 ( .INP(B[8]), .ZN(n301) );
  INVX0 U232 ( .INP(B[14]), .ZN(n276) );
  INVX0 U233 ( .INP(B[7]), .ZN(n328) );
  INVX0 U234 ( .INP(n22), .ZN(n241) );
  NAND2X0 U235 ( .IN1(n151), .IN2(n23), .QN(n150) );
  NAND2X0 U236 ( .IN1(n267), .IN2(n266), .QN(n287) );
  OR2X1 U237 ( .IN1(A[9]), .IN2(B[9]), .Q(n291) );
  NOR2X0 U238 ( .IN1(B[2]), .IN2(A[2]), .QN(n121) );
  NAND2X0 U239 ( .IN1(n21), .IN2(n145), .QN(n141) );
  AND2X1 U240 ( .IN1(n297), .IN2(n111), .Q(n296) );
  NAND2X0 U241 ( .IN1(n298), .IN2(n120), .QN(n111) );
  NAND2X0 U242 ( .IN1(n289), .IN2(n290), .QN(n250) );
  NAND2X0 U243 ( .IN1(n328), .IN2(n329), .QN(n112) );
  INVX0 U244 ( .INP(A[7]), .ZN(n329) );
  NAND2X0 U245 ( .IN1(n332), .IN2(n333), .QN(n113) );
  NAND2X0 U246 ( .IN1(n332), .IN2(n333), .QN(n114) );
  INVX0 U247 ( .INP(A[4]), .ZN(n116) );
  INVX0 U248 ( .INP(n116), .ZN(n117) );
  NOR2X0 U249 ( .IN1(n219), .IN2(n4), .QN(n214) );
  NAND2X0 U250 ( .IN1(n276), .IN2(n277), .QN(n118) );
  INVX0 U251 ( .INP(n120), .ZN(n130) );
  NOR2X0 U252 ( .IN1(n120), .IN2(n129), .QN(n128) );
  NAND2X0 U253 ( .IN1(n139), .IN2(n140), .QN(n136) );
  NAND2X0 U254 ( .IN1(n138), .IN2(n140), .QN(n334) );
  NAND2X0 U255 ( .IN1(B[6]), .IN2(A[6]), .QN(n140) );
  NAND2X0 U256 ( .IN1(n263), .IN2(n264), .QN(n262) );
  INVX0 U257 ( .INP(n264), .ZN(n255) );
  INVX0 U258 ( .INP(B[3]), .ZN(n324) );
  INVX0 U259 ( .INP(n292), .ZN(n134) );
  NAND2X0 U260 ( .IN1(n292), .IN2(n131), .QN(n311) );
  NAND2X0 U261 ( .IN1(n284), .IN2(n285), .QN(n282) );
  INVX0 U262 ( .INP(n285), .ZN(n270) );
  NAND2X0 U263 ( .IN1(B[17]), .IN2(A[17]), .QN(n236) );
  NOR2X0 U264 ( .IN1(n123), .IN2(n304), .QN(n303) );
  NOR2X0 U265 ( .IN1(n123), .IN2(n293), .QN(n289) );
  NAND2X0 U266 ( .IN1(n17), .IN2(n172), .QN(n158) );
  NAND2X0 U267 ( .IN1(n174), .IN2(n17), .QN(n222) );
  INVX0 U268 ( .INP(n171), .ZN(n323) );
  NAND2X0 U269 ( .IN1(B[1]), .IN2(A[1]), .QN(n171) );
  NAND2X0 U270 ( .IN1(B[0]), .IN2(A[0]), .QN(n319) );
  NAND2X0 U271 ( .IN1(B[0]), .IN2(A[0]), .QN(n223) );
  OR2X1 U272 ( .IN1(A[10]), .IN2(B[10]), .Q(n298) );
  NAND2X0 U273 ( .IN1(n308), .IN2(n109), .QN(n307) );
  NAND2X0 U274 ( .IN1(n324), .IN2(n325), .QN(n322) );
  NAND2X0 U275 ( .IN1(n146), .IN2(n114), .QN(n145) );
  AND2X1 U276 ( .IN1(n151), .IN2(n147), .Q(n327) );
  NAND2X0 U277 ( .IN1(n197), .IN2(n198), .QN(n194) );
  NAND2X0 U278 ( .IN1(n141), .IN2(n16), .QN(n139) );
  AND2X1 U279 ( .IN1(n142), .IN2(n248), .Q(n326) );
  INVX0 U280 ( .INP(n115), .ZN(n129) );
  NAND2X0 U281 ( .IN1(n115), .IN2(n127), .QN(n310) );
  AND2X1 U282 ( .IN1(n292), .IN2(n291), .Q(n290) );
  NAND2X0 U283 ( .IN1(n170), .IN2(n322), .QN(n314) );
  NAND2X0 U284 ( .IN1(n252), .IN2(n118), .QN(n251) );
  NAND2X0 U285 ( .IN1(n118), .IN2(n265), .QN(n275) );
  AND2X1 U286 ( .IN1(n264), .IN2(n253), .Q(n269) );
  INVX0 U287 ( .INP(B[11]), .ZN(n305) );
  NAND2X0 U288 ( .IN1(n227), .IN2(n221), .QN(n225) );
  NAND2X0 U289 ( .IN1(n228), .IN2(n229), .QN(n221) );
  INVX0 U290 ( .INP(B[1]), .ZN(n320) );
  NOR2X0 U291 ( .IN1(n170), .IN2(n44), .QN(n169) );
  AND2X1 U292 ( .IN1(n280), .IN2(n285), .Q(n268) );
  NAND2X0 U293 ( .IN1(n305), .IN2(n306), .QN(n266) );
  NAND2X0 U294 ( .IN1(n327), .IN2(n326), .QN(n249) );
  INVX0 U295 ( .INP(A[3]), .ZN(n325) );
  AND2X1 U296 ( .IN1(n268), .IN2(n269), .Q(n126) );
  NAND2X0 U297 ( .IN1(n233), .IN2(n230), .QN(n232) );
  NAND2X0 U298 ( .IN1(n231), .IN2(n230), .QN(n228) );
  NAND2X0 U299 ( .IN1(n234), .IN2(n235), .QN(n230) );
  NOR2X0 U300 ( .IN1(n119), .IN2(n121), .QN(n317) );
  NOR2X0 U301 ( .IN1(n319), .IN2(n124), .QN(n318) );
  NAND2X0 U302 ( .IN1(B[13]), .IN2(A[13]), .QN(n254) );
  INVX0 U303 ( .INP(A[14]), .ZN(n277) );
  NAND2X0 U304 ( .IN1(B[14]), .IN2(A[14]), .QN(n265) );
  NAND2X0 U305 ( .IN1(B[5]), .IN2(A[5]), .QN(n144) );
  INVX0 U306 ( .INP(A[5]), .ZN(n333) );
  NOR2X0 U307 ( .IN1(n300), .IN2(n301), .QN(n299) );
  NAND2X0 U308 ( .IN1(B[12]), .IN2(A[12]), .QN(n283) );
  NAND2X0 U309 ( .IN1(B[15]), .IN2(A[15]), .QN(n245) );
  NOR2X0 U310 ( .IN1(n122), .IN2(n144), .QN(n335) );
  NAND2X0 U311 ( .IN1(n205), .IN2(n202), .QN(n203) );
  NAND2X0 U312 ( .IN1(n199), .IN2(n196), .QN(n197) );
  NAND2X0 U313 ( .IN1(B[2]), .IN2(A[2]), .QN(n156) );
  INVX0 U314 ( .INP(A[11]), .ZN(n306) );
  NAND2X0 U315 ( .IN1(B[11]), .IN2(A[11]), .QN(n295) );
  NAND2X0 U316 ( .IN1(n258), .IN2(n126), .QN(n257) );
  INVX0 U317 ( .INP(A[1]), .ZN(n321) );
  NAND2X0 U318 ( .IN1(n331), .IN2(n330), .QN(n247) );
  NOR2X0 U319 ( .IN1(n335), .IN2(n334), .QN(n330) );
  NAND2X0 U320 ( .IN1(n317), .IN2(n318), .QN(n316) );
  NOR2X0 U321 ( .IN1(n249), .IN2(n250), .QN(n259) );
  NAND2X0 U322 ( .IN1(n214), .IN2(n217), .QN(n215) );
  NAND2X0 U323 ( .IN1(n237), .IN2(n238), .QN(n242) );
  NAND2X0 U324 ( .IN1(n240), .IN2(n237), .QN(n239) );
  NAND2X0 U325 ( .IN1(n236), .IN2(n237), .QN(n234) );
  NAND2X0 U326 ( .IN1(B[16]), .IN2(A[16]), .QN(n237) );
  INVX0 U327 ( .INP(A[8]), .ZN(n300) );
  NAND2X0 U328 ( .IN1(B[8]), .IN2(A[8]), .QN(n135) );
  NAND2X0 U329 ( .IN1(n66), .IN2(n30), .QN(n162) );
  NAND2X0 U330 ( .IN1(B[3]), .IN2(A[3]), .QN(n155) );
  NAND2X0 U331 ( .IN1(B[7]), .IN2(A[7]), .QN(n138) );
  NAND2X0 U332 ( .IN1(n6), .IN2(n1), .QN(n217) );
  NAND2X0 U333 ( .IN1(n97), .IN2(n1), .QN(n233) );
  NAND2X0 U334 ( .IN1(n238), .IN2(n22), .QN(n240) );
  NAND2X0 U335 ( .IN1(n99), .IN2(n1), .QN(n227) );
  NAND2X0 U336 ( .IN1(B[10]), .IN2(A[10]), .QN(n297) );
  NOR2X0 U337 ( .IN1(A[10]), .IN2(B[10]), .QN(n293) );
  NAND2X0 U338 ( .IN1(n178), .IN2(n179), .QN(n177) );
  NAND2X0 U339 ( .IN1(n201), .IN2(n108), .QN(n208) );
  XOR2X1 U340 ( .IN1(n127), .IN2(n128), .Q(SUM[9]) );
  XOR2X1 U341 ( .IN1(n136), .IN2(n137), .Q(SUM[7]) );
  XOR2X1 U342 ( .IN1(n141), .IN2(n143), .Q(SUM[6]) );
  XOR2X1 U343 ( .IN1(n146), .IN2(n148), .Q(SUM[5]) );
  XOR2X1 U344 ( .IN1(n153), .IN2(n154), .Q(SUM[3]) );
  XOR2X1 U345 ( .IN1(n158), .IN2(n169), .Q(SUM[2]) );
  XOR2X1 U346 ( .IN1(n29), .IN2(n181), .Q(SUM[27]) );
  XOR2X1 U347 ( .IN1(n9), .IN2(n184), .Q(SUM[26]) );
  XOR2X1 U348 ( .IN1(n190), .IN2(n191), .Q(SUM[25]) );
  XOR2X1 U349 ( .IN1(n195), .IN2(n104), .Q(SUM[24]) );
  XOR2X1 U350 ( .IN1(n200), .IN2(n103), .Q(SUM[23]) );
  XOR2X1 U351 ( .IN1(n207), .IN2(n101), .Q(SUM[22]) );
  XOR2X1 U352 ( .IN1(n209), .IN2(n210), .Q(SUM[21]) );
  XOR2X1 U353 ( .IN1(n216), .IN2(n215), .Q(SUM[20]) );
  XOR2X1 U354 ( .IN1(n222), .IN2(n223), .Q(SUM[1]) );
  XOR2X1 U355 ( .IN1(n226), .IN2(n225), .Q(SUM[19]) );
  XOR2X1 U356 ( .IN1(n102), .IN2(n232), .Q(SUM[18]) );
  XOR2X1 U357 ( .IN1(n105), .IN2(n239), .Q(SUM[17]) );
  XOR2X1 U358 ( .IN1(n241), .IN2(n242), .Q(SUM[16]) );
  NAND3X0 U359 ( .IN1(n259), .IN2(n126), .IN3(n260), .QN(n256) );
  NAND3X0 U360 ( .IN1(n83), .IN2(n266), .IN3(n126), .QN(n261) );
  XOR2X1 U361 ( .IN1(n272), .IN2(n271), .Q(SUM[15]) );
  XOR2X1 U362 ( .IN1(n8), .IN2(n275), .Q(SUM[14]) );
  XOR2X1 U363 ( .IN1(n279), .IN2(n281), .Q(SUM[13]) );
  XOR2X1 U364 ( .IN1(n302), .IN2(n303), .Q(SUM[11]) );
  XOR2X1 U365 ( .IN1(n308), .IN2(n309), .Q(SUM[10]) );
  NAND4X0 U366 ( .IN1(n316), .IN2(n315), .IN3(n314), .IN4(n155), .QN(n260) );
  NAND4X0 U367 ( .IN1(B[4]), .IN2(n117), .IN3(n114), .IN4(n142), .QN(n331) );
endmodule


module BoothMultiplier ( clk, oClk, rst, oRst, M, Q, P );
  input [31:0] M;
  input [31:0] Q;
  output [63:0] P;
  input clk, oClk, rst, oRst;
  wire   N4, N43, N44, N45, N46, N47, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n161, n164, n168, n171, n172, n173, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442;
  wire   [31:0] Acc;
  wire   [31:0] Q_reg;
  wire   [5:0] count;
  wire   [31:0] M_reg;
  wire   [64:33] case_add;
  wire   [64:33] case_sub;

  LATCHX1 \M_reg_reg[31]  ( .CLK(n382), .D(M[31]), .Q(M_reg[31]) );
  LATCHX1 \M_reg_reg[30]  ( .CLK(n382), .D(M[30]), .Q(M_reg[30]) );
  LATCHX1 \M_reg_reg[29]  ( .CLK(n382), .D(M[29]), .Q(M_reg[29]) );
  LATCHX1 \M_reg_reg[28]  ( .CLK(n382), .D(M[28]), .Q(M_reg[28]) );
  LATCHX1 \M_reg_reg[27]  ( .CLK(n382), .D(M[27]), .Q(M_reg[27]) );
  LATCHX1 \M_reg_reg[26]  ( .CLK(n382), .D(M[26]), .Q(M_reg[26]) );
  LATCHX1 \M_reg_reg[25]  ( .CLK(n382), .D(M[25]), .Q(M_reg[25]) );
  LATCHX1 \M_reg_reg[24]  ( .CLK(n382), .D(M[24]), .Q(M_reg[24]) );
  LATCHX1 \M_reg_reg[23]  ( .CLK(n382), .D(M[23]), .Q(M_reg[23]) );
  LATCHX1 \M_reg_reg[22]  ( .CLK(n382), .D(M[22]), .Q(M_reg[22]) );
  LATCHX1 \M_reg_reg[21]  ( .CLK(n382), .D(M[21]), .Q(M_reg[21]) );
  LATCHX1 \M_reg_reg[20]  ( .CLK(n382), .D(M[20]), .Q(M_reg[20]) );
  LATCHX1 \M_reg_reg[19]  ( .CLK(n382), .D(M[19]), .Q(M_reg[19]) );
  LATCHX1 \M_reg_reg[18]  ( .CLK(n382), .D(M[18]), .Q(M_reg[18]) );
  LATCHX1 \M_reg_reg[17]  ( .CLK(n382), .D(M[17]), .Q(M_reg[17]) );
  LATCHX1 \M_reg_reg[16]  ( .CLK(n382), .D(M[16]), .Q(M_reg[16]) );
  LATCHX1 \M_reg_reg[15]  ( .CLK(n382), .D(M[15]), .Q(M_reg[15]) );
  LATCHX1 \M_reg_reg[14]  ( .CLK(n382), .D(M[14]), .Q(M_reg[14]) );
  LATCHX1 \M_reg_reg[13]  ( .CLK(n382), .D(M[13]), .Q(M_reg[13]) );
  LATCHX1 \M_reg_reg[12]  ( .CLK(n382), .D(M[12]), .Q(M_reg[12]) );
  LATCHX1 \M_reg_reg[11]  ( .CLK(n382), .D(M[11]), .Q(M_reg[11]) );
  LATCHX1 \M_reg_reg[10]  ( .CLK(n382), .D(M[10]), .Q(M_reg[10]) );
  LATCHX1 \M_reg_reg[8]  ( .CLK(n382), .D(M[8]), .Q(M_reg[8]) );
  LATCHX1 \M_reg_reg[6]  ( .CLK(n381), .D(M[6]), .Q(M_reg[6]) );
  LATCHX1 \M_reg_reg[5]  ( .CLK(n381), .D(M[5]), .Q(M_reg[5]) );
  LATCHX1 \M_reg_reg[3]  ( .CLK(n381), .D(M[3]), .Q(M_reg[3]) );
  LATCHX1 \M_reg_reg[1]  ( .CLK(n381), .D(M[1]), .Q(M_reg[1]) );
  LATCHX1 \M_reg_reg[0]  ( .CLK(n381), .D(M[0]), .Q(M_reg[0]) );
  DFFARX1 \P_reg[63]  ( .D(Acc[31]), .CLK(n387), .RSTB(n366), .Q(P[63]) );
  DFFARX1 \P_reg[62]  ( .D(Acc[31]), .CLK(n387), .RSTB(n366), .Q(P[62]) );
  DFFARX1 \P_reg[61]  ( .D(Acc[30]), .CLK(n387), .RSTB(n366), .Q(P[61]) );
  DFFARX1 \P_reg[60]  ( .D(Acc[29]), .CLK(n387), .RSTB(n366), .Q(P[60]) );
  DFFARX1 \P_reg[59]  ( .D(Acc[28]), .CLK(n387), .RSTB(n365), .Q(P[59]) );
  DFFARX1 \P_reg[58]  ( .D(Acc[27]), .CLK(n387), .RSTB(n365), .Q(P[58]) );
  DFFARX1 \P_reg[57]  ( .D(Acc[26]), .CLK(n387), .RSTB(n365), .Q(P[57]) );
  DFFARX1 \P_reg[56]  ( .D(Acc[25]), .CLK(n387), .RSTB(n365), .Q(P[56]) );
  DFFARX1 \P_reg[55]  ( .D(n402), .CLK(n387), .RSTB(n365), .Q(P[55]) );
  DFFARX1 \P_reg[54]  ( .D(Acc[23]), .CLK(n387), .RSTB(n364), .Q(P[54]) );
  DFFARX1 \P_reg[53]  ( .D(Acc[22]), .CLK(n387), .RSTB(n364), .Q(P[53]) );
  DFFARX1 \P_reg[52]  ( .D(n406), .CLK(n387), .RSTB(n364), .Q(P[52]) );
  DFFARX1 \P_reg[51]  ( .D(Acc[20]), .CLK(n388), .RSTB(n364), .Q(P[51]) );
  DFFARX1 \P_reg[50]  ( .D(Acc[19]), .CLK(n388), .RSTB(n364), .Q(P[50]) );
  DFFARX1 \P_reg[49]  ( .D(Acc[18]), .CLK(n388), .RSTB(n363), .Q(P[49]) );
  DFFARX1 \P_reg[48]  ( .D(n411), .CLK(n388), .RSTB(n363), .Q(P[48]) );
  DFFARX1 \P_reg[47]  ( .D(Acc[16]), .CLK(n388), .RSTB(n363), .Q(P[47]) );
  DFFARX1 \P_reg[46]  ( .D(Acc[15]), .CLK(n388), .RSTB(n363), .Q(P[46]) );
  DFFARX1 \P_reg[45]  ( .D(Acc[14]), .CLK(n388), .RSTB(n363), .Q(P[45]) );
  DFFARX1 \P_reg[44]  ( .D(Acc[13]), .CLK(n388), .RSTB(n362), .Q(P[44]) );
  DFFARX1 \P_reg[43]  ( .D(Acc[12]), .CLK(n388), .RSTB(n362), .Q(P[43]) );
  DFFARX1 \P_reg[42]  ( .D(n317), .CLK(n388), .RSTB(n362), .Q(P[42]) );
  DFFARX1 \P_reg[41]  ( .D(n320), .CLK(n388), .RSTB(n362), .Q(P[41]) );
  DFFARX1 \P_reg[40]  ( .D(n319), .CLK(n388), .RSTB(n362), .Q(P[40]) );
  DFFARX1 \P_reg[39]  ( .D(n321), .CLK(n389), .RSTB(n361), .Q(P[39]) );
  DFFARX1 \P_reg[38]  ( .D(n340), .CLK(n389), .RSTB(n361), .Q(P[38]) );
  DFFARX1 \P_reg[37]  ( .D(n424), .CLK(n389), .RSTB(n361), .Q(P[37]) );
  DFFARX1 \P_reg[36]  ( .D(Acc[5]), .CLK(n389), .RSTB(n361), .Q(P[36]) );
  DFFARX1 \P_reg[35]  ( .D(n427), .CLK(n389), .RSTB(n361), .Q(P[35]) );
  DFFARX1 \P_reg[34]  ( .D(n324), .CLK(n389), .RSTB(n360), .Q(P[34]) );
  DFFARX1 \P_reg[33]  ( .D(Acc[2]), .CLK(n389), .RSTB(n360), .Q(P[33]) );
  DFFARX1 \P_reg[32]  ( .D(n325), .CLK(n389), .RSTB(n360), .Q(P[32]) );
  DFFARX1 \P_reg[31]  ( .D(n327), .CLK(n389), .RSTB(n360), .Q(P[31]) );
  DFFARX1 \P_reg[30]  ( .D(Q_reg[31]), .CLK(n389), .RSTB(n360), .Q(P[30]) );
  DFFARX1 \P_reg[29]  ( .D(Q_reg[30]), .CLK(n389), .RSTB(n359), .Q(P[29]) );
  DFFARX1 \P_reg[28]  ( .D(Q_reg[29]), .CLK(n389), .RSTB(n359), .Q(P[28]) );
  DFFARX1 \P_reg[27]  ( .D(Q_reg[28]), .CLK(n390), .RSTB(n359), .Q(P[27]) );
  DFFARX1 \P_reg[26]  ( .D(Q_reg[27]), .CLK(n390), .RSTB(n359), .Q(P[26]) );
  DFFARX1 \P_reg[25]  ( .D(Q_reg[26]), .CLK(n390), .RSTB(n359), .Q(P[25]) );
  DFFARX1 \P_reg[24]  ( .D(Q_reg[25]), .CLK(n390), .RSTB(n358), .Q(P[24]) );
  DFFARX1 \P_reg[23]  ( .D(Q_reg[24]), .CLK(n390), .RSTB(n358), .Q(P[23]) );
  DFFARX1 \P_reg[22]  ( .D(Q_reg[23]), .CLK(n390), .RSTB(n358), .Q(P[22]) );
  DFFARX1 \P_reg[21]  ( .D(Q_reg[22]), .CLK(n390), .RSTB(n358), .Q(P[21]) );
  DFFARX1 \P_reg[20]  ( .D(Q_reg[21]), .CLK(n390), .RSTB(n358), .Q(P[20]) );
  DFFARX1 \P_reg[19]  ( .D(Q_reg[20]), .CLK(n390), .RSTB(n357), .Q(P[19]) );
  DFFARX1 \P_reg[18]  ( .D(Q_reg[19]), .CLK(n390), .RSTB(n357), .Q(P[18]) );
  DFFARX1 \P_reg[17]  ( .D(Q_reg[18]), .CLK(n390), .RSTB(n357), .Q(P[17]) );
  DFFARX1 \P_reg[16]  ( .D(Q_reg[17]), .CLK(n390), .RSTB(n357), .Q(P[16]) );
  DFFARX1 \P_reg[15]  ( .D(Q_reg[16]), .CLK(n391), .RSTB(n357), .Q(P[15]) );
  DFFARX1 \P_reg[14]  ( .D(Q_reg[15]), .CLK(n391), .RSTB(n356), .Q(P[14]) );
  DFFARX1 \P_reg[13]  ( .D(Q_reg[14]), .CLK(n391), .RSTB(n356), .Q(P[13]) );
  DFFARX1 \P_reg[12]  ( .D(Q_reg[13]), .CLK(n391), .RSTB(n356), .Q(P[12]) );
  DFFARX1 \P_reg[11]  ( .D(Q_reg[12]), .CLK(n391), .RSTB(n356), .Q(P[11]) );
  DFFARX1 \P_reg[10]  ( .D(Q_reg[11]), .CLK(n391), .RSTB(n356), .Q(P[10]) );
  DFFARX1 \P_reg[9]  ( .D(Q_reg[10]), .CLK(n391), .RSTB(n355), .Q(P[9]) );
  DFFARX1 \P_reg[8]  ( .D(Q_reg[9]), .CLK(n391), .RSTB(n355), .Q(P[8]) );
  DFFARX1 \P_reg[7]  ( .D(Q_reg[8]), .CLK(n391), .RSTB(n355), .Q(P[7]) );
  DFFARX1 \P_reg[6]  ( .D(Q_reg[7]), .CLK(n391), .RSTB(n355), .Q(P[6]) );
  DFFARX1 \P_reg[5]  ( .D(Q_reg[6]), .CLK(n391), .RSTB(n355), .Q(P[5]) );
  DFFARX1 \P_reg[4]  ( .D(Q_reg[5]), .CLK(n391), .RSTB(n354), .Q(P[4]) );
  DFFARX1 \P_reg[3]  ( .D(Q_reg[4]), .CLK(n392), .RSTB(n354), .Q(P[3]) );
  DFFARX1 \P_reg[2]  ( .D(Q_reg[3]), .CLK(n392), .RSTB(n354), .Q(P[2]) );
  DFFARX1 \P_reg[1]  ( .D(Q_reg[2]), .CLK(n392), .RSTB(n354), .Q(P[1]) );
  DFFARX1 \P_reg[0]  ( .D(Q_reg[1]), .CLK(n392), .RSTB(n354), .Q(P[0]) );
  DFFASX1 \count_reg[0]  ( .D(n310), .CLK(clk), .SETB(n386), .Q(count[0]), 
        .QN(n314) );
  DFFARX1 \count_reg[5]  ( .D(n309), .CLK(clk), .RSTB(n384), .Q(count[5]), 
        .QN(n313) );
  DFFASX1 \count_reg[1]  ( .D(n308), .CLK(clk), .SETB(n386), .Q(count[1]), 
        .QN(n315) );
  DFFASX1 \count_reg[2]  ( .D(n307), .CLK(clk), .SETB(n386), .Q(count[2]) );
  DFFASX1 \count_reg[3]  ( .D(n306), .CLK(clk), .SETB(n386), .Q(count[3]) );
  DFFASX1 \count_reg[4]  ( .D(n305), .CLK(clk), .SETB(n386), .Q(count[4]) );
  DFFASRX1 \Q_reg_reg[0]  ( .D(n304), .CLK(clk), .RSTB(n238), .SETB(n237), .Q(
        n312), .QN(n173) );
  DFFARX1 Q_prev_reg ( .D(n303), .CLK(clk), .RSTB(n383), .Q(n172), .QN(n316)
         );
  DFFARX1 \Acc_reg[31]  ( .D(n302), .CLK(clk), .RSTB(n384), .Q(Acc[31]), .QN(
        n171) );
  DFFARX1 \Acc_reg[30]  ( .D(n301), .CLK(clk), .RSTB(n383), .Q(Acc[30]) );
  DFFARX1 \Acc_reg[29]  ( .D(n300), .CLK(clk), .RSTB(n383), .Q(Acc[29]) );
  DFFARX1 \Acc_reg[28]  ( .D(n299), .CLK(clk), .RSTB(n383), .Q(Acc[28]), .QN(
        n168) );
  DFFARX1 \Acc_reg[27]  ( .D(n298), .CLK(clk), .RSTB(n383), .Q(Acc[27]) );
  DFFARX1 \Acc_reg[26]  ( .D(n297), .CLK(clk), .RSTB(n383), .Q(Acc[26]) );
  DFFARX1 \Acc_reg[25]  ( .D(n296), .CLK(clk), .RSTB(n383), .Q(Acc[25]) );
  DFFARX1 \Acc_reg[24]  ( .D(n295), .CLK(clk), .RSTB(n383), .Q(Acc[24]), .QN(
        n164) );
  DFFARX1 \Acc_reg[23]  ( .D(n294), .CLK(clk), .RSTB(n383), .Q(Acc[23]) );
  DFFARX1 \Acc_reg[22]  ( .D(n293), .CLK(clk), .RSTB(n383), .Q(Acc[22]) );
  DFFARX1 \Acc_reg[21]  ( .D(n292), .CLK(clk), .RSTB(n383), .Q(Acc[21]), .QN(
        n161) );
  DFFARX1 \Acc_reg[20]  ( .D(n291), .CLK(clk), .RSTB(n383), .Q(Acc[20]) );
  DFFARX1 \Acc_reg[19]  ( .D(n290), .CLK(clk), .RSTB(n383), .Q(Acc[19]) );
  DFFARX1 \Acc_reg[18]  ( .D(n289), .CLK(clk), .RSTB(n385), .Q(Acc[18]) );
  DFFARX1 \Acc_reg[17]  ( .D(n288), .CLK(clk), .RSTB(n386), .Q(Acc[17]), .QN(
        n157) );
  DFFARX1 \Acc_reg[16]  ( .D(n287), .CLK(clk), .RSTB(n384), .Q(Acc[16]), .QN(
        n156) );
  DFFARX1 \Acc_reg[15]  ( .D(n286), .CLK(clk), .RSTB(n383), .Q(Acc[15]), .QN(
        n155) );
  DFFARX1 \Acc_reg[14]  ( .D(n285), .CLK(clk), .RSTB(n385), .Q(Acc[14]), .QN(
        n154) );
  DFFARX1 \Acc_reg[13]  ( .D(n284), .CLK(clk), .RSTB(n386), .Q(Acc[13]), .QN(
        n153) );
  DFFARX1 \Acc_reg[12]  ( .D(n283), .CLK(clk), .RSTB(n384), .Q(Acc[12]), .QN(
        n152) );
  DFFARX1 \Acc_reg[11]  ( .D(n282), .CLK(clk), .RSTB(n383), .Q(Acc[11]), .QN(
        n151) );
  DFFARX1 \Acc_reg[10]  ( .D(n281), .CLK(clk), .RSTB(n384), .Q(Acc[10]), .QN(
        n150) );
  DFFARX1 \Acc_reg[9]  ( .D(n280), .CLK(clk), .RSTB(n383), .Q(Acc[9]), .QN(
        n149) );
  DFFARX1 \Acc_reg[8]  ( .D(n279), .CLK(clk), .RSTB(n384), .Q(Acc[8]), .QN(
        n148) );
  DFFARX1 \Acc_reg[7]  ( .D(n278), .CLK(clk), .RSTB(n384), .Q(Acc[7]), .QN(
        n147) );
  DFFARX1 \Acc_reg[6]  ( .D(n277), .CLK(clk), .RSTB(n384), .Q(Acc[6]), .QN(
        n146) );
  DFFARX1 \Acc_reg[5]  ( .D(n276), .CLK(clk), .RSTB(n384), .Q(Acc[5]), .QN(
        n145) );
  DFFARX1 \Acc_reg[4]  ( .D(n275), .CLK(clk), .RSTB(n384), .Q(Acc[4]), .QN(
        n144) );
  DFFARX1 \Acc_reg[3]  ( .D(n274), .CLK(clk), .RSTB(n384), .Q(Acc[3]), .QN(
        n143) );
  DFFARX1 \Acc_reg[2]  ( .D(n273), .CLK(clk), .RSTB(n384), .Q(Acc[2]), .QN(
        n142) );
  DFFARX1 \Acc_reg[1]  ( .D(n272), .CLK(clk), .RSTB(n384), .Q(Acc[1]), .QN(
        n141) );
  DFFARX1 \Acc_reg[0]  ( .D(n271), .CLK(clk), .RSTB(n384), .Q(Acc[0]), .QN(
        n140) );
  DFFASRX1 \Q_reg_reg[31]  ( .D(n270), .CLK(clk), .RSTB(n236), .SETB(n235), 
        .Q(Q_reg[31]) );
  DFFASRX1 \Q_reg_reg[30]  ( .D(n269), .CLK(clk), .RSTB(n234), .SETB(n233), 
        .Q(Q_reg[30]) );
  DFFASRX1 \Q_reg_reg[29]  ( .D(n268), .CLK(clk), .RSTB(n232), .SETB(n231), 
        .Q(Q_reg[29]) );
  DFFASRX1 \Q_reg_reg[28]  ( .D(n267), .CLK(clk), .RSTB(n230), .SETB(n229), 
        .Q(Q_reg[28]) );
  DFFASRX1 \Q_reg_reg[27]  ( .D(n266), .CLK(clk), .RSTB(n228), .SETB(n227), 
        .Q(Q_reg[27]) );
  DFFASRX1 \Q_reg_reg[26]  ( .D(n265), .CLK(clk), .RSTB(n226), .SETB(n225), 
        .Q(Q_reg[26]) );
  DFFASRX1 \Q_reg_reg[25]  ( .D(n264), .CLK(clk), .RSTB(n224), .SETB(n223), 
        .Q(Q_reg[25]) );
  DFFASRX1 \Q_reg_reg[24]  ( .D(n263), .CLK(clk), .RSTB(n222), .SETB(n221), 
        .Q(Q_reg[24]) );
  DFFASRX1 \Q_reg_reg[23]  ( .D(n262), .CLK(clk), .RSTB(n220), .SETB(n219), 
        .Q(Q_reg[23]) );
  DFFASRX1 \Q_reg_reg[22]  ( .D(n261), .CLK(clk), .RSTB(n218), .SETB(n217), 
        .Q(Q_reg[22]) );
  DFFASRX1 \Q_reg_reg[21]  ( .D(n260), .CLK(clk), .RSTB(n216), .SETB(n215), 
        .Q(Q_reg[21]) );
  DFFASRX1 \Q_reg_reg[20]  ( .D(n259), .CLK(clk), .RSTB(n214), .SETB(n213), 
        .Q(Q_reg[20]) );
  DFFASRX1 \Q_reg_reg[19]  ( .D(n258), .CLK(clk), .RSTB(n212), .SETB(n211), 
        .Q(Q_reg[19]) );
  DFFASRX1 \Q_reg_reg[18]  ( .D(n257), .CLK(clk), .RSTB(n210), .SETB(n209), 
        .Q(Q_reg[18]) );
  DFFASRX1 \Q_reg_reg[17]  ( .D(n256), .CLK(clk), .RSTB(n208), .SETB(n207), 
        .Q(Q_reg[17]) );
  DFFASRX1 \Q_reg_reg[16]  ( .D(n255), .CLK(clk), .RSTB(n206), .SETB(n205), 
        .Q(Q_reg[16]) );
  DFFASRX1 \Q_reg_reg[15]  ( .D(n254), .CLK(clk), .RSTB(n204), .SETB(n203), 
        .Q(Q_reg[15]) );
  DFFASRX1 \Q_reg_reg[14]  ( .D(n253), .CLK(clk), .RSTB(n202), .SETB(n201), 
        .Q(Q_reg[14]) );
  DFFASRX1 \Q_reg_reg[13]  ( .D(n252), .CLK(clk), .RSTB(n200), .SETB(n199), 
        .Q(Q_reg[13]) );
  DFFASRX1 \Q_reg_reg[12]  ( .D(n251), .CLK(clk), .RSTB(n198), .SETB(n197), 
        .Q(Q_reg[12]) );
  DFFASRX1 \Q_reg_reg[11]  ( .D(n250), .CLK(clk), .RSTB(n196), .SETB(n195), 
        .Q(Q_reg[11]) );
  DFFASRX1 \Q_reg_reg[10]  ( .D(n249), .CLK(clk), .RSTB(n194), .SETB(n193), 
        .Q(Q_reg[10]) );
  DFFASRX1 \Q_reg_reg[9]  ( .D(n248), .CLK(clk), .RSTB(n192), .SETB(n191), .Q(
        Q_reg[9]) );
  DFFASRX1 \Q_reg_reg[8]  ( .D(n247), .CLK(clk), .RSTB(n190), .SETB(n189), .Q(
        Q_reg[8]) );
  DFFASRX1 \Q_reg_reg[7]  ( .D(n246), .CLK(clk), .RSTB(n188), .SETB(n187), .Q(
        Q_reg[7]) );
  DFFASRX1 \Q_reg_reg[6]  ( .D(n245), .CLK(clk), .RSTB(n186), .SETB(n185), .Q(
        Q_reg[6]) );
  DFFASRX1 \Q_reg_reg[5]  ( .D(n244), .CLK(clk), .RSTB(n184), .SETB(n183), .Q(
        Q_reg[5]) );
  DFFASRX1 \Q_reg_reg[4]  ( .D(n243), .CLK(clk), .RSTB(n182), .SETB(n181), .Q(
        Q_reg[4]) );
  DFFASRX1 \Q_reg_reg[3]  ( .D(n242), .CLK(clk), .RSTB(n180), .SETB(n179), .Q(
        Q_reg[3]) );
  DFFASRX1 \Q_reg_reg[2]  ( .D(n241), .CLK(clk), .RSTB(n178), .SETB(n177), .Q(
        Q_reg[2]) );
  DFFASRX1 \Q_reg_reg[1]  ( .D(n240), .CLK(clk), .RSTB(n176), .SETB(n175), .Q(
        Q_reg[1]) );
  AO22X1 U4 ( .IN1(N47), .IN2(n372), .IN3(n368), .IN4(count[5]), .Q(n309) );
  AO22X1 U5 ( .IN1(N46), .IN2(n372), .IN3(n368), .IN4(count[4]), .Q(n305) );
  AO22X1 U9 ( .IN1(N45), .IN2(n372), .IN3(n368), .IN4(count[3]), .Q(n306) );
  AO22X1 U13 ( .IN1(n372), .IN2(Q_reg[10]), .IN3(n368), .IN4(Q_reg[9]), .Q(
        n248) );
  OR2X1 U15 ( .IN1(n385), .IN2(Q[9]), .Q(n192) );
  AO22X1 U16 ( .IN1(n378), .IN2(Q_reg[9]), .IN3(n368), .IN4(Q_reg[8]), .Q(n247) );
  OR2X1 U19 ( .IN1(n385), .IN2(Q[8]), .Q(n190) );
  AO22X1 U20 ( .IN1(n378), .IN2(Q_reg[8]), .IN3(n368), .IN4(Q_reg[7]), .Q(n246) );
  OR2X1 U23 ( .IN1(n385), .IN2(Q[7]), .Q(n188) );
  AO22X1 U24 ( .IN1(n378), .IN2(Q_reg[7]), .IN3(n368), .IN4(Q_reg[6]), .Q(n245) );
  OR2X1 U27 ( .IN1(n385), .IN2(Q[6]), .Q(n186) );
  AO22X1 U28 ( .IN1(n377), .IN2(Q_reg[6]), .IN3(n368), .IN4(Q_reg[5]), .Q(n244) );
  OR2X1 U31 ( .IN1(n385), .IN2(Q[5]), .Q(n184) );
  AO22X1 U32 ( .IN1(n377), .IN2(Q_reg[5]), .IN3(n368), .IN4(Q_reg[4]), .Q(n243) );
  OR2X1 U35 ( .IN1(n384), .IN2(Q[4]), .Q(n182) );
  AO22X1 U36 ( .IN1(n377), .IN2(Q_reg[4]), .IN3(n368), .IN4(Q_reg[3]), .Q(n242) );
  OR2X1 U39 ( .IN1(n384), .IN2(Q[3]), .Q(n180) );
  OR2X1 U43 ( .IN1(n384), .IN2(Q[31]), .Q(n236) );
  AO22X1 U44 ( .IN1(n377), .IN2(Q_reg[31]), .IN3(n368), .IN4(Q_reg[30]), .Q(
        n269) );
  OR2X1 U47 ( .IN1(n385), .IN2(Q[30]), .Q(n234) );
  AO22X1 U48 ( .IN1(n377), .IN2(Q_reg[3]), .IN3(n368), .IN4(Q_reg[2]), .Q(n241) );
  OR2X1 U51 ( .IN1(n385), .IN2(Q[2]), .Q(n178) );
  AO22X1 U52 ( .IN1(n376), .IN2(Q_reg[30]), .IN3(n368), .IN4(Q_reg[29]), .Q(
        n268) );
  OR2X1 U55 ( .IN1(n385), .IN2(Q[29]), .Q(n232) );
  AO22X1 U56 ( .IN1(n376), .IN2(Q_reg[29]), .IN3(n368), .IN4(Q_reg[28]), .Q(
        n267) );
  OR2X1 U59 ( .IN1(n385), .IN2(Q[28]), .Q(n230) );
  AO22X1 U60 ( .IN1(n376), .IN2(Q_reg[28]), .IN3(n368), .IN4(Q_reg[27]), .Q(
        n266) );
  OR2X1 U63 ( .IN1(n385), .IN2(Q[27]), .Q(n228) );
  AO22X1 U64 ( .IN1(n376), .IN2(Q_reg[27]), .IN3(n367), .IN4(Q_reg[26]), .Q(
        n265) );
  OR2X1 U67 ( .IN1(n385), .IN2(Q[26]), .Q(n226) );
  AO22X1 U68 ( .IN1(n376), .IN2(Q_reg[26]), .IN3(n367), .IN4(Q_reg[25]), .Q(
        n264) );
  OR2X1 U71 ( .IN1(n385), .IN2(Q[25]), .Q(n224) );
  AO22X1 U72 ( .IN1(n375), .IN2(Q_reg[25]), .IN3(n367), .IN4(Q_reg[24]), .Q(
        n263) );
  OR2X1 U75 ( .IN1(n385), .IN2(Q[24]), .Q(n222) );
  AO22X1 U76 ( .IN1(n375), .IN2(Q_reg[24]), .IN3(n367), .IN4(Q_reg[23]), .Q(
        n262) );
  OR2X1 U79 ( .IN1(n385), .IN2(Q[23]), .Q(n220) );
  AO22X1 U80 ( .IN1(n375), .IN2(Q_reg[23]), .IN3(n367), .IN4(Q_reg[22]), .Q(
        n261) );
  OR2X1 U83 ( .IN1(n385), .IN2(Q[22]), .Q(n218) );
  AO22X1 U84 ( .IN1(n375), .IN2(Q_reg[22]), .IN3(n367), .IN4(Q_reg[21]), .Q(
        n260) );
  OR2X1 U87 ( .IN1(n385), .IN2(Q[21]), .Q(n216) );
  AO22X1 U88 ( .IN1(n374), .IN2(Q_reg[21]), .IN3(n367), .IN4(Q_reg[20]), .Q(
        n259) );
  OR2X1 U91 ( .IN1(n386), .IN2(Q[20]), .Q(n214) );
  AO22X1 U92 ( .IN1(n374), .IN2(Q_reg[2]), .IN3(n367), .IN4(Q_reg[1]), .Q(n240) );
  OR2X1 U95 ( .IN1(n386), .IN2(Q[1]), .Q(n176) );
  AO22X1 U96 ( .IN1(n374), .IN2(Q_reg[20]), .IN3(n367), .IN4(Q_reg[19]), .Q(
        n258) );
  OR2X1 U99 ( .IN1(n386), .IN2(Q[19]), .Q(n212) );
  AO22X1 U100 ( .IN1(n374), .IN2(Q_reg[19]), .IN3(n367), .IN4(Q_reg[18]), .Q(
        n257) );
  OR2X1 U103 ( .IN1(n386), .IN2(Q[18]), .Q(n210) );
  AO22X1 U104 ( .IN1(n374), .IN2(Q_reg[18]), .IN3(n367), .IN4(Q_reg[17]), .Q(
        n256) );
  OR2X1 U107 ( .IN1(n386), .IN2(Q[17]), .Q(n208) );
  AO22X1 U108 ( .IN1(n373), .IN2(Q_reg[17]), .IN3(n367), .IN4(Q_reg[16]), .Q(
        n255) );
  OR2X1 U111 ( .IN1(n386), .IN2(Q[16]), .Q(n206) );
  AO22X1 U112 ( .IN1(n373), .IN2(Q_reg[16]), .IN3(n367), .IN4(Q_reg[15]), .Q(
        n254) );
  OR2X1 U115 ( .IN1(n385), .IN2(Q[15]), .Q(n204) );
  AO22X1 U116 ( .IN1(n373), .IN2(Q_reg[15]), .IN3(n367), .IN4(Q_reg[14]), .Q(
        n253) );
  OR2X1 U119 ( .IN1(n386), .IN2(Q[14]), .Q(n202) );
  AO22X1 U120 ( .IN1(n373), .IN2(Q_reg[14]), .IN3(n367), .IN4(Q_reg[13]), .Q(
        n252) );
  OR2X1 U123 ( .IN1(n386), .IN2(Q[13]), .Q(n200) );
  AO22X1 U124 ( .IN1(n373), .IN2(Q_reg[13]), .IN3(n367), .IN4(Q_reg[12]), .Q(
        n251) );
  OR2X1 U127 ( .IN1(n386), .IN2(Q[12]), .Q(n198) );
  AO22X1 U128 ( .IN1(n372), .IN2(Q_reg[12]), .IN3(n367), .IN4(Q_reg[11]), .Q(
        n250) );
  OR2X1 U131 ( .IN1(n386), .IN2(Q[11]), .Q(n196) );
  AO22X1 U132 ( .IN1(n375), .IN2(Q_reg[11]), .IN3(n367), .IN4(Q_reg[10]), .Q(
        n249) );
  OR2X1 U136 ( .IN1(n386), .IN2(Q[10]), .Q(n194) );
  OR2X1 U140 ( .IN1(n386), .IN2(Q[0]), .Q(n238) );
  BoothMultiplier_DW01_sub_1 sub_61 ( .A({Acc[31:17], n328, Acc[15:11], n320, 
        Acc[9:6], n334, Acc[4:3], n326, Acc[1:0]}), .B(M_reg), .CI(1'b0), 
        .DIFF(case_sub) );
  BoothMultiplier_DW01_add_1 add_57 ( .A({Acc[31:25], n402, Acc[23:22], n406, 
        Acc[20:18], n411, Acc[16], n337, n415, n336, n338, Acc[11:10], n339, 
        n318, n340, n335, n323, n342, n343, n341, n344, n327}), .B(M_reg), 
        .CI(1'b0), .SUM(case_add) );
  LATCHX1 \M_reg_reg[2]  ( .CLK(n381), .D(M[2]), .Q(M_reg[2]) );
  LATCHX1 \M_reg_reg[9]  ( .CLK(n381), .D(M[9]), .Q(M_reg[9]) );
  LATCHX1 \M_reg_reg[7]  ( .CLK(n381), .D(M[7]), .Q(M_reg[7]) );
  LATCHX1 \M_reg_reg[4]  ( .CLK(n381), .D(M[4]), .Q(M_reg[4]) );
  NBUFFX4 U246 ( .INP(n320), .Z(n322) );
  INVX0 U247 ( .INP(n433), .ZN(n394) );
  OR2X1 U248 ( .IN1(n329), .IN2(n331), .Q(n302) );
  DELLN1X2 U249 ( .INP(n318), .Z(n321) );
  NBUFFX2 U250 ( .INP(Acc[9]), .Z(n319) );
  NBUFFX2 U251 ( .INP(n343), .Z(n324) );
  NBUFFX2 U252 ( .INP(Acc[1]), .Z(n325) );
  INVX0 U253 ( .INP(n151), .ZN(n317) );
  INVX0 U254 ( .INP(n148), .ZN(n318) );
  INVX0 U255 ( .INP(n150), .ZN(n320) );
  INVX0 U256 ( .INP(n145), .ZN(n323) );
  INVX0 U257 ( .INP(n142), .ZN(n326) );
  INVX0 U258 ( .INP(n140), .ZN(n327) );
  INVX0 U259 ( .INP(n156), .ZN(n328) );
  AO22X1 U260 ( .IN1(case_sub[64]), .IN2(n350), .IN3(case_add[64]), .IN4(n351), 
        .Q(n329) );
  INVX0 U261 ( .INP(n371), .ZN(n367) );
  INVX0 U262 ( .INP(n371), .ZN(n368) );
  INVX0 U263 ( .INP(n371), .ZN(n369) );
  NBUFFX2 U264 ( .INP(n330), .Z(n347) );
  NBUFFX2 U265 ( .INP(n333), .Z(n350) );
  NBUFFX2 U266 ( .INP(N4), .Z(n371) );
  NBUFFX2 U267 ( .INP(n332), .Z(n353) );
  NBUFFX2 U268 ( .INP(N4), .Z(n370) );
  NBUFFX2 U269 ( .INP(N4), .Z(n372) );
  NBUFFX2 U270 ( .INP(N4), .Z(n373) );
  NBUFFX2 U271 ( .INP(N4), .Z(n374) );
  NBUFFX2 U272 ( .INP(N4), .Z(n375) );
  NBUFFX2 U273 ( .INP(N4), .Z(n376) );
  NBUFFX2 U274 ( .INP(N4), .Z(n377) );
  NBUFFX2 U275 ( .INP(N4), .Z(n378) );
  AND2X1 U276 ( .IN1(n394), .IN2(n370), .Q(n330) );
  INVX0 U277 ( .INP(n437), .ZN(n441) );
  INVX0 U278 ( .INP(n435), .ZN(n439) );
  INVX0 U279 ( .INP(n436), .ZN(n440) );
  NBUFFX2 U280 ( .INP(n442), .Z(n354) );
  NBUFFX2 U281 ( .INP(n442), .Z(n355) );
  NBUFFX2 U282 ( .INP(n442), .Z(n356) );
  NBUFFX2 U283 ( .INP(n442), .Z(n357) );
  NBUFFX2 U284 ( .INP(n442), .Z(n358) );
  NBUFFX2 U285 ( .INP(n442), .Z(n359) );
  NBUFFX2 U286 ( .INP(n442), .Z(n360) );
  NBUFFX2 U287 ( .INP(n442), .Z(n361) );
  NBUFFX2 U288 ( .INP(n442), .Z(n362) );
  NBUFFX2 U289 ( .INP(n442), .Z(n363) );
  NBUFFX2 U290 ( .INP(n442), .Z(n364) );
  NBUFFX2 U291 ( .INP(n442), .Z(n365) );
  NBUFFX2 U292 ( .INP(n442), .Z(n366) );
  AOI21X1 U293 ( .IN1(n433), .IN2(n370), .IN3(n171), .QN(n331) );
  NOR2X0 U294 ( .IN1(count[0]), .IN2(n367), .QN(n310) );
  AND3X1 U295 ( .IN1(n172), .IN2(n173), .IN3(n370), .Q(n332) );
  AND3X1 U296 ( .IN1(n370), .IN2(n312), .IN3(n316), .Q(n333) );
  NOR3X0 U297 ( .IN1(count[2]), .IN2(count[3]), .IN3(count[4]), .QN(n393) );
  INVX0 U298 ( .INP(n144), .ZN(n427) );
  INVX0 U299 ( .INP(n146), .ZN(n424) );
  INVX0 U300 ( .INP(n154), .ZN(n415) );
  INVX0 U301 ( .INP(n157), .ZN(n411) );
  INVX0 U302 ( .INP(n161), .ZN(n406) );
  INVX0 U303 ( .INP(n164), .ZN(n402) );
  INVX0 U304 ( .INP(n168), .ZN(n397) );
  NBUFFX2 U305 ( .INP(oClk), .Z(n391) );
  NBUFFX2 U306 ( .INP(oClk), .Z(n390) );
  NBUFFX2 U307 ( .INP(oClk), .Z(n389) );
  NBUFFX2 U308 ( .INP(oClk), .Z(n388) );
  NBUFFX2 U309 ( .INP(oClk), .Z(n387) );
  INVX0 U310 ( .INP(oRst), .ZN(n442) );
  NBUFFX2 U311 ( .INP(oClk), .Z(n392) );
  NBUFFX2 U312 ( .INP(rst), .Z(n381) );
  NBUFFX2 U313 ( .INP(rst), .Z(n380) );
  NBUFFX2 U314 ( .INP(rst), .Z(n379) );
  NBUFFX2 U315 ( .INP(rst), .Z(n382) );
  NAND2X1 U316 ( .IN1(Q[10]), .IN2(n381), .QN(n193) );
  NAND2X1 U317 ( .IN1(Q[11]), .IN2(n381), .QN(n195) );
  NAND2X1 U318 ( .IN1(Q[12]), .IN2(n381), .QN(n197) );
  NAND2X1 U319 ( .IN1(Q[13]), .IN2(n381), .QN(n199) );
  NAND2X1 U320 ( .IN1(Q[14]), .IN2(n381), .QN(n201) );
  NAND2X1 U321 ( .IN1(Q[15]), .IN2(n381), .QN(n203) );
  NAND2X1 U322 ( .IN1(Q[16]), .IN2(n381), .QN(n205) );
  NAND2X1 U323 ( .IN1(Q[0]), .IN2(n381), .QN(n237) );
  NAND2X1 U324 ( .IN1(Q[1]), .IN2(n380), .QN(n175) );
  NAND2X1 U325 ( .IN1(Q[2]), .IN2(n379), .QN(n177) );
  NAND2X1 U326 ( .IN1(Q[3]), .IN2(n379), .QN(n179) );
  NAND2X1 U327 ( .IN1(Q[4]), .IN2(n379), .QN(n181) );
  NAND2X1 U328 ( .IN1(Q[5]), .IN2(n379), .QN(n183) );
  NAND2X1 U329 ( .IN1(Q[6]), .IN2(n379), .QN(n185) );
  NAND2X1 U330 ( .IN1(Q[7]), .IN2(n379), .QN(n187) );
  NAND2X1 U331 ( .IN1(Q[8]), .IN2(n379), .QN(n189) );
  NAND2X1 U332 ( .IN1(Q[9]), .IN2(n379), .QN(n191) );
  NAND2X1 U333 ( .IN1(Q[17]), .IN2(n380), .QN(n207) );
  NAND2X1 U334 ( .IN1(Q[18]), .IN2(n380), .QN(n209) );
  NAND2X1 U335 ( .IN1(Q[19]), .IN2(n380), .QN(n211) );
  NAND2X1 U336 ( .IN1(Q[20]), .IN2(n380), .QN(n213) );
  NAND2X1 U337 ( .IN1(Q[21]), .IN2(n380), .QN(n215) );
  NAND2X1 U338 ( .IN1(Q[22]), .IN2(n380), .QN(n217) );
  NAND2X1 U339 ( .IN1(Q[23]), .IN2(n380), .QN(n219) );
  NAND2X1 U340 ( .IN1(Q[24]), .IN2(n380), .QN(n221) );
  NAND2X1 U341 ( .IN1(Q[25]), .IN2(n380), .QN(n223) );
  NAND2X1 U342 ( .IN1(Q[26]), .IN2(n380), .QN(n225) );
  NAND2X1 U343 ( .IN1(Q[27]), .IN2(n380), .QN(n227) );
  NAND2X1 U344 ( .IN1(Q[28]), .IN2(n379), .QN(n229) );
  NAND2X1 U345 ( .IN1(Q[29]), .IN2(n379), .QN(n231) );
  NAND2X1 U346 ( .IN1(Q[30]), .IN2(n379), .QN(n233) );
  NAND2X1 U347 ( .IN1(Q[31]), .IN2(n379), .QN(n235) );
  INVX0 U348 ( .INP(n145), .ZN(n334) );
  INVX0 U349 ( .INP(n146), .ZN(n335) );
  INVX0 U350 ( .INP(n153), .ZN(n336) );
  INVX0 U351 ( .INP(n155), .ZN(n337) );
  INVX0 U352 ( .INP(n152), .ZN(n338) );
  INVX0 U353 ( .INP(n149), .ZN(n339) );
  INVX0 U354 ( .INP(n147), .ZN(n340) );
  INVX0 U355 ( .INP(n142), .ZN(n341) );
  INVX0 U356 ( .INP(n144), .ZN(n342) );
  INVX0 U357 ( .INP(n143), .ZN(n343) );
  INVX0 U358 ( .INP(n141), .ZN(n344) );
  NBUFFX2 U359 ( .INP(n330), .Z(n345) );
  NBUFFX2 U360 ( .INP(n330), .Z(n346) );
  NBUFFX2 U361 ( .INP(n333), .Z(n348) );
  NBUFFX2 U362 ( .INP(n333), .Z(n349) );
  NBUFFX2 U363 ( .INP(n332), .Z(n351) );
  NBUFFX2 U364 ( .INP(n332), .Z(n352) );
  INVX0 U365 ( .INP(n381), .ZN(n383) );
  INVX0 U366 ( .INP(n381), .ZN(n384) );
  INVX0 U367 ( .INP(n381), .ZN(n385) );
  INVX0 U368 ( .INP(n381), .ZN(n386) );
  NAND4X0 U369 ( .IN1(n314), .IN2(n313), .IN3(n315), .IN4(n393), .QN(N4) );
  AND2X1 U370 ( .IN1(N44), .IN2(n371), .Q(n307) );
  AND2X1 U371 ( .IN1(N43), .IN2(n371), .Q(n308) );
  MUX21X1 U372 ( .IN1(Q_reg[1]), .IN2(n312), .S(n367), .Q(n304) );
  MUX21X1 U373 ( .IN1(n312), .IN2(n172), .S(n367), .Q(n303) );
  XOR2X1 U374 ( .IN1(n312), .IN2(n172), .Q(n433) );
  AO22X1 U375 ( .IN1(n350), .IN2(case_sub[64]), .IN3(n351), .IN4(case_add[64]), 
        .Q(n432) );
  AO221X1 U376 ( .IN1(n345), .IN2(Acc[31]), .IN3(n367), .IN4(Acc[30]), .IN5(
        n432), .Q(n301) );
  AO22X1 U377 ( .IN1(n368), .IN2(Acc[29]), .IN3(n345), .IN4(Acc[30]), .Q(n395)
         );
  AO221X1 U378 ( .IN1(n351), .IN2(case_add[63]), .IN3(case_sub[63]), .IN4(n350), .IN5(n395), .Q(n300) );
  AO22X1 U379 ( .IN1(n369), .IN2(n397), .IN3(n345), .IN4(Acc[29]), .Q(n396) );
  AO221X1 U380 ( .IN1(n351), .IN2(case_add[62]), .IN3(case_sub[62]), .IN4(n350), .IN5(n396), .Q(n299) );
  AO22X1 U381 ( .IN1(n369), .IN2(Acc[27]), .IN3(n345), .IN4(n397), .Q(n398) );
  AO221X1 U382 ( .IN1(n351), .IN2(case_add[61]), .IN3(case_sub[61]), .IN4(n350), .IN5(n398), .Q(n298) );
  AO22X1 U383 ( .IN1(n369), .IN2(Acc[26]), .IN3(n345), .IN4(Acc[27]), .Q(n399)
         );
  AO221X1 U384 ( .IN1(case_add[60]), .IN2(n351), .IN3(case_sub[60]), .IN4(n350), .IN5(n399), .Q(n297) );
  AO22X1 U385 ( .IN1(n369), .IN2(Acc[25]), .IN3(n345), .IN4(Acc[26]), .Q(n400)
         );
  AO221X1 U386 ( .IN1(case_add[59]), .IN2(n351), .IN3(case_sub[59]), .IN4(n350), .IN5(n400), .Q(n296) );
  AO22X1 U387 ( .IN1(n369), .IN2(n402), .IN3(n345), .IN4(Acc[25]), .Q(n401) );
  AO221X1 U388 ( .IN1(case_add[58]), .IN2(n351), .IN3(case_sub[58]), .IN4(n350), .IN5(n401), .Q(n295) );
  AO22X1 U389 ( .IN1(n369), .IN2(Acc[23]), .IN3(n345), .IN4(n402), .Q(n403) );
  AO221X1 U390 ( .IN1(case_add[57]), .IN2(n351), .IN3(case_sub[57]), .IN4(n350), .IN5(n403), .Q(n294) );
  AO22X1 U391 ( .IN1(n369), .IN2(Acc[22]), .IN3(n345), .IN4(Acc[23]), .Q(n404)
         );
  AO221X1 U392 ( .IN1(case_add[56]), .IN2(n351), .IN3(case_sub[56]), .IN4(n349), .IN5(n404), .Q(n293) );
  AO22X1 U393 ( .IN1(n369), .IN2(n406), .IN3(n345), .IN4(Acc[22]), .Q(n405) );
  AO221X1 U394 ( .IN1(case_add[55]), .IN2(n351), .IN3(case_sub[55]), .IN4(n349), .IN5(n405), .Q(n292) );
  AO22X1 U395 ( .IN1(n369), .IN2(Acc[20]), .IN3(n345), .IN4(n406), .Q(n407) );
  AO221X1 U396 ( .IN1(case_add[54]), .IN2(n351), .IN3(case_sub[54]), .IN4(n349), .IN5(n407), .Q(n291) );
  AO22X1 U397 ( .IN1(n369), .IN2(Acc[19]), .IN3(n345), .IN4(Acc[20]), .Q(n408)
         );
  AO221X1 U398 ( .IN1(case_add[53]), .IN2(n351), .IN3(case_sub[53]), .IN4(n349), .IN5(n408), .Q(n290) );
  AO22X1 U399 ( .IN1(n369), .IN2(Acc[18]), .IN3(n345), .IN4(Acc[19]), .Q(n409)
         );
  AO221X1 U400 ( .IN1(case_add[52]), .IN2(n351), .IN3(case_sub[52]), .IN4(n349), .IN5(n409), .Q(n289) );
  AO22X1 U401 ( .IN1(n368), .IN2(n411), .IN3(n346), .IN4(Acc[18]), .Q(n410) );
  AO221X1 U402 ( .IN1(case_add[51]), .IN2(n352), .IN3(case_sub[51]), .IN4(n349), .IN5(n410), .Q(n288) );
  AO22X1 U403 ( .IN1(n369), .IN2(Acc[16]), .IN3(n346), .IN4(n411), .Q(n412) );
  AO221X1 U404 ( .IN1(case_add[50]), .IN2(n352), .IN3(case_sub[50]), .IN4(n349), .IN5(n412), .Q(n287) );
  AO22X1 U405 ( .IN1(n369), .IN2(Acc[15]), .IN3(n346), .IN4(Acc[16]), .Q(n413)
         );
  AO221X1 U406 ( .IN1(case_add[49]), .IN2(n352), .IN3(case_sub[49]), .IN4(n349), .IN5(n413), .Q(n286) );
  AO22X1 U407 ( .IN1(n369), .IN2(n415), .IN3(n346), .IN4(Acc[15]), .Q(n414) );
  AO221X1 U408 ( .IN1(case_add[48]), .IN2(n352), .IN3(case_sub[48]), .IN4(n349), .IN5(n414), .Q(n285) );
  AO22X1 U409 ( .IN1(n369), .IN2(Acc[13]), .IN3(n346), .IN4(n415), .Q(n416) );
  AO221X1 U410 ( .IN1(case_add[47]), .IN2(n352), .IN3(case_sub[47]), .IN4(n349), .IN5(n416), .Q(n284) );
  AO22X1 U411 ( .IN1(n369), .IN2(Acc[12]), .IN3(n346), .IN4(Acc[13]), .Q(n417)
         );
  AO221X1 U412 ( .IN1(case_add[46]), .IN2(n352), .IN3(case_sub[46]), .IN4(n349), .IN5(n417), .Q(n283) );
  AO22X1 U413 ( .IN1(n369), .IN2(n317), .IN3(n346), .IN4(Acc[12]), .Q(n418) );
  AO221X1 U414 ( .IN1(case_add[45]), .IN2(n352), .IN3(case_sub[45]), .IN4(n349), .IN5(n418), .Q(n282) );
  AO22X1 U415 ( .IN1(n369), .IN2(n322), .IN3(n346), .IN4(n317), .Q(n419) );
  AO221X1 U416 ( .IN1(case_add[44]), .IN2(n352), .IN3(case_sub[44]), .IN4(n348), .IN5(n419), .Q(n281) );
  AO22X1 U417 ( .IN1(n369), .IN2(n319), .IN3(n346), .IN4(n322), .Q(n420) );
  AO221X1 U418 ( .IN1(case_add[43]), .IN2(n352), .IN3(case_sub[43]), .IN4(n348), .IN5(n420), .Q(n280) );
  AO22X1 U419 ( .IN1(n369), .IN2(n321), .IN3(n346), .IN4(n319), .Q(n421) );
  AO221X1 U420 ( .IN1(case_add[42]), .IN2(n352), .IN3(case_sub[42]), .IN4(n348), .IN5(n421), .Q(n279) );
  AO22X1 U421 ( .IN1(n369), .IN2(Acc[7]), .IN3(n346), .IN4(n321), .Q(n422) );
  AO221X1 U422 ( .IN1(case_add[41]), .IN2(n352), .IN3(case_sub[41]), .IN4(n348), .IN5(n422), .Q(n278) );
  AO22X1 U423 ( .IN1(n368), .IN2(n424), .IN3(n346), .IN4(Acc[7]), .Q(n423) );
  AO221X1 U424 ( .IN1(case_add[40]), .IN2(n352), .IN3(case_sub[40]), .IN4(n348), .IN5(n423), .Q(n277) );
  AO22X1 U425 ( .IN1(n368), .IN2(Acc[5]), .IN3(n346), .IN4(n424), .Q(n425) );
  AO221X1 U426 ( .IN1(case_add[39]), .IN2(n352), .IN3(case_sub[39]), .IN4(n348), .IN5(n425), .Q(n276) );
  AO22X1 U427 ( .IN1(n368), .IN2(n427), .IN3(n347), .IN4(Acc[5]), .Q(n426) );
  AO221X1 U428 ( .IN1(case_add[38]), .IN2(n353), .IN3(case_sub[38]), .IN4(n348), .IN5(n426), .Q(n275) );
  AO22X1 U429 ( .IN1(n368), .IN2(n324), .IN3(n347), .IN4(n427), .Q(n428) );
  AO221X1 U430 ( .IN1(case_add[37]), .IN2(n353), .IN3(case_sub[37]), .IN4(n348), .IN5(n428), .Q(n274) );
  AO22X1 U431 ( .IN1(n368), .IN2(Acc[2]), .IN3(n347), .IN4(n324), .Q(n429) );
  AO221X1 U432 ( .IN1(case_add[36]), .IN2(n353), .IN3(case_sub[36]), .IN4(n348), .IN5(n429), .Q(n273) );
  AO22X1 U433 ( .IN1(n368), .IN2(n325), .IN3(n347), .IN4(Acc[2]), .Q(n430) );
  AO221X1 U434 ( .IN1(case_add[35]), .IN2(n353), .IN3(case_sub[35]), .IN4(n348), .IN5(n430), .Q(n272) );
  AO22X1 U435 ( .IN1(n368), .IN2(n327), .IN3(n347), .IN4(n325), .Q(n431) );
  AO221X1 U436 ( .IN1(case_add[34]), .IN2(n353), .IN3(case_sub[34]), .IN4(n348), .IN5(n431), .Q(n271) );
  AO22X1 U437 ( .IN1(n368), .IN2(Q_reg[31]), .IN3(n347), .IN4(n327), .Q(n434)
         );
  AO221X1 U438 ( .IN1(case_add[33]), .IN2(n353), .IN3(case_sub[33]), .IN4(n348), .IN5(n434), .Q(n270) );
  NOR2X0 U439 ( .IN1(count[1]), .IN2(count[0]), .QN(n435) );
  AO21X1 U440 ( .IN1(count[1]), .IN2(count[0]), .IN3(n435), .Q(N43) );
  NOR2X0 U441 ( .IN1(n439), .IN2(count[2]), .QN(n436) );
  AO21X1 U442 ( .IN1(count[2]), .IN2(n439), .IN3(n436), .Q(N44) );
  NOR2X0 U443 ( .IN1(n440), .IN2(count[3]), .QN(n437) );
  AO21X1 U444 ( .IN1(count[3]), .IN2(n440), .IN3(n437), .Q(N45) );
  XNOR2X1 U445 ( .IN1(count[4]), .IN2(n441), .Q(N46) );
  NOR2X0 U446 ( .IN1(count[4]), .IN2(n441), .QN(n438) );
  XOR2X1 U447 ( .IN1(count[5]), .IN2(n438), .Q(N47) );
endmodule

