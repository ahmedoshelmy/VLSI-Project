
module BoothMultiplier_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372;

  NAND4X0 U3 ( .IN1(n262), .IN2(n260), .IN3(n261), .IN4(n259), .QN(n55) );
  INVX0 U4 ( .INP(B[31]), .ZN(n31) );
  NAND2X1 U5 ( .IN1(B[10]), .IN2(n318), .QN(n317) );
  OR2X1 U6 ( .IN1(n26), .IN2(n204), .Q(n25) );
  OR2X1 U7 ( .IN1(n22), .IN2(n182), .Q(n21) );
  AND2X1 U8 ( .IN1(n175), .IN2(n176), .Q(n3) );
  XOR3X1 U9 ( .IN1(n149), .IN2(B[29]), .IN3(n57), .Q(DIFF[29]) );
  AND2X1 U10 ( .IN1(n206), .IN2(n207), .Q(n1) );
  AND2X1 U11 ( .IN1(n272), .IN2(n305), .Q(n2) );
  AND2X1 U12 ( .IN1(n169), .IN2(n170), .Q(n4) );
  AND2X1 U13 ( .IN1(n186), .IN2(n187), .Q(n5) );
  AND2X1 U14 ( .IN1(n54), .IN2(n204), .Q(n6) );
  NAND2X1 U15 ( .IN1(n20), .IN2(n21), .QN(n7) );
  NAND2X1 U16 ( .IN1(n306), .IN2(n11), .QN(n8) );
  AND2X1 U17 ( .IN1(n8), .IN2(n9), .Q(n301) );
  OR2X1 U18 ( .IN1(n10), .IN2(n272), .Q(n9) );
  INVX0 U19 ( .INP(n274), .ZN(n10) );
  AND2X1 U20 ( .IN1(n295), .IN2(n274), .Q(n11) );
  NAND2X1 U21 ( .IN1(n159), .IN2(n15), .QN(n12) );
  AND2X1 U22 ( .IN1(n12), .IN2(n13), .Q(n144) );
  OR2X1 U23 ( .IN1(n14), .IN2(n148), .Q(n13) );
  INVX0 U24 ( .INP(n147), .ZN(n14) );
  AND2X1 U25 ( .IN1(n158), .IN2(n147), .Q(n15) );
  XOR3X1 U26 ( .IN1(n145), .IN2(B[30]), .IN3(n144), .Q(DIFF[30]) );
  NAND2X0 U27 ( .IN1(A[27]), .IN2(n168), .QN(n164) );
  NAND2X0 U28 ( .IN1(n170), .IN2(n19), .QN(n16) );
  AND2X1 U29 ( .IN1(n16), .IN2(n17), .Q(n161) );
  OR2X1 U30 ( .IN1(n18), .IN2(n165), .Q(n17) );
  INVX0 U31 ( .INP(n164), .ZN(n18) );
  AND2X1 U32 ( .IN1(n169), .IN2(n164), .Q(n19) );
  NAND2X0 U33 ( .IN1(n181), .IN2(n182), .QN(n183) );
  NAND2X0 U34 ( .IN1(n187), .IN2(n23), .QN(n20) );
  INVX0 U35 ( .INP(n181), .ZN(n22) );
  AND2X1 U36 ( .IN1(n186), .IN2(n181), .Q(n23) );
  NAND2X0 U37 ( .IN1(n55), .IN2(n27), .QN(n24) );
  AND2X1 U38 ( .IN1(n24), .IN2(n25), .Q(n201) );
  INVX0 U39 ( .INP(n202), .ZN(n26) );
  AND2X1 U40 ( .IN1(n1), .IN2(n202), .Q(n27) );
  NAND2X0 U41 ( .IN1(A[28]), .IN2(n163), .QN(n158) );
  XOR3X1 U42 ( .IN1(n162), .IN2(B[28]), .IN3(n161), .Q(DIFF[28]) );
  AND2X1 U43 ( .IN1(n61), .IN2(n44), .Q(n28) );
  NAND2X0 U44 ( .IN1(n33), .IN2(n32), .QN(n29) );
  NAND2X0 U45 ( .IN1(n29), .IN2(n30), .QN(n43) );
  AND2X1 U46 ( .IN1(n46), .IN2(n76), .Q(n30) );
  NAND2X0 U47 ( .IN1(B[25]), .IN2(n179), .QN(n177) );
  NAND2X0 U48 ( .IN1(B[24]), .IN2(n184), .QN(n182) );
  XOR3X1 U49 ( .IN1(A[31]), .IN2(n31), .IN3(n140), .Q(DIFF[31]) );
  NAND2X0 U50 ( .IN1(n175), .IN2(n177), .QN(n178) );
  NAND2X0 U51 ( .IN1(A[25]), .IN2(n180), .QN(n175) );
  NAND2X1 U52 ( .IN1(n39), .IN2(n35), .QN(n32) );
  NAND2X0 U53 ( .IN1(n32), .IN2(n33), .QN(n75) );
  OR2X1 U54 ( .IN1(n34), .IN2(n37), .Q(n33) );
  INVX0 U55 ( .INP(n72), .ZN(n34) );
  AND2X1 U56 ( .IN1(n205), .IN2(n72), .Q(n35) );
  NOR2X0 U57 ( .IN1(n88), .IN2(A[6]), .QN(n36) );
  OR2X1 U58 ( .IN1(n38), .IN2(n40), .Q(n37) );
  INVX0 U59 ( .INP(n66), .ZN(n38) );
  AND2X1 U60 ( .IN1(n42), .IN2(n66), .Q(n39) );
  OR2X1 U61 ( .IN1(n41), .IN2(n64), .Q(n40) );
  INVX0 U62 ( .INP(n62), .ZN(n41) );
  AND2X1 U63 ( .IN1(n204), .IN2(n62), .Q(n42) );
  OR2X1 U64 ( .IN1(n45), .IN2(n48), .Q(n44) );
  INVX0 U65 ( .INP(n158), .ZN(n45) );
  AND2X1 U66 ( .IN1(n50), .IN2(n158), .Q(n46) );
  NAND2X0 U67 ( .IN1(n176), .IN2(n50), .QN(n47) );
  NAND2X0 U68 ( .IN1(n47), .IN2(n48), .QN(n159) );
  OR2X1 U69 ( .IN1(n49), .IN2(n51), .Q(n48) );
  INVX0 U70 ( .INP(n79), .ZN(n49) );
  AND2X1 U71 ( .IN1(n53), .IN2(n79), .Q(n50) );
  OR2X1 U72 ( .IN1(n52), .IN2(n71), .Q(n51) );
  INVX0 U73 ( .INP(n69), .ZN(n52) );
  AND2X1 U74 ( .IN1(n175), .IN2(n69), .Q(n53) );
  NAND2X0 U75 ( .IN1(n1), .IN2(n55), .QN(n54) );
  AND2X1 U76 ( .IN1(n134), .IN2(n338), .Q(n56) );
  NAND2X0 U77 ( .IN1(n1), .IN2(n208), .QN(n205) );
  NAND2X0 U78 ( .IN1(B[20]), .IN2(n224), .QN(n207) );
  NAND2X0 U79 ( .IN1(n158), .IN2(n159), .QN(n57) );
  NAND2X0 U80 ( .IN1(n43), .IN2(n28), .QN(n58) );
  AND2X1 U81 ( .IN1(n58), .IN2(n59), .Q(n142) );
  OR2X1 U82 ( .IN1(n60), .IN2(n147), .Q(n59) );
  INVX0 U83 ( .INP(n143), .ZN(n60) );
  AND2X1 U84 ( .IN1(n148), .IN2(n143), .Q(n61) );
  OR2X1 U85 ( .IN1(n63), .IN2(n200), .Q(n62) );
  INVX0 U86 ( .INP(n68), .ZN(n63) );
  AND2X1 U87 ( .IN1(n202), .IN2(n68), .Q(n64) );
  NAND2X0 U88 ( .IN1(n175), .IN2(n176), .QN(n65) );
  OR2X1 U89 ( .IN1(n67), .IN2(n194), .Q(n66) );
  INVX0 U90 ( .INP(n74), .ZN(n67) );
  AND2X1 U91 ( .IN1(n197), .IN2(n74), .Q(n68) );
  OR2X1 U92 ( .IN1(n70), .IN2(n169), .Q(n69) );
  INVX0 U93 ( .INP(n81), .ZN(n70) );
  AND2X1 U94 ( .IN1(n171), .IN2(n81), .Q(n71) );
  OR2X1 U95 ( .IN1(n73), .IN2(n186), .Q(n72) );
  INVX0 U96 ( .INP(n78), .ZN(n73) );
  AND2X1 U97 ( .IN1(n189), .IN2(n78), .Q(n74) );
  AND2X1 U98 ( .IN1(n75), .IN2(n76), .Q(n176) );
  OR2X1 U99 ( .IN1(n77), .IN2(n181), .Q(n76) );
  INVX0 U100 ( .INP(n177), .ZN(n77) );
  AND2X1 U101 ( .IN1(n182), .IN2(n177), .Q(n78) );
  OR2X1 U102 ( .IN1(n80), .IN2(n164), .Q(n79) );
  INVX0 U103 ( .INP(n160), .ZN(n80) );
  AND2X1 U104 ( .IN1(n165), .IN2(n160), .Q(n81) );
  NAND2X0 U105 ( .IN1(n128), .IN2(n123), .QN(n357) );
  NAND2X0 U106 ( .IN1(n237), .IN2(n236), .QN(n222) );
  NAND2X0 U107 ( .IN1(n221), .IN2(n219), .QN(n209) );
  NAND2X0 U108 ( .IN1(n315), .IN2(n316), .QN(n312) );
  NAND2X0 U109 ( .IN1(n311), .IN2(n277), .QN(n306) );
  NAND2X0 U110 ( .IN1(n328), .IN2(n329), .QN(n327) );
  NAND2X0 U111 ( .IN1(n122), .IN2(n123), .QN(n121) );
  NAND2X0 U112 ( .IN1(n219), .IN2(n217), .QN(n230) );
  NAND2X0 U113 ( .IN1(n236), .IN2(n234), .QN(n241) );
  NAND2X0 U114 ( .IN1(n207), .IN2(n211), .QN(n213) );
  NAND2X0 U115 ( .IN1(n202), .IN2(n200), .QN(n203) );
  NAND2X0 U116 ( .IN1(n194), .IN2(n197), .QN(n199) );
  NAND2X0 U117 ( .IN1(B[18]), .IN2(n250), .QN(n236) );
  NAND2X0 U118 ( .IN1(B[4]), .IN2(n359), .QN(n128) );
  INVX0 U119 ( .INP(B[6]), .ZN(n88) );
  NAND2X0 U120 ( .IN1(B[8]), .IN2(n368), .QN(n109) );
  INVX0 U121 ( .INP(B[11]), .ZN(n89) );
  NAND2X0 U122 ( .IN1(B[9]), .IN2(n369), .QN(n104) );
  NAND2X0 U123 ( .IN1(B[7]), .IN2(n360), .QN(n112) );
  NAND2X0 U124 ( .IN1(B[13]), .IN2(n309), .QN(n295) );
  NAND2X0 U125 ( .IN1(B[17]), .IN2(n257), .QN(n247) );
  INVX0 U126 ( .INP(B[12]), .ZN(n87) );
  INVX0 U127 ( .INP(B[22]), .ZN(n93) );
  INVX0 U128 ( .INP(B[21]), .ZN(n92) );
  INVX0 U129 ( .INP(n129), .ZN(n131) );
  INVX0 U130 ( .INP(n290), .ZN(n276) );
  INVX0 U131 ( .INP(n209), .ZN(n206) );
  INVX0 U132 ( .INP(n291), .ZN(n337) );
  NOR2X0 U133 ( .IN1(n232), .IN2(n218), .QN(n231) );
  NOR2X0 U134 ( .IN1(n220), .IN2(n222), .QN(n232) );
  INVX0 U135 ( .INP(n330), .ZN(n332) );
  INVX0 U136 ( .INP(n306), .ZN(n307) );
  INVX0 U137 ( .INP(n116), .ZN(n118) );
  INVX0 U138 ( .INP(n103), .ZN(n102) );
  INVX0 U139 ( .INP(n122), .ZN(n125) );
  INVX0 U140 ( .INP(n108), .ZN(n107) );
  INVX0 U141 ( .INP(n312), .ZN(n314) );
  INVX0 U142 ( .INP(n156), .ZN(n225) );
  NAND2X0 U143 ( .IN1(n335), .IN2(n336), .QN(n108) );
  NOR2X0 U144 ( .IN1(n154), .IN2(n353), .QN(n350) );
  NOR2X0 U145 ( .IN1(n82), .IN2(n210), .QN(n204) );
  INVX0 U146 ( .INP(n211), .ZN(n210) );
  NAND2X0 U147 ( .IN1(n113), .IN2(n115), .QN(n364) );
  NOR2X0 U148 ( .IN1(n269), .IN2(n270), .QN(n268) );
  INVX0 U149 ( .INP(n271), .ZN(n269) );
  NOR2X0 U150 ( .IN1(n350), .IN2(n351), .QN(n341) );
  INVX0 U151 ( .INP(n135), .ZN(n343) );
  NAND2X0 U152 ( .IN1(n270), .IN2(n301), .QN(n298) );
  NAND2X0 U153 ( .IN1(n96), .IN2(n97), .QN(n82) );
  INVX0 U154 ( .INP(n222), .ZN(n221) );
  NAND2X0 U155 ( .IN1(n312), .IN2(n294), .QN(n311) );
  AND2X1 U156 ( .IN1(n219), .IN2(n207), .Q(n99) );
  INVX0 U157 ( .INP(n277), .ZN(n275) );
  NAND2X0 U158 ( .IN1(n306), .IN2(n295), .QN(n305) );
  NOR2X0 U159 ( .IN1(n255), .IN2(n220), .QN(n253) );
  NOR2X0 U160 ( .IN1(n220), .IN2(n209), .QN(n215) );
  NAND2X0 U161 ( .IN1(n110), .IN2(n334), .QN(n103) );
  NAND2X0 U162 ( .IN1(n109), .IN2(n108), .QN(n334) );
  NAND2X1 U163 ( .IN1(n126), .IN2(n127), .QN(n122) );
  NAND2X0 U164 ( .IN1(n128), .IN2(n129), .QN(n127) );
  NAND2X0 U165 ( .IN1(n114), .IN2(n115), .QN(n111) );
  NAND2X0 U166 ( .IN1(n120), .IN2(n121), .QN(n116) );
  NAND2X0 U167 ( .IN1(n154), .IN2(n155), .QN(n138) );
  NAND2X0 U168 ( .IN1(n136), .IN2(n137), .QN(n133) );
  NAND2X0 U169 ( .IN1(n330), .IN2(n325), .QN(n329) );
  NAND2X1 U170 ( .IN1(n227), .IN2(n228), .QN(n156) );
  INVX0 U171 ( .INP(n95), .ZN(n228) );
  NAND2X0 U172 ( .IN1(n105), .IN2(n333), .QN(n330) );
  NAND2X0 U173 ( .IN1(n104), .IN2(n103), .QN(n333) );
  AND2X1 U174 ( .IN1(n134), .IN2(n135), .Q(n83) );
  NAND2X0 U175 ( .IN1(n294), .IN2(n277), .QN(n313) );
  NOR2X0 U176 ( .IN1(n152), .IN2(n153), .QN(n151) );
  INVX0 U177 ( .INP(n136), .ZN(n152) );
  NAND2X0 U178 ( .IN1(n123), .IN2(n120), .QN(n124) );
  NAND2X0 U179 ( .IN1(n104), .IN2(n105), .QN(n101) );
  NAND2X1 U180 ( .IN1(n109), .IN2(n110), .QN(n106) );
  NAND2X1 U181 ( .IN1(n128), .IN2(n126), .QN(n130) );
  NAND2X0 U182 ( .IN1(n325), .IN2(n328), .QN(n331) );
  NAND2X0 U183 ( .IN1(n272), .IN2(n295), .QN(n308) );
  AND2X1 U184 ( .IN1(n278), .IN2(n320), .Q(n84) );
  NAND2X0 U185 ( .IN1(n247), .IN2(n245), .QN(n251) );
  AND2X1 U186 ( .IN1(n271), .IN2(n260), .Q(n85) );
  NAND2X1 U187 ( .IN1(n186), .IN2(n189), .QN(n191) );
  NAND2X1 U188 ( .IN1(n169), .IN2(n171), .QN(n172) );
  NAND2X1 U189 ( .IN1(n164), .IN2(n165), .QN(n166) );
  AND2X1 U190 ( .IN1(n112), .IN2(n113), .Q(n86) );
  INVX0 U191 ( .INP(B[9]), .ZN(n370) );
  INVX0 U192 ( .INP(B[5]), .ZN(n366) );
  INVX0 U193 ( .INP(B[13]), .ZN(n310) );
  INVX0 U194 ( .INP(B[14]), .ZN(n304) );
  INVX0 U195 ( .INP(B[2]), .ZN(n352) );
  INVX0 U196 ( .INP(B[7]), .ZN(n367) );
  INVX0 U197 ( .INP(B[1]), .ZN(n356) );
  INVX0 U198 ( .INP(B[17]), .ZN(n256) );
  OR2X1 U199 ( .IN1(n87), .IN2(A[12]), .Q(n294) );
  INVX0 U200 ( .INP(B[28]), .ZN(n163) );
  NAND2X1 U201 ( .IN1(A[29]), .IN2(n150), .QN(n147) );
  INVX0 U202 ( .INP(B[29]), .ZN(n150) );
  INVX0 U203 ( .INP(B[3]), .ZN(n349) );
  OR2X1 U204 ( .IN1(n88), .IN2(A[6]), .Q(n117) );
  NAND2X1 U205 ( .IN1(B[5]), .IN2(n363), .QN(n123) );
  INVX0 U206 ( .INP(B[16]), .ZN(n296) );
  NAND2X1 U207 ( .IN1(A[30]), .IN2(n146), .QN(n141) );
  INVX0 U208 ( .INP(B[30]), .ZN(n146) );
  NAND3X0 U209 ( .IN1(A[0]), .IN2(n157), .IN3(n139), .QN(n345) );
  NAND2X1 U210 ( .IN1(B[19]), .IN2(n240), .QN(n219) );
  INVX0 U211 ( .INP(A[19]), .ZN(n240) );
  INVX0 U212 ( .INP(A[18]), .ZN(n250) );
  INVX0 U213 ( .INP(A[20]), .ZN(n224) );
  OR2X1 U214 ( .IN1(n89), .IN2(A[11]), .Q(n278) );
  NAND2X0 U215 ( .IN1(A[19]), .IN2(n239), .QN(n217) );
  INVX0 U216 ( .INP(B[19]), .ZN(n239) );
  NAND2X0 U217 ( .IN1(A[18]), .IN2(n249), .QN(n234) );
  INVX0 U218 ( .INP(B[18]), .ZN(n249) );
  NOR2X0 U219 ( .IN1(n90), .IN2(n91), .QN(n284) );
  NAND2X0 U220 ( .IN1(n109), .IN2(n104), .QN(n90) );
  NAND2X0 U221 ( .IN1(n317), .IN2(n278), .QN(n91) );
  INVX0 U222 ( .INP(A[28]), .ZN(n162) );
  NAND2X0 U223 ( .IN1(A[20]), .IN2(n223), .QN(n211) );
  INVX0 U224 ( .INP(B[20]), .ZN(n223) );
  OR2X1 U225 ( .IN1(n92), .IN2(A[21]), .Q(n202) );
  OR2X1 U226 ( .IN1(n93), .IN2(A[22]), .Q(n197) );
  NAND2X1 U227 ( .IN1(B[26]), .IN2(n173), .QN(n171) );
  INVX0 U228 ( .INP(A[26]), .ZN(n173) );
  NAND2X0 U229 ( .IN1(A[21]), .IN2(n92), .QN(n200) );
  NAND2X1 U230 ( .IN1(A[23]), .IN2(n193), .QN(n186) );
  INVX0 U231 ( .INP(B[23]), .ZN(n193) );
  NAND2X0 U232 ( .IN1(A[22]), .IN2(n93), .QN(n194) );
  NAND2X1 U233 ( .IN1(A[24]), .IN2(n185), .QN(n181) );
  INVX0 U234 ( .INP(B[24]), .ZN(n185) );
  INVX0 U235 ( .INP(B[25]), .ZN(n180) );
  NAND2X1 U236 ( .IN1(A[26]), .IN2(n174), .QN(n169) );
  INVX0 U237 ( .INP(B[26]), .ZN(n174) );
  INVX0 U238 ( .INP(B[27]), .ZN(n168) );
  NAND2X0 U239 ( .IN1(A[15]), .IN2(n299), .QN(n260) );
  INVX0 U240 ( .INP(B[15]), .ZN(n299) );
  INVX0 U241 ( .INP(A[24]), .ZN(n184) );
  NAND2X1 U242 ( .IN1(B[23]), .IN2(n192), .QN(n189) );
  INVX0 U243 ( .INP(A[23]), .ZN(n192) );
  INVX0 U244 ( .INP(A[25]), .ZN(n179) );
  NAND2X1 U245 ( .IN1(B[27]), .IN2(n167), .QN(n165) );
  INVX0 U246 ( .INP(A[27]), .ZN(n167) );
  NAND2X1 U247 ( .IN1(B[28]), .IN2(n162), .QN(n160) );
  INVX0 U248 ( .INP(B[10]), .ZN(n371) );
  INVX0 U249 ( .INP(A[29]), .ZN(n149) );
  INVX0 U250 ( .INP(A[30]), .ZN(n145) );
  NAND2X0 U251 ( .IN1(A[0]), .IN2(n347), .QN(n227) );
  NAND2X1 U252 ( .IN1(B[30]), .IN2(n145), .QN(n143) );
  NAND2X1 U253 ( .IN1(B[29]), .IN2(n149), .QN(n148) );
  INVX0 U254 ( .INP(B[0]), .ZN(n347) );
  INVX0 U255 ( .INP(B[4]), .ZN(n132) );
  INVX0 U256 ( .INP(B[8]), .ZN(n326) );
  INVX0 U257 ( .INP(n188), .ZN(n190) );
  NAND2X1 U258 ( .IN1(B[15]), .IN2(n300), .QN(n271) );
  INVX0 U259 ( .INP(n238), .ZN(n237) );
  NOR2X0 U260 ( .IN1(n220), .IN2(n238), .QN(n243) );
  INVX0 U261 ( .INP(n55), .ZN(n220) );
  NAND2X0 U262 ( .IN1(n265), .IN2(n266), .QN(n264) );
  NAND2X0 U263 ( .IN1(n289), .IN2(n129), .QN(n336) );
  NOR2X0 U264 ( .IN1(n357), .IN2(n358), .QN(n289) );
  AND2X1 U265 ( .IN1(n279), .IN2(n94), .Q(n263) );
  AND2X1 U266 ( .IN1(n276), .IN2(n278), .Q(n94) );
  NAND2X0 U267 ( .IN1(n156), .IN2(n157), .QN(n155) );
  NAND2X0 U268 ( .IN1(n154), .IN2(n157), .QN(n226) );
  NAND2X0 U269 ( .IN1(B[1]), .IN2(n348), .QN(n157) );
  OR2X1 U270 ( .IN1(n347), .IN2(A[0]), .Q(n229) );
  NOR2X0 U271 ( .IN1(n340), .IN2(n136), .QN(n351) );
  NAND2X0 U272 ( .IN1(n116), .IN2(n117), .QN(n114) );
  NAND2X0 U273 ( .IN1(n115), .IN2(n117), .QN(n119) );
  NAND2X0 U274 ( .IN1(n112), .IN2(n117), .QN(n358) );
  INVX0 U275 ( .INP(A[16]), .ZN(n297) );
  NAND2X0 U276 ( .IN1(A[16]), .IN2(n296), .QN(n254) );
  NAND2X0 U277 ( .IN1(n279), .IN2(n278), .QN(n315) );
  NAND2X0 U278 ( .IN1(n138), .IN2(n139), .QN(n137) );
  INVX0 U279 ( .INP(n139), .ZN(n153) );
  NAND2X1 U280 ( .IN1(B[2]), .IN2(n355), .QN(n139) );
  NAND2X0 U281 ( .IN1(B[0]), .IN2(n372), .QN(n95) );
  INVX0 U282 ( .INP(A[1]), .ZN(n348) );
  NAND2X0 U283 ( .IN1(n218), .IN2(n99), .QN(n96) );
  OR2X1 U284 ( .IN1(n98), .IN2(n217), .Q(n97) );
  INVX0 U285 ( .INP(n207), .ZN(n98) );
  NAND2X0 U286 ( .IN1(n337), .IN2(n288), .QN(n129) );
  NAND2X0 U287 ( .IN1(A[5]), .IN2(n366), .QN(n120) );
  INVX0 U288 ( .INP(A[5]), .ZN(n363) );
  NAND2X0 U289 ( .IN1(n248), .IN2(n254), .QN(n258) );
  INVX0 U290 ( .INP(n248), .ZN(n255) );
  NAND2X0 U291 ( .IN1(n248), .IN2(n247), .QN(n238) );
  NAND2X1 U292 ( .IN1(B[16]), .IN2(n297), .QN(n248) );
  NAND2X0 U293 ( .IN1(n361), .IN2(n362), .QN(n100) );
  NAND2X0 U294 ( .IN1(n134), .IN2(n338), .QN(n288) );
  NOR2X0 U295 ( .IN1(n339), .IN2(n153), .QN(n338) );
  INVX0 U296 ( .INP(A[4]), .ZN(n359) );
  NAND2X0 U297 ( .IN1(A[4]), .IN2(n132), .QN(n126) );
  NAND2X0 U298 ( .IN1(n100), .IN2(n112), .QN(n335) );
  NAND2X0 U299 ( .IN1(n361), .IN2(n362), .QN(n285) );
  NAND2X0 U300 ( .IN1(n139), .IN2(n134), .QN(n353) );
  INVX0 U301 ( .INP(n134), .ZN(n340) );
  NAND2X0 U302 ( .IN1(n134), .IN2(n347), .QN(n346) );
  NAND2X1 U303 ( .IN1(B[3]), .IN2(n354), .QN(n134) );
  NAND2X0 U304 ( .IN1(n244), .IN2(n245), .QN(n235) );
  NAND2X0 U305 ( .IN1(A[9]), .IN2(n370), .QN(n105) );
  INVX0 U306 ( .INP(A[9]), .ZN(n369) );
  INVX0 U307 ( .INP(A[7]), .ZN(n360) );
  NAND2X0 U308 ( .IN1(A[7]), .IN2(n367), .QN(n113) );
  NAND2X0 U309 ( .IN1(n291), .IN2(n292), .QN(n259) );
  NOR2X0 U310 ( .IN1(n263), .IN2(n264), .QN(n262) );
  NAND2X0 U311 ( .IN1(A[8]), .IN2(n326), .QN(n110) );
  INVX0 U312 ( .INP(A[8]), .ZN(n368) );
  NAND2X0 U313 ( .IN1(n157), .IN2(n229), .QN(n339) );
  NAND2X1 U314 ( .IN1(n95), .IN2(n227), .QN(DIFF[0]) );
  NAND2X1 U315 ( .IN1(n341), .IN2(n342), .QN(n291) );
  NOR2X0 U316 ( .IN1(n343), .IN2(n344), .QN(n342) );
  NOR2X0 U317 ( .IN1(n345), .IN2(n346), .QN(n344) );
  NAND2X0 U318 ( .IN1(n274), .IN2(n271), .QN(n273) );
  NAND2X0 U319 ( .IN1(n270), .IN2(n274), .QN(n302) );
  NAND2X1 U320 ( .IN1(B[14]), .IN2(n303), .QN(n274) );
  NOR2X0 U321 ( .IN1(n267), .IN2(n268), .QN(n266) );
  NOR2X0 U322 ( .IN1(n272), .IN2(n273), .QN(n267) );
  INVX0 U323 ( .INP(A[2]), .ZN(n355) );
  NAND2X0 U324 ( .IN1(A[2]), .IN2(n352), .QN(n136) );
  NAND2X0 U325 ( .IN1(n216), .IN2(n217), .QN(n212) );
  NOR2X0 U326 ( .IN1(n253), .IN2(n246), .QN(n252) );
  NAND2X0 U327 ( .IN1(n246), .IN2(n247), .QN(n244) );
  NOR2X0 U328 ( .IN1(n287), .IN2(n286), .QN(n280) );
  INVX0 U329 ( .INP(n254), .ZN(n246) );
  INVX0 U330 ( .INP(A[14]), .ZN(n303) );
  NOR2X0 U331 ( .IN1(n324), .IN2(n105), .QN(n322) );
  INVX0 U332 ( .INP(A[3]), .ZN(n354) );
  NAND2X0 U333 ( .IN1(A[3]), .IN2(n349), .QN(n135) );
  NAND2X0 U334 ( .IN1(A[13]), .IN2(n310), .QN(n272) );
  INVX0 U335 ( .INP(A[13]), .ZN(n309) );
  INVX0 U336 ( .INP(A[15]), .ZN(n300) );
  NOR2X0 U337 ( .IN1(n365), .IN2(n364), .QN(n361) );
  NOR2X0 U338 ( .IN1(n36), .IN2(n120), .QN(n365) );
  NOR2X0 U339 ( .IN1(n293), .IN2(n290), .QN(n292) );
  NAND2X0 U340 ( .IN1(n276), .IN2(n289), .QN(n286) );
  NAND2X0 U341 ( .IN1(n275), .IN2(n276), .QN(n265) );
  NAND2X0 U342 ( .IN1(n284), .IN2(n108), .QN(n316) );
  NAND2X0 U343 ( .IN1(n284), .IN2(n56), .QN(n287) );
  NAND2X0 U344 ( .IN1(n284), .IN2(n276), .QN(n283) );
  NAND2X0 U345 ( .IN1(n284), .IN2(n289), .QN(n293) );
  NAND2X0 U346 ( .IN1(A[11]), .IN2(n89), .QN(n320) );
  INVX0 U347 ( .INP(A[17]), .ZN(n257) );
  NAND2X0 U348 ( .IN1(n218), .IN2(n219), .QN(n216) );
  NOR2X0 U349 ( .IN1(n322), .IN2(n323), .QN(n321) );
  NOR2X0 U350 ( .IN1(n282), .IN2(n283), .QN(n281) );
  NAND2X0 U351 ( .IN1(A[12]), .IN2(n87), .QN(n277) );
  INVX0 U352 ( .INP(A[10]), .ZN(n318) );
  INVX0 U353 ( .INP(n325), .ZN(n324) );
  NAND2X0 U354 ( .IN1(A[6]), .IN2(n88), .QN(n115) );
  NOR2X0 U355 ( .IN1(n215), .IN2(n212), .QN(n214) );
  NAND2X1 U356 ( .IN1(n233), .IN2(n234), .QN(n218) );
  NOR2X0 U357 ( .IN1(n280), .IN2(n281), .QN(n261) );
  INVX0 U358 ( .INP(A[0]), .ZN(n372) );
  INVX0 U359 ( .INP(n196), .ZN(n198) );
  NAND2X0 U360 ( .IN1(A[1]), .IN2(n356), .QN(n154) );
  NAND2X0 U361 ( .IN1(A[10]), .IN2(n371), .QN(n328) );
  NOR2X0 U362 ( .IN1(B[10]), .IN2(n318), .QN(n323) );
  NAND2X1 U363 ( .IN1(B[10]), .IN2(n318), .QN(n325) );
  NAND2X0 U364 ( .IN1(n285), .IN2(n112), .QN(n282) );
  NAND2X0 U365 ( .IN1(A[14]), .IN2(n304), .QN(n270) );
  NAND2X0 U366 ( .IN1(n200), .IN2(n201), .QN(n196) );
  NAND2X0 U367 ( .IN1(n188), .IN2(n189), .QN(n187) );
  NOR2X0 U368 ( .IN1(n243), .IN2(n235), .QN(n242) );
  NAND2X0 U369 ( .IN1(n194), .IN2(n195), .QN(n188) );
  NAND2X0 U370 ( .IN1(n236), .IN2(n235), .QN(n233) );
  NAND2X0 U371 ( .IN1(n196), .IN2(n197), .QN(n195) );
  NAND2X0 U372 ( .IN1(A[17]), .IN2(n256), .QN(n245) );
  NAND2X0 U373 ( .IN1(n65), .IN2(n171), .QN(n170) );
  NAND2X0 U374 ( .IN1(n141), .IN2(n142), .QN(n140) );
  XOR2X1 U375 ( .IN1(n101), .IN2(n102), .Q(DIFF[9]) );
  XOR2X1 U376 ( .IN1(n106), .IN2(n107), .Q(DIFF[8]) );
  XOR2X1 U377 ( .IN1(n111), .IN2(n86), .Q(DIFF[7]) );
  XOR2X1 U378 ( .IN1(n118), .IN2(n119), .Q(DIFF[6]) );
  XOR2X1 U379 ( .IN1(n124), .IN2(n125), .Q(DIFF[5]) );
  XOR2X1 U380 ( .IN1(n130), .IN2(n131), .Q(DIFF[4]) );
  XOR2X1 U381 ( .IN1(n133), .IN2(n83), .Q(DIFF[3]) );
  XOR2X1 U382 ( .IN1(n138), .IN2(n151), .Q(DIFF[2]) );
  XOR2X1 U383 ( .IN1(n4), .IN2(n166), .Q(DIFF[27]) );
  XOR2X1 U384 ( .IN1(n3), .IN2(n172), .Q(DIFF[26]) );
  XOR2X1 U385 ( .IN1(n7), .IN2(n178), .Q(DIFF[25]) );
  XOR2X1 U386 ( .IN1(n5), .IN2(n183), .Q(DIFF[24]) );
  XOR2X1 U387 ( .IN1(n190), .IN2(n191), .Q(DIFF[23]) );
  XOR2X1 U388 ( .IN1(n198), .IN2(n199), .Q(DIFF[22]) );
  XOR2X1 U389 ( .IN1(n203), .IN2(n6), .Q(DIFF[21]) );
  XOR2X1 U390 ( .IN1(n213), .IN2(n214), .Q(DIFF[20]) );
  XOR2X1 U391 ( .IN1(n225), .IN2(n226), .Q(DIFF[1]) );
  XOR2X1 U392 ( .IN1(n230), .IN2(n231), .Q(DIFF[19]) );
  XOR2X1 U393 ( .IN1(n241), .IN2(n242), .Q(DIFF[18]) );
  XOR2X1 U394 ( .IN1(n251), .IN2(n252), .Q(DIFF[17]) );
  XOR2X1 U395 ( .IN1(n258), .IN2(n220), .Q(DIFF[16]) );
  NAND4X0 U396 ( .IN1(n262), .IN2(n260), .IN3(n261), .IN4(n259), .QN(n208) );
  NAND4X0 U397 ( .IN1(n294), .IN2(n295), .IN3(n274), .IN4(n271), .QN(n290) );
  XOR2X1 U398 ( .IN1(n298), .IN2(n85), .Q(DIFF[15]) );
  XOR2X1 U399 ( .IN1(n2), .IN2(n302), .Q(DIFF[14]) );
  XOR2X1 U400 ( .IN1(n307), .IN2(n308), .Q(DIFF[13]) );
  XOR2X1 U401 ( .IN1(n313), .IN2(n314), .Q(DIFF[12]) );
  NAND3X0 U402 ( .IN1(n321), .IN2(n320), .IN3(n319), .QN(n279) );
  NAND4X0 U403 ( .IN1(A[8]), .IN2(n325), .IN3(n104), .IN4(n326), .QN(n319) );
  XOR2X1 U404 ( .IN1(n327), .IN2(n84), .Q(DIFF[11]) );
  XOR2X1 U405 ( .IN1(n331), .IN2(n332), .Q(DIFF[10]) );
  NAND4X0 U406 ( .IN1(A[4]), .IN2(n117), .IN3(n123), .IN4(n132), .QN(n362) );
endmodule


module BoothMultiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313;

  AND2X1 U2 ( .IN1(B[28]), .IN2(A[28]), .Q(n22) );
  AND2X1 U3 ( .IN1(n33), .IN2(n34), .Q(n23) );
  AND2X1 U4 ( .IN1(n190), .IN2(n198), .Q(n62) );
  AND2X1 U5 ( .IN1(n165), .IN2(n162), .Q(n58) );
  OR2X1 U6 ( .IN1(A[10]), .IN2(B[10]), .Q(n282) );
  AND2X1 U7 ( .IN1(B[16]), .IN2(A[16]), .Q(n66) );
  NBUFFX2 U8 ( .INP(n228), .Z(n60) );
  OR2X1 U9 ( .IN1(B[25]), .IN2(A[25]), .Q(n170) );
  INVX0 U10 ( .INP(n164), .ZN(n28) );
  AND2X1 U11 ( .IN1(n31), .IN2(n282), .Q(n289) );
  XOR3X1 U12 ( .IN1(B[29]), .IN2(A[29]), .IN3(n149), .Q(SUM[29]) );
  XOR3X1 U13 ( .IN1(B[30]), .IN2(A[30]), .IN3(n143), .Q(SUM[30]) );
  AND2X1 U14 ( .IN1(n167), .IN2(n168), .Q(n1) );
  AND2X1 U15 ( .IN1(n182), .IN2(n183), .Q(n2) );
  AND2X1 U16 ( .IN1(B[1]), .IN2(A[1]), .Q(n3) );
  AND2X1 U17 ( .IN1(n212), .IN2(n211), .Q(SUM[0]) );
  NAND2X0 U18 ( .IN1(B[1]), .IN2(A[1]), .QN(n5) );
  OR2X1 U19 ( .IN1(A[3]), .IN2(B[3]), .Q(n6) );
  OR2X1 U20 ( .IN1(B[8]), .IN2(A[8]), .Q(n109) );
  OR2X1 U21 ( .IN1(A[3]), .IN2(B[3]), .Q(n303) );
  NOR2X0 U22 ( .IN1(A[1]), .IN2(B[1]), .QN(n95) );
  NAND2X0 U23 ( .IN1(n105), .IN2(n109), .QN(n7) );
  NOR2X0 U24 ( .IN1(n8), .IN2(n9), .QN(n195) );
  NAND2X0 U25 ( .IN1(n70), .IN2(n71), .QN(n8) );
  NOR2X0 U26 ( .IN1(n98), .IN2(n206), .QN(n9) );
  AND2X1 U27 ( .IN1(n165), .IN2(n170), .Q(n10) );
  NAND2X0 U28 ( .IN1(n165), .IN2(n82), .QN(n11) );
  AND2X1 U29 ( .IN1(n34), .IN2(n14), .Q(n12) );
  NOR2X0 U30 ( .IN1(n12), .IN2(n13), .QN(n51) );
  AND2X1 U31 ( .IN1(n54), .IN2(n22), .Q(n13) );
  AND2X1 U32 ( .IN1(n33), .IN2(n54), .Q(n14) );
  NAND2X0 U33 ( .IN1(n160), .IN2(n162), .QN(n163) );
  NAND2X0 U34 ( .IN1(B[27]), .IN2(A[27]), .QN(n160) );
  OR2X1 U35 ( .IN1(B[28]), .IN2(A[28]), .Q(n158) );
  NAND2X0 U36 ( .IN1(n184), .IN2(n87), .QN(n15) );
  NAND2X0 U37 ( .IN1(n15), .IN2(n16), .QN(n59) );
  AND2X1 U38 ( .IN1(n178), .IN2(n85), .Q(n16) );
  NAND3X1 U39 ( .IN1(n139), .IN2(n6), .IN3(n3), .QN(n296) );
  NOR2X0 U40 ( .IN1(n90), .IN2(n91), .QN(n17) );
  NAND2X1 U41 ( .IN1(n225), .IN2(n226), .QN(n218) );
  NAND2X0 U42 ( .IN1(n208), .IN2(n198), .QN(n18) );
  INVX0 U43 ( .INP(A[19]), .ZN(n19) );
  INVX0 U44 ( .INP(n19), .ZN(n20) );
  NOR2X0 U45 ( .IN1(A[6]), .IN2(B[6]), .QN(n100) );
  AND2X1 U46 ( .IN1(n141), .IN2(n52), .Q(n21) );
  OR2X1 U47 ( .IN1(n22), .IN2(n23), .Q(n149) );
  INVX0 U48 ( .INP(n98), .ZN(n24) );
  NAND2X0 U49 ( .IN1(n312), .IN2(n313), .QN(n117) );
  INVX0 U50 ( .INP(n88), .ZN(n25) );
  NAND2X0 U51 ( .IN1(n168), .IN2(n29), .QN(n26) );
  NAND2X0 U52 ( .IN1(n26), .IN2(n27), .QN(n32) );
  OR2X1 U53 ( .IN1(n28), .IN2(n165), .Q(n27) );
  AND2X1 U54 ( .IN1(n167), .IN2(n164), .Q(n29) );
  XOR3X1 U55 ( .IN1(B[28]), .IN2(A[28]), .IN3(n159), .Q(SUM[28]) );
  AND2X1 U56 ( .IN1(n30), .IN2(n31), .Q(n281) );
  NAND2X0 U57 ( .IN1(n278), .IN2(n73), .QN(n30) );
  NAND2X0 U58 ( .IN1(B[10]), .IN2(A[10]), .QN(n31) );
  NAND2X0 U59 ( .IN1(B[25]), .IN2(A[25]), .QN(n167) );
  NAND2X0 U60 ( .IN1(n179), .IN2(n36), .QN(n33) );
  OR2X1 U61 ( .IN1(n35), .IN2(n37), .Q(n34) );
  INVX0 U62 ( .INP(n80), .ZN(n35) );
  AND2X1 U63 ( .IN1(n39), .IN2(n80), .Q(n36) );
  OR2X1 U64 ( .IN1(n38), .IN2(n40), .Q(n37) );
  INVX0 U65 ( .INP(n74), .ZN(n38) );
  AND2X1 U66 ( .IN1(n42), .IN2(n74), .Q(n39) );
  OR2X1 U67 ( .IN1(n41), .IN2(n44), .Q(n40) );
  INVX0 U68 ( .INP(n68), .ZN(n41) );
  AND2X1 U69 ( .IN1(n46), .IN2(n68), .Q(n42) );
  NAND2X0 U70 ( .IN1(n195), .IN2(n196), .QN(n43) );
  AND2X1 U71 ( .IN1(n303), .IN2(n139), .Q(n298) );
  OR2X1 U72 ( .IN1(n45), .IN2(n65), .Q(n44) );
  INVX0 U73 ( .INP(n63), .ZN(n45) );
  AND2X1 U74 ( .IN1(n178), .IN2(n63), .Q(n46) );
  XOR3X1 U75 ( .IN1(B[31]), .IN2(A[31]), .IN3(n140), .Q(SUM[31]) );
  NAND2X1 U76 ( .IN1(n237), .IN2(n238), .QN(n236) );
  NAND2X0 U77 ( .IN1(n169), .IN2(n50), .QN(n47) );
  AND2X1 U78 ( .IN1(n47), .IN2(n48), .Q(n55) );
  OR2X1 U79 ( .IN1(n49), .IN2(n167), .Q(n48) );
  INVX0 U80 ( .INP(n58), .ZN(n49) );
  AND2X1 U81 ( .IN1(n170), .IN2(n58), .Q(n50) );
  OR2X1 U82 ( .IN1(n53), .IN2(n146), .Q(n52) );
  INVX0 U83 ( .INP(n142), .ZN(n53) );
  AND2X1 U84 ( .IN1(n148), .IN2(n142), .Q(n54) );
  AND2X1 U85 ( .IN1(n55), .IN2(n56), .Q(n161) );
  OR2X1 U86 ( .IN1(n57), .IN2(n164), .Q(n56) );
  INVX0 U87 ( .INP(n162), .ZN(n57) );
  NOR2X0 U88 ( .IN1(n209), .IN2(n88), .QN(n61) );
  NAND2X0 U89 ( .IN1(n61), .IN2(n62), .QN(n79) );
  OR2X1 U90 ( .IN1(n64), .IN2(n173), .Q(n63) );
  INVX0 U91 ( .INP(n69), .ZN(n64) );
  AND2X1 U92 ( .IN1(n175), .IN2(n69), .Q(n65) );
  NAND2X0 U93 ( .IN1(n188), .IN2(n189), .QN(n67) );
  OR2X1 U94 ( .IN1(n11), .IN2(n167), .Q(n68) );
  AND2X1 U95 ( .IN1(n82), .IN2(n10), .Q(n69) );
  NAND2X0 U96 ( .IN1(n218), .IN2(n72), .QN(n70) );
  OR2X1 U97 ( .IN1(n18), .IN2(n217), .Q(n71) );
  AND2X1 U98 ( .IN1(n219), .IN2(n99), .Q(n72) );
  AND2X1 U99 ( .IN1(A[9]), .IN2(B[9]), .Q(n73) );
  OR2X1 U100 ( .IN1(n75), .IN2(n164), .Q(n74) );
  INVX0 U101 ( .INP(n82), .ZN(n75) );
  NOR2X0 U102 ( .IN1(n199), .IN2(n79), .QN(n76) );
  NOR2X0 U103 ( .IN1(n76), .IN2(n77), .QN(n189) );
  AND2X1 U104 ( .IN1(n78), .IN2(n194), .Q(n77) );
  INVX0 U105 ( .INP(n83), .ZN(n78) );
  OR2X1 U106 ( .IN1(B[21]), .IN2(A[21]), .Q(n190) );
  NAND2X0 U107 ( .IN1(n195), .IN2(n196), .QN(n194) );
  OR2X1 U108 ( .IN1(n81), .IN2(n160), .Q(n80) );
  INVX0 U109 ( .INP(n158), .ZN(n81) );
  AND2X1 U110 ( .IN1(n162), .IN2(n158), .Q(n82) );
  NOR2X0 U111 ( .IN1(B[21]), .IN2(A[21]), .QN(n83) );
  NAND2X0 U112 ( .IN1(n278), .IN2(n246), .QN(n91) );
  NAND2X0 U113 ( .IN1(n105), .IN2(n102), .QN(n290) );
  NAND2X0 U114 ( .IN1(n114), .IN2(n115), .QN(n111) );
  NAND2X0 U115 ( .IN1(n288), .IN2(n282), .QN(n287) );
  NAND2X0 U116 ( .IN1(n25), .IN2(n206), .QN(n213) );
  NAND2X0 U117 ( .IN1(n190), .IN2(n188), .QN(n192) );
  NAND2X0 U118 ( .IN1(n185), .IN2(n182), .QN(n186) );
  NAND2X0 U119 ( .IN1(n24), .IN2(n196), .QN(n202) );
  NAND2X0 U120 ( .IN1(n219), .IN2(n217), .QN(n222) );
  NAND2X0 U121 ( .IN1(n126), .IN2(n128), .QN(n130) );
  NAND2X0 U122 ( .IN1(B[19]), .IN2(n20), .QN(n206) );
  NAND2X0 U123 ( .IN1(n184), .IN2(n87), .QN(n84) );
  AND2X1 U124 ( .IN1(n84), .IN2(n85), .Q(n179) );
  OR2X1 U125 ( .IN1(n86), .IN2(n182), .Q(n85) );
  INVX0 U126 ( .INP(n180), .ZN(n86) );
  AND2X1 U127 ( .IN1(n185), .IN2(n180), .Q(n87) );
  NOR2X0 U128 ( .IN1(B[19]), .IN2(n20), .QN(n88) );
  AND2X1 U129 ( .IN1(n251), .IN2(n252), .Q(n89) );
  INVX0 U130 ( .INP(n294), .ZN(n129) );
  INVX0 U131 ( .INP(n122), .ZN(n124) );
  NAND2X0 U132 ( .IN1(n123), .IN2(n128), .QN(n304) );
  INVX0 U133 ( .INP(n263), .ZN(n260) );
  AND2X1 U134 ( .IN1(n208), .IN2(n198), .Q(n99) );
  INVX0 U135 ( .INP(n267), .ZN(n258) );
  INVX0 U136 ( .INP(n136), .ZN(n153) );
  NOR2X0 U137 ( .IN1(n7), .IN2(n91), .QN(n240) );
  NAND2X0 U138 ( .IN1(n105), .IN2(n109), .QN(n90) );
  OR2X1 U139 ( .IN1(n209), .IN2(n88), .Q(n201) );
  NAND2X0 U140 ( .IN1(n61), .IN2(n24), .QN(n200) );
  NAND2X0 U141 ( .IN1(n255), .IN2(n256), .QN(n248) );
  NAND3X0 U142 ( .IN1(n257), .IN2(n258), .IN3(n259), .QN(n256) );
  NAND2X0 U143 ( .IN1(n260), .IN2(n257), .QN(n255) );
  NAND2X0 U144 ( .IN1(n272), .IN2(n250), .QN(n269) );
  NAND2X0 U145 ( .IN1(n292), .IN2(n293), .QN(n107) );
  NAND2X1 U146 ( .IN1(n126), .IN2(n127), .QN(n122) );
  NAND2X0 U147 ( .IN1(n128), .IN2(n129), .QN(n127) );
  NAND2X1 U148 ( .IN1(n110), .IN2(n291), .QN(n102) );
  NAND2X0 U149 ( .IN1(n109), .IN2(n107), .QN(n291) );
  NOR2X0 U150 ( .IN1(n231), .IN2(n66), .QN(n230) );
  INVX0 U151 ( .INP(n60), .ZN(n233) );
  NOR2X0 U152 ( .IN1(n204), .IN2(n197), .QN(n203) );
  NAND2X0 U153 ( .IN1(n276), .IN2(n277), .QN(n273) );
  NAND2X0 U154 ( .IN1(n120), .IN2(n121), .QN(n116) );
  NAND2X1 U155 ( .IN1(n122), .IN2(n97), .QN(n121) );
  NAND2X0 U156 ( .IN1(n31), .IN2(n287), .QN(n286) );
  NAND2X0 U157 ( .IN1(n263), .IN2(n264), .QN(n261) );
  NAND2X0 U158 ( .IN1(n267), .IN2(n268), .QN(n265) );
  NAND2X0 U159 ( .IN1(n269), .IN2(n270), .QN(n268) );
  INVX0 U160 ( .INP(n135), .ZN(n133) );
  INVX0 U161 ( .INP(n211), .ZN(n156) );
  NAND2X0 U162 ( .IN1(n157), .IN2(n5), .QN(n210) );
  NOR2X0 U163 ( .IN1(n119), .IN2(n100), .QN(n118) );
  INVX0 U164 ( .INP(n115), .ZN(n119) );
  NAND2X0 U165 ( .IN1(n120), .IN2(n96), .QN(n125) );
  NAND2X0 U166 ( .IN1(n301), .IN2(n302), .QN(n157) );
  NOR2X0 U167 ( .IN1(n260), .IN2(n253), .QN(n266) );
  NOR2X0 U168 ( .IN1(n73), .IN2(n104), .QN(n103) );
  INVX0 U169 ( .INP(n105), .ZN(n104) );
  AND2X1 U170 ( .IN1(n110), .IN2(n109), .Q(n108) );
  AND2X1 U171 ( .IN1(n238), .IN2(n257), .Q(n262) );
  NAND2X0 U172 ( .IN1(n136), .IN2(n137), .QN(n131) );
  NOR2X0 U173 ( .IN1(n258), .IN2(n254), .QN(n271) );
  INVX0 U174 ( .INP(n270), .ZN(n254) );
  NAND2X0 U175 ( .IN1(n5), .IN2(n155), .QN(n138) );
  NAND2X1 U176 ( .IN1(n156), .IN2(n157), .QN(n155) );
  AND2X1 U177 ( .IN1(n250), .IN2(n274), .Q(n275) );
  NAND2X1 U178 ( .IN1(n178), .IN2(n180), .QN(n181) );
  NAND2X1 U179 ( .IN1(n173), .IN2(n175), .QN(n177) );
  NAND2X1 U180 ( .IN1(n167), .IN2(n170), .QN(n172) );
  NAND2X1 U181 ( .IN1(n164), .IN2(n165), .QN(n166) );
  AND2X1 U182 ( .IN1(n112), .IN2(n113), .Q(n92) );
  AND2X1 U183 ( .IN1(n246), .IN2(n280), .Q(n93) );
  OR2X1 U184 ( .IN1(B[15]), .IN2(A[15]), .Q(n257) );
  NAND2X0 U185 ( .IN1(n113), .IN2(n115), .QN(n310) );
  OR2X1 U186 ( .IN1(B[13]), .IN2(A[13]), .Q(n270) );
  OR2X1 U187 ( .IN1(A[10]), .IN2(B[10]), .Q(n278) );
  OR2X1 U188 ( .IN1(B[4]), .IN2(A[4]), .Q(n128) );
  OR2X1 U189 ( .IN1(B[16]), .IN2(A[16]), .Q(n228) );
  NAND2X1 U190 ( .IN1(B[29]), .IN2(A[29]), .QN(n146) );
  NAND2X1 U191 ( .IN1(n150), .IN2(n151), .QN(n148) );
  NAND2X1 U192 ( .IN1(B[30]), .IN2(A[30]), .QN(n141) );
  NAND2X1 U193 ( .IN1(n144), .IN2(n145), .QN(n142) );
  OR2X1 U194 ( .IN1(B[14]), .IN2(A[14]), .Q(n259) );
  OR2X1 U195 ( .IN1(B[12]), .IN2(A[12]), .Q(n274) );
  OR2X1 U196 ( .IN1(A[20]), .IN2(B[20]), .Q(n198) );
  OR2X1 U197 ( .IN1(B[9]), .IN2(A[9]), .Q(n105) );
  OR2X1 U198 ( .IN1(B[7]), .IN2(A[7]), .Q(n112) );
  NAND2X0 U199 ( .IN1(B[18]), .IN2(A[18]), .QN(n217) );
  OR2X1 U200 ( .IN1(B[11]), .IN2(A[11]), .Q(n246) );
  OR2X1 U201 ( .IN1(B[18]), .IN2(A[18]), .Q(n219) );
  OR2X1 U202 ( .IN1(B[19]), .IN2(A[19]), .Q(n208) );
  OR2X1 U203 ( .IN1(A[2]), .IN2(B[2]), .Q(n139) );
  OR2X1 U204 ( .IN1(A[17]), .IN2(B[17]), .Q(n227) );
  NAND2X0 U205 ( .IN1(B[20]), .IN2(A[20]), .QN(n196) );
  NAND2X0 U206 ( .IN1(B[22]), .IN2(A[22]), .QN(n182) );
  NAND2X0 U207 ( .IN1(B[21]), .IN2(A[21]), .QN(n188) );
  NAND2X1 U208 ( .IN1(B[23]), .IN2(A[23]), .QN(n178) );
  NAND2X1 U209 ( .IN1(B[24]), .IN2(A[24]), .QN(n173) );
  NAND2X1 U210 ( .IN1(B[26]), .IN2(A[26]), .QN(n164) );
  OR2X1 U211 ( .IN1(B[26]), .IN2(A[26]), .Q(n165) );
  OR2X1 U212 ( .IN1(B[24]), .IN2(A[24]), .Q(n175) );
  OR2X1 U213 ( .IN1(B[23]), .IN2(A[23]), .Q(n180) );
  OR2X1 U214 ( .IN1(B[27]), .IN2(A[27]), .Q(n162) );
  OR2X1 U215 ( .IN1(B[22]), .IN2(A[22]), .Q(n185) );
  OR2X1 U216 ( .IN1(B[0]), .IN2(A[0]), .Q(n212) );
  INVX0 U217 ( .INP(A[30]), .ZN(n145) );
  INVX0 U218 ( .INP(A[29]), .ZN(n151) );
  INVX0 U219 ( .INP(B[30]), .ZN(n144) );
  INVX0 U220 ( .INP(B[29]), .ZN(n150) );
  INVX0 U221 ( .INP(B[8]), .ZN(n285) );
  INVX0 U222 ( .INP(B[5]), .ZN(n308) );
  NAND3X0 U223 ( .IN1(n242), .IN2(n243), .IN3(n244), .QN(n235) );
  INVX0 U224 ( .INP(n59), .ZN(n176) );
  NOR2X0 U225 ( .IN1(n235), .IN2(n236), .QN(n94) );
  NAND2X0 U226 ( .IN1(B[0]), .IN2(A[0]), .QN(n300) );
  NAND2X0 U227 ( .IN1(B[0]), .IN2(A[0]), .QN(n211) );
  NOR2X0 U228 ( .IN1(n133), .IN2(n134), .QN(n132) );
  NAND2X0 U229 ( .IN1(n239), .IN2(n129), .QN(n293) );
  NOR2X0 U230 ( .IN1(n304), .IN2(n305), .QN(n239) );
  NOR2X0 U231 ( .IN1(n153), .IN2(n154), .QN(n152) );
  NAND2X0 U232 ( .IN1(n106), .IN2(n290), .QN(n288) );
  NAND2X0 U233 ( .IN1(B[9]), .IN2(A[9]), .QN(n106) );
  INVX0 U234 ( .INP(n6), .ZN(n134) );
  NAND2X0 U235 ( .IN1(n153), .IN2(n6), .QN(n295) );
  NAND2X0 U236 ( .IN1(n265), .IN2(n259), .QN(n264) );
  INVX0 U237 ( .INP(n259), .ZN(n253) );
  AND2X1 U238 ( .IN1(n257), .IN2(n259), .Q(n252) );
  NAND2X0 U239 ( .IN1(n138), .IN2(n139), .QN(n137) );
  INVX0 U240 ( .INP(n139), .ZN(n154) );
  NOR2X0 U241 ( .IN1(n120), .IN2(n100), .QN(n311) );
  NAND2X0 U242 ( .IN1(B[5]), .IN2(A[5]), .QN(n120) );
  INVX0 U243 ( .INP(B[1]), .ZN(n301) );
  INVX0 U244 ( .INP(A[1]), .ZN(n302) );
  NAND2X0 U245 ( .IN1(n17), .IN2(n107), .QN(n277) );
  NAND2X0 U246 ( .IN1(n308), .IN2(n309), .QN(n96) );
  NAND2X0 U247 ( .IN1(n308), .IN2(n309), .QN(n97) );
  NAND2X0 U248 ( .IN1(n308), .IN2(n309), .QN(n123) );
  INVX0 U249 ( .INP(A[5]), .ZN(n309) );
  INVX0 U250 ( .INP(n198), .ZN(n98) );
  NAND2X0 U251 ( .IN1(B[4]), .IN2(A[4]), .QN(n126) );
  NOR2X0 U252 ( .IN1(n284), .IN2(n285), .QN(n283) );
  AND2X1 U253 ( .IN1(n270), .IN2(n274), .Q(n251) );
  NAND2X1 U254 ( .IN1(n205), .IN2(n206), .QN(n197) );
  NOR2X0 U255 ( .IN1(n95), .IN2(n300), .QN(n299) );
  NAND2X0 U256 ( .IN1(B[7]), .IN2(A[7]), .QN(n113) );
  INVX0 U257 ( .INP(B[6]), .ZN(n312) );
  NAND2X0 U258 ( .IN1(B[8]), .IN2(A[8]), .QN(n110) );
  INVX0 U259 ( .INP(A[8]), .ZN(n284) );
  NAND2X0 U260 ( .IN1(n251), .IN2(n252), .QN(n101) );
  NAND2X0 U261 ( .IN1(n220), .IN2(n219), .QN(n209) );
  INVX0 U262 ( .INP(n221), .ZN(n220) );
  NAND2X0 U263 ( .IN1(B[2]), .IN2(A[2]), .QN(n136) );
  NOR2X0 U264 ( .IN1(n235), .IN2(n236), .QN(n199) );
  NAND2X0 U265 ( .IN1(n247), .IN2(n246), .QN(n276) );
  NAND2X0 U266 ( .IN1(B[3]), .IN2(A[3]), .QN(n135) );
  NAND2X0 U267 ( .IN1(B[13]), .IN2(A[13]), .QN(n267) );
  NOR2X0 U268 ( .IN1(n311), .IN2(n310), .QN(n306) );
  NAND2X0 U269 ( .IN1(B[15]), .IN2(A[15]), .QN(n238) );
  NOR2X0 U270 ( .IN1(n215), .IN2(n207), .QN(n214) );
  NAND2X0 U271 ( .IN1(n207), .IN2(n25), .QN(n205) );
  NAND2X0 U272 ( .IN1(n216), .IN2(n217), .QN(n207) );
  NAND2X0 U273 ( .IN1(n298), .IN2(n299), .QN(n297) );
  NAND2X0 U274 ( .IN1(n306), .IN2(n307), .QN(n245) );
  INVX0 U275 ( .INP(n241), .ZN(n294) );
  NAND2X0 U276 ( .IN1(B[11]), .IN2(A[11]), .QN(n280) );
  NOR2X0 U277 ( .IN1(n249), .IN2(n248), .QN(n242) );
  NAND2X0 U278 ( .IN1(n245), .IN2(n112), .QN(n292) );
  INVX0 U279 ( .INP(n67), .ZN(n187) );
  NAND2X0 U280 ( .IN1(n273), .IN2(n274), .QN(n272) );
  NOR2X0 U281 ( .IN1(n101), .IN2(n250), .QN(n249) );
  NAND2X0 U282 ( .IN1(B[12]), .IN2(A[12]), .QN(n250) );
  INVX0 U283 ( .INP(n169), .ZN(n171) );
  NAND2X0 U284 ( .IN1(n116), .IN2(n117), .QN(n114) );
  NAND2X0 U285 ( .IN1(n169), .IN2(n170), .QN(n168) );
  NAND2X0 U286 ( .IN1(n112), .IN2(n117), .QN(n305) );
  NAND2X0 U287 ( .IN1(n173), .IN2(n174), .QN(n169) );
  NOR2X0 U288 ( .IN1(n224), .IN2(n218), .QN(n223) );
  NAND2X0 U289 ( .IN1(n59), .IN2(n175), .QN(n174) );
  NAND2X0 U290 ( .IN1(n218), .IN2(n219), .QN(n216) );
  INVX0 U291 ( .INP(A[6]), .ZN(n313) );
  NAND2X0 U292 ( .IN1(B[14]), .IN2(A[14]), .QN(n263) );
  NAND2X0 U293 ( .IN1(n60), .IN2(n232), .QN(n234) );
  NAND2X0 U294 ( .IN1(n188), .IN2(n189), .QN(n184) );
  NAND2X0 U295 ( .IN1(n67), .IN2(n185), .QN(n183) );
  NAND2X0 U296 ( .IN1(B[6]), .IN2(A[6]), .QN(n115) );
  NAND2X0 U297 ( .IN1(n160), .IN2(n161), .QN(n159) );
  NOR2X0 U298 ( .IN1(n94), .IN2(n201), .QN(n204) );
  NOR2X0 U299 ( .IN1(n94), .IN2(n209), .QN(n215) );
  NOR2X0 U300 ( .IN1(n94), .IN2(n221), .QN(n224) );
  NOR2X0 U301 ( .IN1(n233), .IN2(n94), .QN(n231) );
  NOR2X0 U302 ( .IN1(n193), .IN2(n43), .QN(n191) );
  NAND2X0 U303 ( .IN1(n227), .IN2(n226), .QN(n229) );
  NAND2X0 U304 ( .IN1(n51), .IN2(n21), .QN(n140) );
  NAND2X0 U305 ( .IN1(n228), .IN2(n227), .QN(n221) );
  NAND2X0 U306 ( .IN1(n66), .IN2(n227), .QN(n225) );
  NAND2X0 U307 ( .IN1(B[17]), .IN2(A[17]), .QN(n226) );
  NAND2X0 U308 ( .IN1(n146), .IN2(n147), .QN(n143) );
  NAND2X0 U309 ( .IN1(B[16]), .IN2(A[16]), .QN(n232) );
  NAND2X0 U310 ( .IN1(n148), .IN2(n149), .QN(n147) );
  NOR2X0 U311 ( .IN1(n94), .IN2(n200), .QN(n193) );
  XOR2X1 U312 ( .IN1(n102), .IN2(n103), .Q(SUM[9]) );
  XOR2X1 U313 ( .IN1(n107), .IN2(n108), .Q(SUM[8]) );
  XOR2X1 U314 ( .IN1(n111), .IN2(n92), .Q(SUM[7]) );
  XOR2X1 U315 ( .IN1(n116), .IN2(n118), .Q(SUM[6]) );
  XOR2X1 U316 ( .IN1(n124), .IN2(n125), .Q(SUM[5]) );
  XOR2X1 U317 ( .IN1(n294), .IN2(n130), .Q(SUM[4]) );
  XOR2X1 U318 ( .IN1(n131), .IN2(n132), .Q(SUM[3]) );
  XOR2X1 U319 ( .IN1(n138), .IN2(n152), .Q(SUM[2]) );
  XOR2X1 U320 ( .IN1(n32), .IN2(n163), .Q(SUM[27]) );
  XOR2X1 U321 ( .IN1(n1), .IN2(n166), .Q(SUM[26]) );
  XOR2X1 U322 ( .IN1(n171), .IN2(n172), .Q(SUM[25]) );
  XOR2X1 U323 ( .IN1(n176), .IN2(n177), .Q(SUM[24]) );
  XOR2X1 U324 ( .IN1(n2), .IN2(n181), .Q(SUM[23]) );
  XOR2X1 U325 ( .IN1(n186), .IN2(n187), .Q(SUM[22]) );
  XOR2X1 U326 ( .IN1(n192), .IN2(n191), .Q(SUM[21]) );
  XOR2X1 U327 ( .IN1(n202), .IN2(n203), .Q(SUM[20]) );
  XOR2X1 U328 ( .IN1(n210), .IN2(n211), .Q(SUM[1]) );
  XOR2X1 U329 ( .IN1(n213), .IN2(n214), .Q(SUM[19]) );
  XOR2X1 U330 ( .IN1(n222), .IN2(n223), .Q(SUM[18]) );
  XOR2X1 U331 ( .IN1(n229), .IN2(n230), .Q(SUM[17]) );
  XOR2X1 U332 ( .IN1(n234), .IN2(n94), .Q(SUM[16]) );
  NAND4X0 U333 ( .IN1(n241), .IN2(n89), .IN3(n17), .IN4(n239), .QN(n237) );
  NAND4X0 U334 ( .IN1(n240), .IN2(n89), .IN3(n245), .IN4(n112), .QN(n244) );
  NAND3X0 U335 ( .IN1(n89), .IN2(n246), .IN3(n247), .QN(n243) );
  XOR2X1 U336 ( .IN1(n261), .IN2(n262), .Q(SUM[15]) );
  XOR2X1 U337 ( .IN1(n265), .IN2(n266), .Q(SUM[14]) );
  XOR2X1 U338 ( .IN1(n269), .IN2(n271), .Q(SUM[13]) );
  XOR2X1 U339 ( .IN1(n273), .IN2(n275), .Q(SUM[12]) );
  NAND3X0 U340 ( .IN1(n281), .IN2(n280), .IN3(n279), .QN(n247) );
  NAND3X0 U341 ( .IN1(n282), .IN2(n105), .IN3(n283), .QN(n279) );
  XOR2X1 U342 ( .IN1(n286), .IN2(n93), .Q(SUM[11]) );
  XOR2X1 U343 ( .IN1(n288), .IN2(n289), .Q(SUM[10]) );
  NAND4X0 U344 ( .IN1(n297), .IN2(n296), .IN3(n295), .IN4(n135), .QN(n241) );
  NAND4X0 U345 ( .IN1(B[4]), .IN2(A[4]), .IN3(n96), .IN4(n117), .QN(n307) );
endmodule


module BoothMultiplier ( clk, oClk, rst, oRst, M, Q, P );
  input [31:0] M;
  input [31:0] Q;
  output [63:0] P;
  input clk, oClk, rst, oRst;
  wire   N4, N43, N44, N45, N46, N47, n140, n141, n142, n143, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n159,
         n160, n164, n165, n171, n172, n173, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433;
  wire   [31:0] Acc;
  wire   [31:0] Q_reg;
  wire   [5:0] count;
  wire   [31:0] M_reg;
  wire   [64:33] case_add;
  wire   [64:33] case_sub;

  LATCHX1 \M_reg_reg[31]  ( .CLK(n375), .D(M[31]), .Q(M_reg[31]) );
  LATCHX1 \M_reg_reg[30]  ( .CLK(n375), .D(M[30]), .Q(M_reg[30]) );
  LATCHX1 \M_reg_reg[29]  ( .CLK(n375), .D(M[29]), .Q(M_reg[29]) );
  LATCHX1 \M_reg_reg[28]  ( .CLK(n375), .D(M[28]), .Q(M_reg[28]) );
  LATCHX1 \M_reg_reg[27]  ( .CLK(n375), .D(M[27]), .Q(M_reg[27]) );
  LATCHX1 \M_reg_reg[26]  ( .CLK(n375), .D(M[26]), .Q(M_reg[26]) );
  LATCHX1 \M_reg_reg[25]  ( .CLK(n375), .D(M[25]), .Q(M_reg[25]) );
  LATCHX1 \M_reg_reg[24]  ( .CLK(n375), .D(M[24]), .Q(M_reg[24]) );
  LATCHX1 \M_reg_reg[23]  ( .CLK(n375), .D(M[23]), .Q(M_reg[23]) );
  LATCHX1 \M_reg_reg[22]  ( .CLK(n375), .D(M[22]), .Q(M_reg[22]) );
  LATCHX1 \M_reg_reg[21]  ( .CLK(n375), .D(M[21]), .Q(M_reg[21]) );
  LATCHX1 \M_reg_reg[20]  ( .CLK(n375), .D(M[20]), .Q(M_reg[20]) );
  LATCHX1 \M_reg_reg[19]  ( .CLK(n375), .D(M[19]), .Q(M_reg[19]) );
  LATCHX1 \M_reg_reg[18]  ( .CLK(n375), .D(M[18]), .Q(M_reg[18]) );
  LATCHX1 \M_reg_reg[17]  ( .CLK(n375), .D(M[17]), .Q(M_reg[17]) );
  LATCHX1 \M_reg_reg[16]  ( .CLK(n375), .D(M[16]), .Q(M_reg[16]) );
  LATCHX1 \M_reg_reg[15]  ( .CLK(n375), .D(M[15]), .Q(M_reg[15]) );
  LATCHX1 \M_reg_reg[14]  ( .CLK(n375), .D(M[14]), .Q(M_reg[14]) );
  LATCHX1 \M_reg_reg[13]  ( .CLK(n375), .D(M[13]), .Q(M_reg[13]) );
  LATCHX1 \M_reg_reg[12]  ( .CLK(n375), .D(M[12]), .Q(M_reg[12]) );
  LATCHX1 \M_reg_reg[11]  ( .CLK(n375), .D(M[11]), .Q(M_reg[11]) );
  LATCHX1 \M_reg_reg[10]  ( .CLK(n375), .D(M[10]), .Q(M_reg[10]) );
  LATCHX1 \M_reg_reg[9]  ( .CLK(n374), .D(M[9]), .Q(M_reg[9]) );
  LATCHX1 \M_reg_reg[8]  ( .CLK(n375), .D(M[8]), .Q(M_reg[8]) );
  LATCHX1 \M_reg_reg[7]  ( .CLK(n374), .D(M[7]), .Q(M_reg[7]) );
  LATCHX1 \M_reg_reg[6]  ( .CLK(n374), .D(M[6]), .Q(M_reg[6]) );
  LATCHX1 \M_reg_reg[5]  ( .CLK(n374), .D(M[5]), .Q(M_reg[5]) );
  LATCHX1 \M_reg_reg[4]  ( .CLK(n374), .D(M[4]), .Q(M_reg[4]) );
  LATCHX1 \M_reg_reg[3]  ( .CLK(n374), .D(M[3]), .Q(M_reg[3]) );
  LATCHX1 \M_reg_reg[2]  ( .CLK(n374), .D(M[2]), .Q(M_reg[2]) );
  LATCHX1 \M_reg_reg[1]  ( .CLK(n374), .D(M[1]), .Q(M_reg[1]) );
  LATCHX1 \M_reg_reg[0]  ( .CLK(n374), .D(M[0]), .Q(M_reg[0]) );
  DFFARX1 \P_reg[63]  ( .D(Acc[31]), .CLK(oClk), .RSTB(n359), .Q(P[63]) );
  DFFARX1 \P_reg[62]  ( .D(Acc[31]), .CLK(oClk), .RSTB(n359), .Q(P[62]) );
  DFFARX1 \P_reg[61]  ( .D(Acc[30]), .CLK(oClk), .RSTB(n359), .Q(P[61]) );
  DFFARX1 \P_reg[60]  ( .D(Acc[29]), .CLK(oClk), .RSTB(n359), .Q(P[60]) );
  DFFARX1 \P_reg[59]  ( .D(Acc[28]), .CLK(oClk), .RSTB(n358), .Q(P[59]) );
  DFFARX1 \P_reg[58]  ( .D(Acc[27]), .CLK(oClk), .RSTB(n358), .Q(P[58]) );
  DFFARX1 \P_reg[57]  ( .D(Acc[26]), .CLK(oClk), .RSTB(n358), .Q(P[57]) );
  DFFARX1 \P_reg[56]  ( .D(Acc[25]), .CLK(oClk), .RSTB(n358), .Q(P[56]) );
  DFFARX1 \P_reg[55]  ( .D(Acc[24]), .CLK(oClk), .RSTB(n358), .Q(P[55]) );
  DFFARX1 \P_reg[54]  ( .D(Acc[23]), .CLK(oClk), .RSTB(n357), .Q(P[54]) );
  DFFARX1 \P_reg[53]  ( .D(Acc[22]), .CLK(oClk), .RSTB(n357), .Q(P[53]) );
  DFFARX1 \P_reg[52]  ( .D(Acc[21]), .CLK(oClk), .RSTB(n357), .Q(P[52]) );
  DFFARX1 \P_reg[51]  ( .D(Acc[20]), .CLK(oClk), .RSTB(n357), .Q(P[51]) );
  DFFARX1 \P_reg[50]  ( .D(n394), .CLK(oClk), .RSTB(n357), .Q(P[50]) );
  DFFARX1 \P_reg[49]  ( .D(Acc[18]), .CLK(oClk), .RSTB(n356), .Q(P[49]) );
  DFFARX1 \P_reg[48]  ( .D(Acc[17]), .CLK(oClk), .RSTB(n356), .Q(P[48]) );
  DFFARX1 \P_reg[47]  ( .D(Acc[16]), .CLK(oClk), .RSTB(n356), .Q(P[47]) );
  DFFARX1 \P_reg[46]  ( .D(Acc[15]), .CLK(oClk), .RSTB(n356), .Q(P[46]) );
  DFFARX1 \P_reg[45]  ( .D(n402), .CLK(oClk), .RSTB(n356), .Q(P[45]) );
  DFFARX1 \P_reg[44]  ( .D(n333), .CLK(oClk), .RSTB(n355), .Q(P[44]) );
  DFFARX1 \P_reg[43]  ( .D(n336), .CLK(oClk), .RSTB(n355), .Q(P[43]) );
  DFFARX1 \P_reg[42]  ( .D(n332), .CLK(oClk), .RSTB(n355), .Q(P[42]) );
  DFFARX1 \P_reg[41]  ( .D(n407), .CLK(oClk), .RSTB(n355), .Q(P[41]) );
  DFFARX1 \P_reg[40]  ( .D(n320), .CLK(oClk), .RSTB(n355), .Q(P[40]) );
  DFFARX1 \P_reg[39]  ( .D(Acc[8]), .CLK(oClk), .RSTB(n354), .Q(P[39]) );
  DFFARX1 \P_reg[38]  ( .D(Acc[7]), .CLK(oClk), .RSTB(n354), .Q(P[38]) );
  DFFARX1 \P_reg[37]  ( .D(Acc[6]), .CLK(oClk), .RSTB(n354), .Q(P[37]) );
  DFFARX1 \P_reg[36]  ( .D(Acc[5]), .CLK(oClk), .RSTB(n354), .Q(P[36]) );
  DFFARX1 \P_reg[35]  ( .D(Acc[4]), .CLK(oClk), .RSTB(n354), .Q(P[35]) );
  DFFARX1 \P_reg[34]  ( .D(n330), .CLK(oClk), .RSTB(n353), .Q(P[34]) );
  DFFARX1 \P_reg[33]  ( .D(n419), .CLK(oClk), .RSTB(n353), .Q(P[33]) );
  DFFARX1 \P_reg[32]  ( .D(n335), .CLK(oClk), .RSTB(n353), .Q(P[32]) );
  DFFARX1 \P_reg[31]  ( .D(Acc[0]), .CLK(oClk), .RSTB(n353), .Q(P[31]) );
  DFFARX1 \P_reg[30]  ( .D(Q_reg[31]), .CLK(oClk), .RSTB(n353), .Q(P[30]) );
  DFFARX1 \P_reg[29]  ( .D(Q_reg[30]), .CLK(oClk), .RSTB(n352), .Q(P[29]) );
  DFFARX1 \P_reg[28]  ( .D(Q_reg[29]), .CLK(oClk), .RSTB(n352), .Q(P[28]) );
  DFFARX1 \P_reg[27]  ( .D(Q_reg[28]), .CLK(oClk), .RSTB(n352), .Q(P[27]) );
  DFFARX1 \P_reg[26]  ( .D(Q_reg[27]), .CLK(oClk), .RSTB(n352), .Q(P[26]) );
  DFFARX1 \P_reg[25]  ( .D(Q_reg[26]), .CLK(oClk), .RSTB(n352), .Q(P[25]) );
  DFFARX1 \P_reg[24]  ( .D(Q_reg[25]), .CLK(oClk), .RSTB(n351), .Q(P[24]) );
  DFFARX1 \P_reg[23]  ( .D(Q_reg[24]), .CLK(oClk), .RSTB(n351), .Q(P[23]) );
  DFFARX1 \P_reg[22]  ( .D(Q_reg[23]), .CLK(oClk), .RSTB(n351), .Q(P[22]) );
  DFFARX1 \P_reg[21]  ( .D(Q_reg[22]), .CLK(oClk), .RSTB(n351), .Q(P[21]) );
  DFFARX1 \P_reg[20]  ( .D(Q_reg[21]), .CLK(oClk), .RSTB(n351), .Q(P[20]) );
  DFFARX1 \P_reg[19]  ( .D(Q_reg[20]), .CLK(oClk), .RSTB(n350), .Q(P[19]) );
  DFFARX1 \P_reg[18]  ( .D(Q_reg[19]), .CLK(oClk), .RSTB(n350), .Q(P[18]) );
  DFFARX1 \P_reg[17]  ( .D(Q_reg[18]), .CLK(oClk), .RSTB(n350), .Q(P[17]) );
  DFFARX1 \P_reg[16]  ( .D(Q_reg[17]), .CLK(oClk), .RSTB(n350), .Q(P[16]) );
  DFFARX1 \P_reg[15]  ( .D(Q_reg[16]), .CLK(oClk), .RSTB(n350), .Q(P[15]) );
  DFFARX1 \P_reg[14]  ( .D(Q_reg[15]), .CLK(oClk), .RSTB(n349), .Q(P[14]) );
  DFFARX1 \P_reg[13]  ( .D(Q_reg[14]), .CLK(oClk), .RSTB(n349), .Q(P[13]) );
  DFFARX1 \P_reg[12]  ( .D(Q_reg[13]), .CLK(oClk), .RSTB(n349), .Q(P[12]) );
  DFFARX1 \P_reg[11]  ( .D(Q_reg[12]), .CLK(oClk), .RSTB(n349), .Q(P[11]) );
  DFFARX1 \P_reg[10]  ( .D(Q_reg[11]), .CLK(oClk), .RSTB(n349), .Q(P[10]) );
  DFFARX1 \P_reg[9]  ( .D(Q_reg[10]), .CLK(oClk), .RSTB(n348), .Q(P[9]) );
  DFFARX1 \P_reg[8]  ( .D(Q_reg[9]), .CLK(oClk), .RSTB(n348), .Q(P[8]) );
  DFFARX1 \P_reg[7]  ( .D(Q_reg[8]), .CLK(oClk), .RSTB(n348), .Q(P[7]) );
  DFFARX1 \P_reg[6]  ( .D(Q_reg[7]), .CLK(oClk), .RSTB(n348), .Q(P[6]) );
  DFFARX1 \P_reg[5]  ( .D(Q_reg[6]), .CLK(oClk), .RSTB(n348), .Q(P[5]) );
  DFFARX1 \P_reg[4]  ( .D(Q_reg[5]), .CLK(oClk), .RSTB(n347), .Q(P[4]) );
  DFFARX1 \P_reg[3]  ( .D(Q_reg[4]), .CLK(oClk), .RSTB(n347), .Q(P[3]) );
  DFFARX1 \P_reg[2]  ( .D(Q_reg[3]), .CLK(oClk), .RSTB(n347), .Q(P[2]) );
  DFFARX1 \P_reg[1]  ( .D(Q_reg[2]), .CLK(oClk), .RSTB(n347), .Q(P[1]) );
  DFFARX1 \P_reg[0]  ( .D(Q_reg[1]), .CLK(oClk), .RSTB(n347), .Q(P[0]) );
  DFFASX1 \count_reg[0]  ( .D(n310), .CLK(clk), .SETB(n376), .Q(count[0]), 
        .QN(n312) );
  DFFARX1 \count_reg[5]  ( .D(n309), .CLK(clk), .RSTB(n377), .Q(count[5]), 
        .QN(n317) );
  DFFASX1 \count_reg[1]  ( .D(n308), .CLK(clk), .SETB(n378), .Q(count[1]), 
        .QN(n315) );
  DFFASX1 \count_reg[2]  ( .D(n307), .CLK(clk), .SETB(n379), .Q(count[2]) );
  DFFASX1 \count_reg[3]  ( .D(n306), .CLK(clk), .SETB(n377), .Q(count[3]) );
  DFFASX1 \count_reg[4]  ( .D(n305), .CLK(clk), .SETB(n376), .Q(count[4]) );
  DFFASRX1 \Q_reg_reg[0]  ( .D(n304), .CLK(clk), .RSTB(n238), .SETB(n237), .Q(
        n314), .QN(n173) );
  DFFARX1 Q_prev_reg ( .D(n303), .CLK(clk), .RSTB(n376), .Q(n172), .QN(n318)
         );
  DFFARX1 \Acc_reg[31]  ( .D(n302), .CLK(clk), .RSTB(n378), .Q(Acc[31]), .QN(
        n171) );
  DFFARX1 \Acc_reg[30]  ( .D(n301), .CLK(clk), .RSTB(n376), .Q(Acc[30]) );
  DFFARX1 \Acc_reg[29]  ( .D(n300), .CLK(clk), .RSTB(n376), .Q(Acc[29]) );
  DFFARX1 \Acc_reg[28]  ( .D(n299), .CLK(clk), .RSTB(n376), .Q(Acc[28]) );
  DFFARX1 \Acc_reg[27]  ( .D(n298), .CLK(clk), .RSTB(n376), .Q(Acc[27]) );
  DFFARX1 \Acc_reg[26]  ( .D(n297), .CLK(clk), .RSTB(n376), .Q(Acc[26]) );
  DFFARX1 \Acc_reg[25]  ( .D(n296), .CLK(clk), .RSTB(n376), .Q(Acc[25]), .QN(
        n165) );
  DFFARX1 \Acc_reg[24]  ( .D(n295), .CLK(clk), .RSTB(n376), .Q(Acc[24]), .QN(
        n164) );
  DFFARX1 \Acc_reg[23]  ( .D(n294), .CLK(clk), .RSTB(n376), .Q(Acc[23]) );
  DFFARX1 \Acc_reg[22]  ( .D(n293), .CLK(clk), .RSTB(n376), .Q(Acc[22]) );
  DFFARX1 \Acc_reg[21]  ( .D(n292), .CLK(clk), .RSTB(n376), .Q(Acc[21]) );
  DFFARX1 \Acc_reg[20]  ( .D(n291), .CLK(clk), .RSTB(n376), .Q(Acc[20]), .QN(
        n160) );
  DFFARX1 \Acc_reg[19]  ( .D(n290), .CLK(clk), .RSTB(n377), .Q(Acc[19]), .QN(
        n159) );
  DFFARX1 \Acc_reg[18]  ( .D(n289), .CLK(clk), .RSTB(n377), .Q(Acc[18]) );
  DFFARX1 \Acc_reg[17]  ( .D(n288), .CLK(clk), .RSTB(n377), .Q(Acc[17]), .QN(
        n157) );
  DFFARX1 \Acc_reg[16]  ( .D(n287), .CLK(clk), .RSTB(n377), .Q(Acc[16]), .QN(
        n156) );
  DFFARX1 \Acc_reg[15]  ( .D(n286), .CLK(clk), .RSTB(n377), .Q(Acc[15]), .QN(
        n155) );
  DFFARX1 \Acc_reg[14]  ( .D(n285), .CLK(clk), .RSTB(n377), .Q(Acc[14]), .QN(
        n154) );
  DFFARX1 \Acc_reg[13]  ( .D(n284), .CLK(clk), .RSTB(n377), .Q(Acc[13]), .QN(
        n153) );
  DFFARX1 \Acc_reg[12]  ( .D(n283), .CLK(clk), .RSTB(n377), .Q(Acc[12]), .QN(
        n152) );
  DFFARX1 \Acc_reg[11]  ( .D(n282), .CLK(clk), .RSTB(n377), .Q(Acc[11]), .QN(
        n151) );
  DFFARX1 \Acc_reg[10]  ( .D(n281), .CLK(clk), .RSTB(n377), .Q(Acc[10]), .QN(
        n150) );
  DFFARX1 \Acc_reg[9]  ( .D(n280), .CLK(clk), .RSTB(n377), .Q(Acc[9]), .QN(
        n149) );
  DFFARX1 \Acc_reg[8]  ( .D(n279), .CLK(clk), .RSTB(n378), .Q(Acc[8]), .QN(
        n148) );
  DFFARX1 \Acc_reg[7]  ( .D(n278), .CLK(clk), .RSTB(n378), .Q(Acc[7]), .QN(
        n147) );
  DFFARX1 \Acc_reg[6]  ( .D(n277), .CLK(clk), .RSTB(n378), .Q(Acc[6]), .QN(
        n146) );
  DFFARX1 \Acc_reg[5]  ( .D(n276), .CLK(clk), .RSTB(n378), .Q(Acc[5]), .QN(
        n145) );
  DFFARX1 \Acc_reg[4]  ( .D(n275), .CLK(clk), .RSTB(n378), .Q(Acc[4]) );
  DFFARX1 \Acc_reg[3]  ( .D(n274), .CLK(clk), .RSTB(n378), .Q(Acc[3]), .QN(
        n143) );
  DFFARX1 \Acc_reg[2]  ( .D(n273), .CLK(clk), .RSTB(n378), .Q(Acc[2]), .QN(
        n142) );
  DFFARX1 \Acc_reg[1]  ( .D(n272), .CLK(clk), .RSTB(n378), .Q(Acc[1]), .QN(
        n141) );
  DFFARX1 \Acc_reg[0]  ( .D(n271), .CLK(clk), .RSTB(n378), .Q(Acc[0]), .QN(
        n140) );
  DFFASRX1 \Q_reg_reg[31]  ( .D(n270), .CLK(clk), .RSTB(n236), .SETB(n235), 
        .Q(Q_reg[31]) );
  DFFASRX1 \Q_reg_reg[30]  ( .D(n269), .CLK(clk), .RSTB(n234), .SETB(n233), 
        .Q(Q_reg[30]) );
  DFFASRX1 \Q_reg_reg[29]  ( .D(n268), .CLK(clk), .RSTB(n232), .SETB(n231), 
        .Q(Q_reg[29]) );
  DFFASRX1 \Q_reg_reg[28]  ( .D(n267), .CLK(clk), .RSTB(n230), .SETB(n229), 
        .Q(Q_reg[28]) );
  DFFASRX1 \Q_reg_reg[27]  ( .D(n266), .CLK(clk), .RSTB(n228), .SETB(n227), 
        .Q(Q_reg[27]) );
  DFFASRX1 \Q_reg_reg[26]  ( .D(n265), .CLK(clk), .RSTB(n226), .SETB(n225), 
        .Q(Q_reg[26]) );
  DFFASRX1 \Q_reg_reg[25]  ( .D(n264), .CLK(clk), .RSTB(n224), .SETB(n223), 
        .Q(Q_reg[25]) );
  DFFASRX1 \Q_reg_reg[24]  ( .D(n263), .CLK(clk), .RSTB(n222), .SETB(n221), 
        .Q(Q_reg[24]) );
  DFFASRX1 \Q_reg_reg[23]  ( .D(n262), .CLK(clk), .RSTB(n220), .SETB(n219), 
        .Q(Q_reg[23]) );
  DFFASRX1 \Q_reg_reg[22]  ( .D(n261), .CLK(clk), .RSTB(n218), .SETB(n217), 
        .Q(Q_reg[22]) );
  DFFASRX1 \Q_reg_reg[21]  ( .D(n260), .CLK(clk), .RSTB(n216), .SETB(n215), 
        .Q(Q_reg[21]) );
  DFFASRX1 \Q_reg_reg[20]  ( .D(n259), .CLK(clk), .RSTB(n214), .SETB(n213), 
        .Q(Q_reg[20]) );
  DFFASRX1 \Q_reg_reg[19]  ( .D(n258), .CLK(clk), .RSTB(n212), .SETB(n211), 
        .Q(Q_reg[19]) );
  DFFASRX1 \Q_reg_reg[18]  ( .D(n257), .CLK(clk), .RSTB(n210), .SETB(n209), 
        .Q(Q_reg[18]) );
  DFFASRX1 \Q_reg_reg[17]  ( .D(n256), .CLK(clk), .RSTB(n208), .SETB(n207), 
        .Q(Q_reg[17]) );
  DFFASRX1 \Q_reg_reg[16]  ( .D(n255), .CLK(clk), .RSTB(n206), .SETB(n205), 
        .Q(Q_reg[16]) );
  DFFASRX1 \Q_reg_reg[15]  ( .D(n254), .CLK(clk), .RSTB(n204), .SETB(n203), 
        .Q(Q_reg[15]) );
  DFFASRX1 \Q_reg_reg[14]  ( .D(n253), .CLK(clk), .RSTB(n202), .SETB(n201), 
        .Q(Q_reg[14]) );
  DFFASRX1 \Q_reg_reg[13]  ( .D(n252), .CLK(clk), .RSTB(n200), .SETB(n199), 
        .Q(Q_reg[13]) );
  DFFASRX1 \Q_reg_reg[12]  ( .D(n251), .CLK(clk), .RSTB(n198), .SETB(n197), 
        .Q(Q_reg[12]) );
  DFFASRX1 \Q_reg_reg[11]  ( .D(n250), .CLK(clk), .RSTB(n196), .SETB(n195), 
        .Q(Q_reg[11]) );
  DFFASRX1 \Q_reg_reg[10]  ( .D(n249), .CLK(clk), .RSTB(n194), .SETB(n193), 
        .Q(Q_reg[10]) );
  DFFASRX1 \Q_reg_reg[9]  ( .D(n248), .CLK(clk), .RSTB(n192), .SETB(n191), .Q(
        Q_reg[9]) );
  DFFASRX1 \Q_reg_reg[8]  ( .D(n247), .CLK(clk), .RSTB(n190), .SETB(n189), .Q(
        Q_reg[8]) );
  DFFASRX1 \Q_reg_reg[7]  ( .D(n246), .CLK(clk), .RSTB(n188), .SETB(n187), .Q(
        Q_reg[7]) );
  DFFASRX1 \Q_reg_reg[6]  ( .D(n245), .CLK(clk), .RSTB(n186), .SETB(n185), .Q(
        Q_reg[6]) );
  DFFASRX1 \Q_reg_reg[5]  ( .D(n244), .CLK(clk), .RSTB(n184), .SETB(n183), .Q(
        Q_reg[5]) );
  DFFASRX1 \Q_reg_reg[4]  ( .D(n243), .CLK(clk), .RSTB(n182), .SETB(n181), .Q(
        Q_reg[4]) );
  DFFASRX1 \Q_reg_reg[3]  ( .D(n242), .CLK(clk), .RSTB(n180), .SETB(n179), .Q(
        Q_reg[3]) );
  DFFASRX1 \Q_reg_reg[2]  ( .D(n241), .CLK(clk), .RSTB(n178), .SETB(n177), .Q(
        Q_reg[2]) );
  DFFASRX1 \Q_reg_reg[1]  ( .D(n240), .CLK(clk), .RSTB(n176), .SETB(n175), .Q(
        Q_reg[1]) );
  AO22X1 U4 ( .IN1(N47), .IN2(n365), .IN3(n361), .IN4(count[5]), .Q(n309) );
  AO22X1 U5 ( .IN1(N46), .IN2(n365), .IN3(n361), .IN4(count[4]), .Q(n305) );
  AO22X1 U9 ( .IN1(N45), .IN2(n365), .IN3(n361), .IN4(count[3]), .Q(n306) );
  AO22X1 U13 ( .IN1(n365), .IN2(Q_reg[10]), .IN3(n361), .IN4(Q_reg[9]), .Q(
        n248) );
  OR2X1 U15 ( .IN1(n379), .IN2(Q[9]), .Q(n192) );
  AO22X1 U16 ( .IN1(n371), .IN2(Q_reg[9]), .IN3(n361), .IN4(Q_reg[8]), .Q(n247) );
  OR2X1 U19 ( .IN1(n379), .IN2(Q[8]), .Q(n190) );
  AO22X1 U20 ( .IN1(n371), .IN2(Q_reg[8]), .IN3(n361), .IN4(Q_reg[7]), .Q(n246) );
  OR2X1 U23 ( .IN1(n379), .IN2(Q[7]), .Q(n188) );
  AO22X1 U24 ( .IN1(n371), .IN2(Q_reg[7]), .IN3(n361), .IN4(Q_reg[6]), .Q(n245) );
  OR2X1 U27 ( .IN1(n379), .IN2(Q[6]), .Q(n186) );
  AO22X1 U28 ( .IN1(n370), .IN2(Q_reg[6]), .IN3(n361), .IN4(Q_reg[5]), .Q(n244) );
  OR2X1 U31 ( .IN1(n379), .IN2(Q[5]), .Q(n184) );
  AO22X1 U32 ( .IN1(n370), .IN2(Q_reg[5]), .IN3(n361), .IN4(Q_reg[4]), .Q(n243) );
  OR2X1 U35 ( .IN1(n378), .IN2(Q[4]), .Q(n182) );
  AO22X1 U36 ( .IN1(n370), .IN2(Q_reg[4]), .IN3(n361), .IN4(Q_reg[3]), .Q(n242) );
  OR2X1 U39 ( .IN1(n378), .IN2(Q[3]), .Q(n180) );
  OR2X1 U43 ( .IN1(n378), .IN2(Q[31]), .Q(n236) );
  AO22X1 U44 ( .IN1(n370), .IN2(Q_reg[31]), .IN3(n361), .IN4(Q_reg[30]), .Q(
        n269) );
  OR2X1 U47 ( .IN1(n379), .IN2(Q[30]), .Q(n234) );
  AO22X1 U48 ( .IN1(n370), .IN2(Q_reg[3]), .IN3(n361), .IN4(Q_reg[2]), .Q(n241) );
  OR2X1 U51 ( .IN1(n379), .IN2(Q[2]), .Q(n178) );
  AO22X1 U52 ( .IN1(n369), .IN2(Q_reg[30]), .IN3(n361), .IN4(Q_reg[29]), .Q(
        n268) );
  OR2X1 U55 ( .IN1(n379), .IN2(Q[29]), .Q(n232) );
  AO22X1 U56 ( .IN1(n369), .IN2(Q_reg[29]), .IN3(n361), .IN4(Q_reg[28]), .Q(
        n267) );
  OR2X1 U59 ( .IN1(n379), .IN2(Q[28]), .Q(n230) );
  AO22X1 U60 ( .IN1(n369), .IN2(Q_reg[28]), .IN3(n361), .IN4(Q_reg[27]), .Q(
        n266) );
  OR2X1 U63 ( .IN1(n379), .IN2(Q[27]), .Q(n228) );
  AO22X1 U64 ( .IN1(n369), .IN2(Q_reg[27]), .IN3(n360), .IN4(Q_reg[26]), .Q(
        n265) );
  OR2X1 U67 ( .IN1(n379), .IN2(Q[26]), .Q(n226) );
  AO22X1 U68 ( .IN1(n369), .IN2(Q_reg[26]), .IN3(n360), .IN4(Q_reg[25]), .Q(
        n264) );
  OR2X1 U71 ( .IN1(n379), .IN2(Q[25]), .Q(n224) );
  AO22X1 U72 ( .IN1(n368), .IN2(Q_reg[25]), .IN3(n360), .IN4(Q_reg[24]), .Q(
        n263) );
  OR2X1 U75 ( .IN1(n379), .IN2(Q[24]), .Q(n222) );
  AO22X1 U76 ( .IN1(n368), .IN2(Q_reg[24]), .IN3(n360), .IN4(Q_reg[23]), .Q(
        n262) );
  OR2X1 U79 ( .IN1(n379), .IN2(Q[23]), .Q(n220) );
  AO22X1 U80 ( .IN1(n368), .IN2(Q_reg[23]), .IN3(n360), .IN4(Q_reg[22]), .Q(
        n261) );
  OR2X1 U83 ( .IN1(n379), .IN2(Q[22]), .Q(n218) );
  AO22X1 U84 ( .IN1(n368), .IN2(Q_reg[22]), .IN3(n360), .IN4(Q_reg[21]), .Q(
        n260) );
  OR2X1 U87 ( .IN1(n379), .IN2(Q[21]), .Q(n216) );
  AO22X1 U88 ( .IN1(n367), .IN2(Q_reg[21]), .IN3(n360), .IN4(Q_reg[20]), .Q(
        n259) );
  OR2X1 U91 ( .IN1(n379), .IN2(Q[20]), .Q(n214) );
  AO22X1 U92 ( .IN1(n367), .IN2(Q_reg[2]), .IN3(n360), .IN4(Q_reg[1]), .Q(n240) );
  OR2X1 U95 ( .IN1(n377), .IN2(Q[1]), .Q(n176) );
  AO22X1 U96 ( .IN1(n367), .IN2(Q_reg[20]), .IN3(n360), .IN4(Q_reg[19]), .Q(
        n258) );
  OR2X1 U99 ( .IN1(n376), .IN2(Q[19]), .Q(n212) );
  AO22X1 U100 ( .IN1(n367), .IN2(Q_reg[19]), .IN3(n360), .IN4(Q_reg[18]), .Q(
        n257) );
  OR2X1 U103 ( .IN1(n378), .IN2(Q[18]), .Q(n210) );
  AO22X1 U104 ( .IN1(n367), .IN2(Q_reg[18]), .IN3(n360), .IN4(Q_reg[17]), .Q(
        n256) );
  OR2X1 U107 ( .IN1(n379), .IN2(Q[17]), .Q(n208) );
  AO22X1 U108 ( .IN1(n366), .IN2(Q_reg[17]), .IN3(n360), .IN4(Q_reg[16]), .Q(
        n255) );
  OR2X1 U111 ( .IN1(n377), .IN2(Q[16]), .Q(n206) );
  AO22X1 U112 ( .IN1(n366), .IN2(Q_reg[16]), .IN3(n360), .IN4(Q_reg[15]), .Q(
        n254) );
  OR2X1 U115 ( .IN1(n379), .IN2(Q[15]), .Q(n204) );
  AO22X1 U116 ( .IN1(n366), .IN2(Q_reg[15]), .IN3(n360), .IN4(Q_reg[14]), .Q(
        n253) );
  OR2X1 U119 ( .IN1(n378), .IN2(Q[14]), .Q(n202) );
  AO22X1 U120 ( .IN1(n366), .IN2(Q_reg[14]), .IN3(n360), .IN4(Q_reg[13]), .Q(
        n252) );
  OR2X1 U123 ( .IN1(n378), .IN2(Q[13]), .Q(n200) );
  AO22X1 U124 ( .IN1(n366), .IN2(Q_reg[13]), .IN3(n360), .IN4(Q_reg[12]), .Q(
        n251) );
  OR2X1 U127 ( .IN1(n379), .IN2(Q[12]), .Q(n198) );
  AO22X1 U128 ( .IN1(n365), .IN2(Q_reg[12]), .IN3(n360), .IN4(Q_reg[11]), .Q(
        n250) );
  OR2X1 U131 ( .IN1(n377), .IN2(Q[11]), .Q(n196) );
  AO22X1 U132 ( .IN1(n368), .IN2(Q_reg[11]), .IN3(n360), .IN4(Q_reg[10]), .Q(
        n249) );
  OR2X1 U136 ( .IN1(n376), .IN2(Q[10]), .Q(n194) );
  OR2X1 U140 ( .IN1(n376), .IN2(Q[0]), .Q(n238) );
  BoothMultiplier_DW01_sub_1 sub_61 ( .A({Acc[31:20], n394, Acc[18:15], n402, 
        n333, n336, n332, Acc[10], n320, Acc[8:4], n330, Acc[2], n335, Acc[0]}), .B(M_reg), .CI(1'b0), .DIFF(case_sub) );
  BoothMultiplier_DW01_add_1 add_57 ( .A({Acc[31:21], n392, Acc[19:18], n397, 
        n399, n334, Acc[14:11], n337, Acc[9:7], n329, Acc[5:3], n331, Acc[1:0]}), .B(M_reg), .CI(1'b0), .SUM(case_add) );
  INVX0 U246 ( .INP(n423), .ZN(n381) );
  OR2X1 U247 ( .IN1(n422), .IN2(n326), .Q(n302) );
  AOI22X1 U248 ( .IN1(n362), .IN2(Acc[26]), .IN3(n338), .IN4(Acc[27]), .QN(
        n313) );
  AOI22X1 U249 ( .IN1(n362), .IN2(Acc[27]), .IN3(n338), .IN4(Acc[28]), .QN(
        n316) );
  INVX0 U250 ( .INP(Acc[2]), .ZN(n319) );
  INVX0 U251 ( .INP(n149), .ZN(n320) );
  INVX0 U252 ( .INP(n150), .ZN(n337) );
  NAND2X0 U253 ( .IN1(n344), .IN2(case_add[61]), .QN(n321) );
  NAND2X1 U254 ( .IN1(case_sub[61]), .IN2(n343), .QN(n322) );
  NAND3X0 U255 ( .IN1(n321), .IN2(n322), .IN3(n316), .QN(n298) );
  NBUFFX2 U256 ( .INP(n327), .Z(n344) );
  NAND2X0 U257 ( .IN1(case_add[60]), .IN2(n344), .QN(n323) );
  NAND2X1 U258 ( .IN1(case_sub[60]), .IN2(n343), .QN(n324) );
  NAND3X0 U259 ( .IN1(n323), .IN2(n324), .IN3(n313), .QN(n297) );
  INVX0 U260 ( .INP(n364), .ZN(n360) );
  INVX0 U261 ( .INP(n364), .ZN(n361) );
  INVX0 U262 ( .INP(n364), .ZN(n362) );
  NBUFFX2 U263 ( .INP(n325), .Z(n340) );
  NBUFFX2 U264 ( .INP(n328), .Z(n343) );
  NBUFFX2 U265 ( .INP(N4), .Z(n364) );
  NBUFFX2 U266 ( .INP(n327), .Z(n346) );
  NBUFFX2 U267 ( .INP(N4), .Z(n363) );
  AND2X1 U268 ( .IN1(n381), .IN2(n363), .Q(n325) );
  NBUFFX2 U269 ( .INP(N4), .Z(n365) );
  NBUFFX2 U270 ( .INP(N4), .Z(n366) );
  NBUFFX2 U271 ( .INP(N4), .Z(n367) );
  NBUFFX2 U272 ( .INP(N4), .Z(n368) );
  NBUFFX2 U273 ( .INP(N4), .Z(n369) );
  NBUFFX2 U274 ( .INP(N4), .Z(n370) );
  NBUFFX2 U275 ( .INP(N4), .Z(n371) );
  INVX0 U276 ( .INP(n428), .ZN(n432) );
  INVX0 U277 ( .INP(n426), .ZN(n430) );
  INVX0 U278 ( .INP(n427), .ZN(n431) );
  NBUFFX2 U279 ( .INP(n433), .Z(n347) );
  NBUFFX2 U280 ( .INP(n433), .Z(n348) );
  NBUFFX2 U281 ( .INP(n433), .Z(n349) );
  NBUFFX2 U282 ( .INP(n433), .Z(n350) );
  NBUFFX2 U283 ( .INP(n433), .Z(n351) );
  NBUFFX2 U284 ( .INP(n433), .Z(n352) );
  NBUFFX2 U285 ( .INP(n433), .Z(n353) );
  NBUFFX2 U286 ( .INP(n433), .Z(n354) );
  NBUFFX2 U287 ( .INP(n433), .Z(n355) );
  NBUFFX2 U288 ( .INP(n433), .Z(n356) );
  NBUFFX2 U289 ( .INP(n433), .Z(n357) );
  NBUFFX2 U290 ( .INP(n433), .Z(n358) );
  NBUFFX2 U291 ( .INP(n433), .Z(n359) );
  AOI21X1 U292 ( .IN1(n423), .IN2(n363), .IN3(n171), .QN(n326) );
  AND3X1 U293 ( .IN1(n172), .IN2(n173), .IN3(n363), .Q(n327) );
  NOR2X0 U294 ( .IN1(count[0]), .IN2(n360), .QN(n310) );
  AND3X1 U295 ( .IN1(n363), .IN2(n314), .IN3(n318), .Q(n328) );
  NOR3X0 U296 ( .IN1(count[2]), .IN2(count[3]), .IN3(count[4]), .QN(n380) );
  INVX0 U297 ( .INP(n157), .ZN(n397) );
  INVX0 U298 ( .INP(n140), .ZN(n424) );
  INVX0 U299 ( .INP(n145), .ZN(n415) );
  INVX0 U300 ( .INP(n147), .ZN(n412) );
  INVX0 U301 ( .INP(n148), .ZN(n410) );
  INVX0 U302 ( .INP(n154), .ZN(n402) );
  INVX0 U303 ( .INP(n156), .ZN(n399) );
  INVX0 U304 ( .INP(n159), .ZN(n394) );
  INVX0 U305 ( .INP(n160), .ZN(n392) );
  INVX0 U306 ( .INP(n164), .ZN(n387) );
  INVX0 U307 ( .INP(n165), .ZN(n385) );
  INVX0 U308 ( .INP(oRst), .ZN(n433) );
  NBUFFX2 U309 ( .INP(rst), .Z(n374) );
  NBUFFX2 U310 ( .INP(rst), .Z(n373) );
  NBUFFX2 U311 ( .INP(rst), .Z(n372) );
  NBUFFX2 U312 ( .INP(rst), .Z(n375) );
  NAND2X1 U313 ( .IN1(Q[10]), .IN2(n374), .QN(n193) );
  NAND2X1 U314 ( .IN1(Q[11]), .IN2(n374), .QN(n195) );
  NAND2X1 U315 ( .IN1(Q[12]), .IN2(n374), .QN(n197) );
  NAND2X1 U316 ( .IN1(Q[13]), .IN2(n374), .QN(n199) );
  NAND2X1 U317 ( .IN1(Q[14]), .IN2(n374), .QN(n201) );
  NAND2X1 U318 ( .IN1(Q[15]), .IN2(n374), .QN(n203) );
  NAND2X1 U319 ( .IN1(Q[16]), .IN2(n374), .QN(n205) );
  NAND2X1 U320 ( .IN1(Q[0]), .IN2(n374), .QN(n237) );
  NAND2X1 U321 ( .IN1(Q[1]), .IN2(n373), .QN(n175) );
  NAND2X1 U322 ( .IN1(Q[2]), .IN2(n372), .QN(n177) );
  NAND2X1 U323 ( .IN1(Q[3]), .IN2(n372), .QN(n179) );
  NAND2X1 U324 ( .IN1(Q[4]), .IN2(n372), .QN(n181) );
  NAND2X1 U325 ( .IN1(Q[5]), .IN2(n372), .QN(n183) );
  NAND2X1 U326 ( .IN1(Q[6]), .IN2(n372), .QN(n185) );
  NAND2X1 U327 ( .IN1(Q[7]), .IN2(n372), .QN(n187) );
  NAND2X1 U328 ( .IN1(Q[8]), .IN2(n372), .QN(n189) );
  NAND2X1 U329 ( .IN1(Q[9]), .IN2(n372), .QN(n191) );
  NAND2X1 U330 ( .IN1(Q[17]), .IN2(n373), .QN(n207) );
  NAND2X1 U331 ( .IN1(Q[18]), .IN2(n373), .QN(n209) );
  NAND2X1 U332 ( .IN1(Q[19]), .IN2(n373), .QN(n211) );
  NAND2X1 U333 ( .IN1(Q[20]), .IN2(n373), .QN(n213) );
  NAND2X1 U334 ( .IN1(Q[21]), .IN2(n373), .QN(n215) );
  NAND2X1 U335 ( .IN1(Q[22]), .IN2(n373), .QN(n217) );
  NAND2X1 U336 ( .IN1(Q[23]), .IN2(n373), .QN(n219) );
  NAND2X1 U337 ( .IN1(Q[24]), .IN2(n373), .QN(n221) );
  NAND2X1 U338 ( .IN1(Q[25]), .IN2(n373), .QN(n223) );
  NAND2X1 U339 ( .IN1(Q[26]), .IN2(n373), .QN(n225) );
  NAND2X1 U340 ( .IN1(Q[27]), .IN2(n373), .QN(n227) );
  NAND2X1 U341 ( .IN1(Q[28]), .IN2(n372), .QN(n229) );
  NAND2X1 U342 ( .IN1(Q[29]), .IN2(n372), .QN(n231) );
  NAND2X1 U343 ( .IN1(Q[30]), .IN2(n372), .QN(n233) );
  NAND2X1 U344 ( .IN1(Q[31]), .IN2(n372), .QN(n235) );
  INVX0 U345 ( .INP(n319), .ZN(n419) );
  INVX0 U346 ( .INP(n146), .ZN(n329) );
  INVX0 U347 ( .INP(n143), .ZN(n330) );
  INVX0 U348 ( .INP(n142), .ZN(n331) );
  INVX0 U349 ( .INP(n151), .ZN(n332) );
  INVX0 U350 ( .INP(n153), .ZN(n333) );
  INVX0 U351 ( .INP(n155), .ZN(n334) );
  INVX0 U352 ( .INP(n141), .ZN(n335) );
  INVX0 U353 ( .INP(n152), .ZN(n336) );
  INVX0 U354 ( .INP(n150), .ZN(n407) );
  NBUFFX2 U355 ( .INP(n325), .Z(n338) );
  NBUFFX2 U356 ( .INP(n325), .Z(n339) );
  NBUFFX2 U357 ( .INP(n328), .Z(n341) );
  NBUFFX2 U358 ( .INP(n328), .Z(n342) );
  NBUFFX2 U359 ( .INP(n327), .Z(n345) );
  INVX0 U360 ( .INP(n374), .ZN(n376) );
  INVX0 U361 ( .INP(n374), .ZN(n377) );
  INVX0 U362 ( .INP(n374), .ZN(n378) );
  INVX0 U363 ( .INP(n374), .ZN(n379) );
  NAND4X0 U364 ( .IN1(n312), .IN2(n317), .IN3(n315), .IN4(n380), .QN(N4) );
  AND2X1 U365 ( .IN1(N44), .IN2(n364), .Q(n307) );
  AND2X1 U366 ( .IN1(N43), .IN2(n364), .Q(n308) );
  MUX21X1 U367 ( .IN1(Q_reg[1]), .IN2(n314), .S(n360), .Q(n304) );
  MUX21X1 U368 ( .IN1(n314), .IN2(n172), .S(n360), .Q(n303) );
  XOR2X1 U369 ( .IN1(n314), .IN2(n172), .Q(n423) );
  AO22X1 U370 ( .IN1(n343), .IN2(case_sub[64]), .IN3(n344), .IN4(case_add[64]), 
        .Q(n422) );
  AO221X1 U371 ( .IN1(n338), .IN2(Acc[31]), .IN3(n360), .IN4(Acc[30]), .IN5(
        n422), .Q(n301) );
  AO22X1 U372 ( .IN1(n361), .IN2(Acc[29]), .IN3(n338), .IN4(Acc[30]), .Q(n382)
         );
  AO221X1 U373 ( .IN1(case_add[63]), .IN2(n344), .IN3(case_sub[63]), .IN4(n343), .IN5(n382), .Q(n300) );
  AO22X1 U374 ( .IN1(n362), .IN2(Acc[28]), .IN3(n338), .IN4(Acc[29]), .Q(n383)
         );
  AO221X1 U375 ( .IN1(case_add[62]), .IN2(n344), .IN3(case_sub[62]), .IN4(n343), .IN5(n383), .Q(n299) );
  AO22X1 U376 ( .IN1(n362), .IN2(n385), .IN3(n338), .IN4(Acc[26]), .Q(n384) );
  AO221X1 U377 ( .IN1(case_add[59]), .IN2(n344), .IN3(case_sub[59]), .IN4(n343), .IN5(n384), .Q(n296) );
  AO22X1 U378 ( .IN1(n362), .IN2(n387), .IN3(n338), .IN4(n385), .Q(n386) );
  AO221X1 U379 ( .IN1(case_add[58]), .IN2(n344), .IN3(case_sub[58]), .IN4(n343), .IN5(n386), .Q(n295) );
  AO22X1 U380 ( .IN1(n362), .IN2(Acc[23]), .IN3(n338), .IN4(n387), .Q(n388) );
  AO221X1 U381 ( .IN1(case_add[57]), .IN2(n344), .IN3(case_sub[57]), .IN4(n343), .IN5(n388), .Q(n294) );
  AO22X1 U382 ( .IN1(n362), .IN2(Acc[22]), .IN3(n338), .IN4(Acc[23]), .Q(n389)
         );
  AO221X1 U383 ( .IN1(case_add[56]), .IN2(n344), .IN3(case_sub[56]), .IN4(n342), .IN5(n389), .Q(n293) );
  AO22X1 U384 ( .IN1(n362), .IN2(Acc[21]), .IN3(n338), .IN4(Acc[22]), .Q(n390)
         );
  AO221X1 U385 ( .IN1(case_add[55]), .IN2(n344), .IN3(case_sub[55]), .IN4(n342), .IN5(n390), .Q(n292) );
  AO22X1 U386 ( .IN1(n362), .IN2(Acc[20]), .IN3(n338), .IN4(Acc[21]), .Q(n391)
         );
  AO221X1 U387 ( .IN1(case_add[54]), .IN2(n344), .IN3(case_sub[54]), .IN4(n342), .IN5(n391), .Q(n291) );
  AO22X1 U388 ( .IN1(n362), .IN2(n394), .IN3(n338), .IN4(Acc[20]), .Q(n393) );
  AO221X1 U389 ( .IN1(case_add[53]), .IN2(n344), .IN3(case_sub[53]), .IN4(n342), .IN5(n393), .Q(n290) );
  AO22X1 U390 ( .IN1(n362), .IN2(Acc[18]), .IN3(n338), .IN4(n394), .Q(n395) );
  AO221X1 U391 ( .IN1(case_add[52]), .IN2(n344), .IN3(case_sub[52]), .IN4(n342), .IN5(n395), .Q(n289) );
  AO22X1 U392 ( .IN1(n361), .IN2(n397), .IN3(n339), .IN4(Acc[18]), .Q(n396) );
  AO221X1 U393 ( .IN1(case_add[51]), .IN2(n345), .IN3(case_sub[51]), .IN4(n342), .IN5(n396), .Q(n288) );
  AO22X1 U394 ( .IN1(n362), .IN2(n399), .IN3(n339), .IN4(n397), .Q(n398) );
  AO221X1 U395 ( .IN1(case_add[50]), .IN2(n345), .IN3(case_sub[50]), .IN4(n342), .IN5(n398), .Q(n287) );
  AO22X1 U396 ( .IN1(n362), .IN2(Acc[15]), .IN3(n339), .IN4(n399), .Q(n400) );
  AO221X1 U397 ( .IN1(case_add[49]), .IN2(n345), .IN3(case_sub[49]), .IN4(n342), .IN5(n400), .Q(n286) );
  AO22X1 U398 ( .IN1(n362), .IN2(n402), .IN3(n339), .IN4(Acc[15]), .Q(n401) );
  AO221X1 U399 ( .IN1(case_add[48]), .IN2(n345), .IN3(case_sub[48]), .IN4(n342), .IN5(n401), .Q(n285) );
  AO22X1 U400 ( .IN1(n362), .IN2(n333), .IN3(n339), .IN4(n402), .Q(n403) );
  AO221X1 U401 ( .IN1(case_add[47]), .IN2(n345), .IN3(case_sub[47]), .IN4(n342), .IN5(n403), .Q(n284) );
  AO22X1 U402 ( .IN1(n362), .IN2(n336), .IN3(n339), .IN4(n333), .Q(n404) );
  AO221X1 U403 ( .IN1(case_add[46]), .IN2(n345), .IN3(case_sub[46]), .IN4(n342), .IN5(n404), .Q(n283) );
  AO22X1 U404 ( .IN1(n362), .IN2(n332), .IN3(n339), .IN4(n336), .Q(n405) );
  AO221X1 U405 ( .IN1(case_add[45]), .IN2(n345), .IN3(case_sub[45]), .IN4(n342), .IN5(n405), .Q(n282) );
  AO22X1 U406 ( .IN1(n362), .IN2(n407), .IN3(n339), .IN4(n332), .Q(n406) );
  AO221X1 U407 ( .IN1(case_add[44]), .IN2(n345), .IN3(case_sub[44]), .IN4(n341), .IN5(n406), .Q(n281) );
  AO22X1 U408 ( .IN1(n362), .IN2(n320), .IN3(n339), .IN4(n407), .Q(n408) );
  AO221X1 U409 ( .IN1(case_add[43]), .IN2(n345), .IN3(case_sub[43]), .IN4(n341), .IN5(n408), .Q(n280) );
  AO22X1 U410 ( .IN1(n362), .IN2(n410), .IN3(n339), .IN4(n320), .Q(n409) );
  AO221X1 U411 ( .IN1(case_add[42]), .IN2(n345), .IN3(case_sub[42]), .IN4(n341), .IN5(n409), .Q(n279) );
  AO22X1 U412 ( .IN1(n362), .IN2(n412), .IN3(n339), .IN4(n410), .Q(n411) );
  AO221X1 U413 ( .IN1(case_add[41]), .IN2(n345), .IN3(case_sub[41]), .IN4(n341), .IN5(n411), .Q(n278) );
  AO22X1 U414 ( .IN1(n361), .IN2(Acc[6]), .IN3(n339), .IN4(n412), .Q(n413) );
  AO221X1 U415 ( .IN1(case_add[40]), .IN2(n345), .IN3(case_sub[40]), .IN4(n341), .IN5(n413), .Q(n277) );
  AO22X1 U416 ( .IN1(n361), .IN2(n415), .IN3(n339), .IN4(Acc[6]), .Q(n414) );
  AO221X1 U417 ( .IN1(case_add[39]), .IN2(n345), .IN3(case_sub[39]), .IN4(n341), .IN5(n414), .Q(n276) );
  AO22X1 U418 ( .IN1(n361), .IN2(Acc[4]), .IN3(n340), .IN4(n415), .Q(n416) );
  AO221X1 U419 ( .IN1(case_add[38]), .IN2(n346), .IN3(case_sub[38]), .IN4(n341), .IN5(n416), .Q(n275) );
  AO22X1 U420 ( .IN1(n361), .IN2(n330), .IN3(n340), .IN4(Acc[4]), .Q(n417) );
  AO221X1 U421 ( .IN1(case_add[37]), .IN2(n346), .IN3(case_sub[37]), .IN4(n341), .IN5(n417), .Q(n274) );
  AO22X1 U422 ( .IN1(n361), .IN2(n419), .IN3(n340), .IN4(n330), .Q(n418) );
  AO221X1 U423 ( .IN1(case_add[36]), .IN2(n346), .IN3(case_sub[36]), .IN4(n341), .IN5(n418), .Q(n273) );
  AO22X1 U424 ( .IN1(n361), .IN2(n335), .IN3(n340), .IN4(n419), .Q(n420) );
  AO221X1 U425 ( .IN1(case_add[35]), .IN2(n346), .IN3(case_sub[35]), .IN4(n341), .IN5(n420), .Q(n272) );
  AO22X1 U426 ( .IN1(n361), .IN2(n424), .IN3(n340), .IN4(n335), .Q(n421) );
  AO221X1 U427 ( .IN1(case_add[34]), .IN2(n346), .IN3(case_sub[34]), .IN4(n341), .IN5(n421), .Q(n271) );
  AO22X1 U428 ( .IN1(n361), .IN2(Q_reg[31]), .IN3(n340), .IN4(n424), .Q(n425)
         );
  AO221X1 U429 ( .IN1(case_add[33]), .IN2(n346), .IN3(case_sub[33]), .IN4(n341), .IN5(n425), .Q(n270) );
  NOR2X0 U430 ( .IN1(count[1]), .IN2(count[0]), .QN(n426) );
  AO21X1 U431 ( .IN1(count[1]), .IN2(count[0]), .IN3(n426), .Q(N43) );
  NOR2X0 U432 ( .IN1(n430), .IN2(count[2]), .QN(n427) );
  AO21X1 U433 ( .IN1(count[2]), .IN2(n430), .IN3(n427), .Q(N44) );
  NOR2X0 U434 ( .IN1(n431), .IN2(count[3]), .QN(n428) );
  AO21X1 U435 ( .IN1(count[3]), .IN2(n431), .IN3(n428), .Q(N45) );
  XNOR2X1 U436 ( .IN1(count[4]), .IN2(n432), .Q(N46) );
  NOR2X0 U437 ( .IN1(count[4]), .IN2(n432), .QN(n429) );
  XOR2X1 U438 ( .IN1(count[5]), .IN2(n429), .Q(N47) );
endmodule

