
module FP_MULTIPLIER_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[7]), .B(A[7]), .Z(SUM[7]) );
endmodule


module FP_MULTIPLIER_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [46:0] A;
  input [4:0] SH;
  output [46:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][46] , \ML_int[1][45] , \ML_int[1][44] , \ML_int[1][43] ,
         \ML_int[1][42] , \ML_int[1][41] , \ML_int[1][40] , \ML_int[1][39] ,
         \ML_int[1][38] , \ML_int[1][37] , \ML_int[1][36] , \ML_int[1][35] ,
         \ML_int[1][34] , \ML_int[1][33] , \ML_int[1][32] , \ML_int[1][31] ,
         \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] , \ML_int[1][27] ,
         \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] , \ML_int[1][23] ,
         \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] , \ML_int[1][19] ,
         \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] , \ML_int[1][15] ,
         \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] , \ML_int[1][11] ,
         \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] , \ML_int[1][7] ,
         \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] , \ML_int[1][3] ,
         \ML_int[1][2] , \ML_int[1][1] , \ML_int[2][46] , \ML_int[2][45] ,
         \ML_int[2][44] , \ML_int[2][43] , \ML_int[2][42] , \ML_int[2][41] ,
         \ML_int[2][40] , \ML_int[2][39] , \ML_int[2][38] , \ML_int[2][37] ,
         \ML_int[2][36] , \ML_int[2][35] , \ML_int[2][34] , \ML_int[2][33] ,
         \ML_int[2][32] , \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] ,
         \ML_int[2][28] , \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] ,
         \ML_int[2][24] , \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] ,
         \ML_int[2][20] , \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] ,
         \ML_int[2][16] , \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] ,
         \ML_int[2][12] , \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] ,
         \ML_int[2][8] , \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] ,
         \ML_int[2][4] , \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] ,
         \ML_int[2][0] , \ML_int[3][46] , \ML_int[3][45] , \ML_int[3][44] ,
         \ML_int[3][43] , \ML_int[3][42] , \ML_int[3][41] , \ML_int[3][40] ,
         \ML_int[3][39] , \ML_int[3][38] , \ML_int[3][37] , \ML_int[3][36] ,
         \ML_int[3][35] , \ML_int[3][34] , \ML_int[3][33] , \ML_int[3][32] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][46] , \ML_int[4][45] , \ML_int[4][44] , \ML_int[4][43] ,
         \ML_int[4][42] , \ML_int[4][41] , \ML_int[4][40] , \ML_int[4][39] ,
         \ML_int[4][38] , \ML_int[4][37] , \ML_int[4][36] , \ML_int[4][35] ,
         \ML_int[4][34] , \ML_int[4][33] , \ML_int[4][32] , \ML_int[4][31] ,
         \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] , \ML_int[4][27] ,
         \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] , \ML_int[4][23] ,
         \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] , \ML_int[4][19] ,
         \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] , \ML_int[4][15] ,
         \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] , \ML_int[4][11] ,
         \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] , \ML_int[5][46] ,
         \ML_int[5][45] , \ML_int[5][44] , \ML_int[5][43] , \ML_int[5][42] ,
         \ML_int[5][41] , \ML_int[5][40] , \ML_int[5][39] , \ML_int[5][38] ,
         \ML_int[5][37] , \ML_int[5][36] , \ML_int[5][35] , \ML_int[5][34] ,
         \ML_int[5][33] , \ML_int[5][32] , \ML_int[5][31] , \ML_int[5][30] ,
         \ML_int[5][29] , \ML_int[5][28] , \ML_int[5][27] , \ML_int[5][26] ,
         \ML_int[5][25] , \ML_int[5][24] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65;
  assign B[46] = \ML_int[5][46] ;
  assign B[45] = \ML_int[5][45] ;
  assign B[44] = \ML_int[5][44] ;
  assign B[43] = \ML_int[5][43] ;
  assign B[42] = \ML_int[5][42] ;
  assign B[41] = \ML_int[5][41] ;
  assign B[40] = \ML_int[5][40] ;
  assign B[39] = \ML_int[5][39] ;
  assign B[38] = \ML_int[5][38] ;
  assign B[37] = \ML_int[5][37] ;
  assign B[36] = \ML_int[5][36] ;
  assign B[35] = \ML_int[5][35] ;
  assign B[34] = \ML_int[5][34] ;
  assign B[33] = \ML_int[5][33] ;
  assign B[32] = \ML_int[5][32] ;
  assign B[31] = \ML_int[5][31] ;
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;

  MUX2_X1 M1_4_44 ( .A(\ML_int[4][44] ), .B(\ML_int[4][28] ), .S(n60), .Z(
        \ML_int[5][44] ) );
  MUX2_X1 M1_4_43 ( .A(\ML_int[4][43] ), .B(\ML_int[4][27] ), .S(n60), .Z(
        \ML_int[5][43] ) );
  MUX2_X1 M1_4_42 ( .A(\ML_int[4][42] ), .B(\ML_int[4][26] ), .S(n60), .Z(
        \ML_int[5][42] ) );
  MUX2_X1 M1_4_41 ( .A(\ML_int[4][41] ), .B(\ML_int[4][25] ), .S(n60), .Z(
        \ML_int[5][41] ) );
  MUX2_X1 M1_4_40 ( .A(\ML_int[4][40] ), .B(\ML_int[4][24] ), .S(n60), .Z(
        \ML_int[5][40] ) );
  MUX2_X1 M1_4_39 ( .A(\ML_int[4][39] ), .B(\ML_int[4][23] ), .S(n60), .Z(
        \ML_int[5][39] ) );
  MUX2_X1 M1_4_36 ( .A(\ML_int[4][36] ), .B(\ML_int[4][20] ), .S(n60), .Z(
        \ML_int[5][36] ) );
  MUX2_X1 M1_4_35 ( .A(\ML_int[4][35] ), .B(\ML_int[4][19] ), .S(n60), .Z(
        \ML_int[5][35] ) );
  MUX2_X1 M1_4_34 ( .A(\ML_int[4][34] ), .B(\ML_int[4][18] ), .S(n61), .Z(
        \ML_int[5][34] ) );
  MUX2_X1 M1_4_33 ( .A(\ML_int[4][33] ), .B(\ML_int[4][17] ), .S(n61), .Z(
        \ML_int[5][33] ) );
  MUX2_X1 M1_4_32 ( .A(\ML_int[4][32] ), .B(\ML_int[4][16] ), .S(n61), .Z(
        \ML_int[5][32] ) );
  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n61), .Z(
        \ML_int[5][31] ) );
  MUX2_X1 M1_4_30 ( .A(n27), .B(\ML_int[4][14] ), .S(n61), .Z(\ML_int[5][30] )
         );
  MUX2_X1 M1_4_29 ( .A(n28), .B(\ML_int[4][13] ), .S(n61), .Z(\ML_int[5][29] )
         );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n61), .Z(
        \ML_int[5][28] ) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n61), .Z(
        \ML_int[5][27] ) );
  MUX2_X1 M1_4_26 ( .A(n18), .B(\ML_int[4][10] ), .S(n61), .Z(\ML_int[5][26] )
         );
  MUX2_X1 M1_4_25 ( .A(n13), .B(\ML_int[4][9] ), .S(n61), .Z(\ML_int[5][25] )
         );
  MUX2_X1 M1_4_24 ( .A(n19), .B(\ML_int[4][8] ), .S(n61), .Z(\ML_int[5][24] )
         );
  MUX2_X1 M1_3_46 ( .A(\ML_int[3][46] ), .B(\ML_int[3][38] ), .S(n59), .Z(
        \ML_int[4][46] ) );
  MUX2_X1 M1_3_45 ( .A(\ML_int[3][45] ), .B(\ML_int[3][37] ), .S(n59), .Z(
        \ML_int[4][45] ) );
  MUX2_X1 M1_3_44 ( .A(\ML_int[3][44] ), .B(\ML_int[3][36] ), .S(n59), .Z(
        \ML_int[4][44] ) );
  MUX2_X1 M1_3_43 ( .A(\ML_int[3][43] ), .B(\ML_int[3][35] ), .S(n58), .Z(
        \ML_int[4][43] ) );
  MUX2_X1 M1_3_42 ( .A(\ML_int[3][42] ), .B(\ML_int[3][34] ), .S(n58), .Z(
        \ML_int[4][42] ) );
  MUX2_X1 M1_3_41 ( .A(\ML_int[3][41] ), .B(\ML_int[3][33] ), .S(n58), .Z(
        \ML_int[4][41] ) );
  MUX2_X1 M1_3_40 ( .A(\ML_int[3][40] ), .B(\ML_int[3][32] ), .S(n58), .Z(
        \ML_int[4][40] ) );
  MUX2_X1 M1_3_39 ( .A(\ML_int[3][39] ), .B(\ML_int[3][31] ), .S(n58), .Z(
        \ML_int[4][39] ) );
  MUX2_X1 M1_3_38 ( .A(\ML_int[3][38] ), .B(\ML_int[3][30] ), .S(n58), .Z(
        \ML_int[4][38] ) );
  MUX2_X1 M1_3_37 ( .A(\ML_int[3][37] ), .B(\ML_int[3][29] ), .S(n58), .Z(
        \ML_int[4][37] ) );
  MUX2_X1 M1_3_36 ( .A(\ML_int[3][36] ), .B(\ML_int[3][28] ), .S(n58), .Z(
        \ML_int[4][36] ) );
  MUX2_X1 M1_3_35 ( .A(\ML_int[3][35] ), .B(\ML_int[3][27] ), .S(n58), .Z(
        \ML_int[4][35] ) );
  MUX2_X1 M1_3_34 ( .A(\ML_int[3][34] ), .B(\ML_int[3][26] ), .S(n58), .Z(
        \ML_int[4][34] ) );
  MUX2_X1 M1_3_33 ( .A(\ML_int[3][33] ), .B(\ML_int[3][25] ), .S(n58), .Z(
        \ML_int[4][33] ) );
  MUX2_X1 M1_3_32 ( .A(\ML_int[3][32] ), .B(\ML_int[3][24] ), .S(n58), .Z(
        \ML_int[4][32] ) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n57), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n57), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n57), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n57), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n57), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n57), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n56), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n56), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(n20), .B(\ML_int[3][9] ), .S(n56), .Z(\ML_int[4][17] )
         );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n56), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n56), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n56), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n56), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n56), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n56), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n56), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n56), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n56), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M1_2_46 ( .A(\ML_int[2][46] ), .B(\ML_int[2][42] ), .S(n54), .Z(
        \ML_int[3][46] ) );
  MUX2_X1 M1_2_45 ( .A(\ML_int[2][45] ), .B(\ML_int[2][41] ), .S(n51), .Z(
        \ML_int[3][45] ) );
  MUX2_X1 M1_2_44 ( .A(\ML_int[2][44] ), .B(\ML_int[2][40] ), .S(n53), .Z(
        \ML_int[3][44] ) );
  MUX2_X1 M1_2_43 ( .A(\ML_int[2][43] ), .B(\ML_int[2][39] ), .S(n53), .Z(
        \ML_int[3][43] ) );
  MUX2_X1 M1_2_42 ( .A(\ML_int[2][42] ), .B(\ML_int[2][38] ), .S(n51), .Z(
        \ML_int[3][42] ) );
  MUX2_X1 M1_2_41 ( .A(\ML_int[2][41] ), .B(\ML_int[2][37] ), .S(n53), .Z(
        \ML_int[3][41] ) );
  MUX2_X1 M1_2_40 ( .A(\ML_int[2][40] ), .B(\ML_int[2][36] ), .S(n54), .Z(
        \ML_int[3][40] ) );
  MUX2_X1 M1_2_39 ( .A(\ML_int[2][39] ), .B(\ML_int[2][35] ), .S(n53), .Z(
        \ML_int[3][39] ) );
  MUX2_X1 M1_2_38 ( .A(\ML_int[2][38] ), .B(\ML_int[2][34] ), .S(n53), .Z(
        \ML_int[3][38] ) );
  MUX2_X1 M1_2_37 ( .A(\ML_int[2][37] ), .B(\ML_int[2][33] ), .S(n54), .Z(
        \ML_int[3][37] ) );
  MUX2_X1 M1_2_36 ( .A(\ML_int[2][36] ), .B(\ML_int[2][32] ), .S(n51), .Z(
        \ML_int[3][36] ) );
  MUX2_X1 M1_2_35 ( .A(\ML_int[2][35] ), .B(\ML_int[2][31] ), .S(n53), .Z(
        \ML_int[3][35] ) );
  MUX2_X1 M1_2_34 ( .A(\ML_int[2][34] ), .B(\ML_int[2][30] ), .S(n53), .Z(
        \ML_int[3][34] ) );
  MUX2_X1 M1_2_33 ( .A(\ML_int[2][33] ), .B(\ML_int[2][29] ), .S(n54), .Z(
        \ML_int[3][33] ) );
  MUX2_X1 M1_2_32 ( .A(\ML_int[2][32] ), .B(\ML_int[2][28] ), .S(n51), .Z(
        \ML_int[3][32] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n54), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n52), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n51), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n52), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n52), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n52), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n53), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n52), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n54), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n52), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n51), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n51), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n54), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n54), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n51), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n53), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n51), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n53), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n54), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n51), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M1_1_46 ( .A(\ML_int[1][46] ), .B(\ML_int[1][44] ), .S(n49), .Z(
        \ML_int[2][46] ) );
  MUX2_X1 M1_1_45 ( .A(\ML_int[1][45] ), .B(\ML_int[1][43] ), .S(n11), .Z(
        \ML_int[2][45] ) );
  MUX2_X1 M1_1_44 ( .A(\ML_int[1][44] ), .B(\ML_int[1][42] ), .S(n11), .Z(
        \ML_int[2][44] ) );
  MUX2_X1 M1_1_43 ( .A(\ML_int[1][43] ), .B(\ML_int[1][41] ), .S(n47), .Z(
        \ML_int[2][43] ) );
  MUX2_X1 M1_1_42 ( .A(\ML_int[1][42] ), .B(\ML_int[1][40] ), .S(n11), .Z(
        \ML_int[2][42] ) );
  MUX2_X1 M1_1_41 ( .A(\ML_int[1][41] ), .B(\ML_int[1][39] ), .S(n11), .Z(
        \ML_int[2][41] ) );
  MUX2_X1 M1_1_40 ( .A(\ML_int[1][40] ), .B(\ML_int[1][38] ), .S(n49), .Z(
        \ML_int[2][40] ) );
  MUX2_X1 M1_1_39 ( .A(\ML_int[1][39] ), .B(\ML_int[1][37] ), .S(n49), .Z(
        \ML_int[2][39] ) );
  MUX2_X1 M1_1_38 ( .A(\ML_int[1][38] ), .B(\ML_int[1][36] ), .S(n47), .Z(
        \ML_int[2][38] ) );
  MUX2_X1 M1_1_37 ( .A(\ML_int[1][37] ), .B(\ML_int[1][35] ), .S(n46), .Z(
        \ML_int[2][37] ) );
  MUX2_X1 M1_1_36 ( .A(\ML_int[1][36] ), .B(\ML_int[1][34] ), .S(n46), .Z(
        \ML_int[2][36] ) );
  MUX2_X1 M1_1_35 ( .A(\ML_int[1][35] ), .B(\ML_int[1][33] ), .S(n21), .Z(
        \ML_int[2][35] ) );
  MUX2_X1 M1_1_34 ( .A(\ML_int[1][34] ), .B(\ML_int[1][32] ), .S(n46), .Z(
        \ML_int[2][34] ) );
  MUX2_X1 M1_1_33 ( .A(\ML_int[1][33] ), .B(\ML_int[1][31] ), .S(n21), .Z(
        \ML_int[2][33] ) );
  MUX2_X1 M1_1_32 ( .A(\ML_int[1][32] ), .B(\ML_int[1][30] ), .S(n22), .Z(
        \ML_int[2][32] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n21), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n47), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n22), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n22), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n48), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n46), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n22), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n47), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n48), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n21), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(n24), .B(\ML_int[1][16] ), .S(n47), .Z(\ML_int[2][18] )
         );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n48), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n22), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n48), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n21), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n48), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n21), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n46), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n47), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n46), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n21), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n46), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n49), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(n62), .S(n49), .Z(\ML_int[2][2] ) );
  MUX2_X1 M1_0_46 ( .A(A[46]), .B(A[45]), .S(n16), .Z(\ML_int[1][46] ) );
  MUX2_X1 M1_0_45 ( .A(A[45]), .B(A[44]), .S(n16), .Z(\ML_int[1][45] ) );
  MUX2_X1 M1_0_44 ( .A(A[44]), .B(A[43]), .S(n44), .Z(\ML_int[1][44] ) );
  MUX2_X1 M1_0_43 ( .A(A[43]), .B(A[42]), .S(n16), .Z(\ML_int[1][43] ) );
  MUX2_X1 M1_0_42 ( .A(A[42]), .B(A[41]), .S(n16), .Z(\ML_int[1][42] ) );
  MUX2_X1 M1_0_41 ( .A(A[41]), .B(A[40]), .S(n44), .Z(\ML_int[1][41] ) );
  MUX2_X1 M1_0_40 ( .A(A[40]), .B(A[39]), .S(n44), .Z(\ML_int[1][40] ) );
  MUX2_X1 M1_0_39 ( .A(A[39]), .B(A[38]), .S(n16), .Z(\ML_int[1][39] ) );
  MUX2_X1 M1_0_38 ( .A(A[38]), .B(A[37]), .S(n16), .Z(\ML_int[1][38] ) );
  MUX2_X1 M1_0_37 ( .A(A[37]), .B(A[36]), .S(n44), .Z(\ML_int[1][37] ) );
  MUX2_X1 M1_0_36 ( .A(A[36]), .B(A[35]), .S(n25), .Z(\ML_int[1][36] ) );
  MUX2_X1 M1_0_35 ( .A(A[35]), .B(A[34]), .S(n37), .Z(\ML_int[1][35] ) );
  MUX2_X1 M1_0_34 ( .A(A[34]), .B(A[33]), .S(n34), .Z(\ML_int[1][34] ) );
  MUX2_X1 M1_0_33 ( .A(A[33]), .B(A[32]), .S(n33), .Z(\ML_int[1][33] ) );
  MUX2_X1 M1_0_32 ( .A(A[32]), .B(A[31]), .S(n33), .Z(\ML_int[1][32] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n25), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n33), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n37), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n34), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n25), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n41), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n37), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n32), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n44), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n36), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n35), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n32), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n44), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n39), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n38), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n44), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n38), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n44), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n36), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n35), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n44), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n26), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n32), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n39), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n26), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n44), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n16), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n44), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n34), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n36), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n44), .Z(\ML_int[1][1] ) );
  BUF_X1 U3 ( .A(SH[4]), .Z(n60) );
  NAND2_X1 U4 ( .A1(\ML_int[2][29] ), .A2(n10), .ZN(n1) );
  NAND2_X1 U5 ( .A1(\ML_int[2][25] ), .A2(n52), .ZN(n2) );
  NAND2_X1 U6 ( .A1(n1), .A2(n2), .ZN(\ML_int[3][29] ) );
  MUX2_X1 U7 ( .A(\ML_int[1][28] ), .B(\ML_int[1][30] ), .S(n12), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 U8 ( .A(\ML_int[1][27] ), .B(\ML_int[1][29] ), .S(n50), .Z(
        \ML_int[2][29] ) );
  NAND2_X1 U9 ( .A1(\ML_int[1][25] ), .A2(n12), .ZN(n3) );
  NAND2_X1 U10 ( .A1(\ML_int[1][23] ), .A2(n47), .ZN(n4) );
  NAND2_X1 U11 ( .A1(n3), .A2(n4), .ZN(\ML_int[2][25] ) );
  MUX2_X1 U12 ( .A(\ML_int[4][30] ), .B(\ML_int[4][46] ), .S(n5), .Z(
        \ML_int[5][46] ) );
  MUX2_X1 U13 ( .A(\ML_int[4][29] ), .B(\ML_int[4][45] ), .S(n5), .Z(
        \ML_int[5][45] ) );
  NAND2_X1 U14 ( .A1(\ML_int[4][38] ), .A2(n5), .ZN(n6) );
  NAND2_X1 U15 ( .A1(\ML_int[4][22] ), .A2(n60), .ZN(n7) );
  NAND2_X1 U16 ( .A1(n6), .A2(n7), .ZN(\ML_int[5][38] ) );
  INV_X1 U17 ( .A(n60), .ZN(n5) );
  NAND2_X1 U18 ( .A1(\ML_int[4][37] ), .A2(n5), .ZN(n8) );
  NAND2_X1 U19 ( .A1(\ML_int[4][21] ), .A2(n60), .ZN(n9) );
  NAND2_X1 U20 ( .A1(n8), .A2(n9), .ZN(\ML_int[5][37] ) );
  INV_X2 U21 ( .A(SH[2]), .ZN(n10) );
  INV_X1 U22 ( .A(SH[2]), .ZN(n55) );
  INV_X1 U23 ( .A(n40), .ZN(n46) );
  INV_X1 U24 ( .A(n12), .ZN(n11) );
  INV_X1 U25 ( .A(n12), .ZN(n49) );
  INV_X1 U26 ( .A(SH[1]), .ZN(n12) );
  MUX2_X1 U27 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n59), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 U28 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n57), .Z(n13) );
  NAND2_X1 U29 ( .A1(\ML_int[3][28] ), .A2(n29), .ZN(n14) );
  NAND2_X1 U30 ( .A1(\ML_int[3][20] ), .A2(n57), .ZN(n15) );
  NAND2_X1 U31 ( .A1(n14), .A2(n15), .ZN(\ML_int[4][28] ) );
  BUF_X1 U32 ( .A(n42), .Z(n36) );
  INV_X1 U33 ( .A(SH[1]), .ZN(n50) );
  INV_X1 U34 ( .A(n23), .ZN(n16) );
  INV_X1 U35 ( .A(n16), .ZN(n17) );
  BUF_X1 U36 ( .A(n41), .Z(n39) );
  BUF_X1 U37 ( .A(n42), .Z(n38) );
  INV_X2 U38 ( .A(n23), .ZN(n44) );
  MUX2_X1 U39 ( .A(\ML_int[3][14] ), .B(\ML_int[3][22] ), .S(n29), .Z(
        \ML_int[4][22] ) );
  BUF_X2 U40 ( .A(SH[3]), .Z(n57) );
  MUX2_X1 U41 ( .A(\ML_int[2][8] ), .B(\ML_int[2][12] ), .S(n10), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 U42 ( .A(\ML_int[2][6] ), .B(\ML_int[2][10] ), .S(n10), .Z(
        \ML_int[3][10] ) );
  INV_X1 U43 ( .A(n55), .ZN(n51) );
  MUX2_X1 U44 ( .A(\ML_int[2][24] ), .B(\ML_int[2][28] ), .S(n10), .Z(
        \ML_int[3][28] ) );
  INV_X1 U45 ( .A(n55), .ZN(n53) );
  MUX2_X1 U46 ( .A(\ML_int[3][13] ), .B(\ML_int[3][21] ), .S(n29), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 U47 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n57), .Z(n18) );
  MUX2_X1 U48 ( .A(\ML_int[2][11] ), .B(\ML_int[2][15] ), .S(n10), .Z(
        \ML_int[3][15] ) );
  INV_X1 U49 ( .A(n40), .ZN(n47) );
  MUX2_X1 U50 ( .A(\ML_int[2][12] ), .B(\ML_int[2][16] ), .S(n10), .Z(
        \ML_int[3][16] ) );
  INV_X1 U51 ( .A(n55), .ZN(n52) );
  MUX2_X1 U52 ( .A(\ML_int[1][12] ), .B(\ML_int[1][14] ), .S(n12), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 U53 ( .A(\ML_int[2][17] ), .B(\ML_int[2][21] ), .S(n10), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 U54 ( .A(\ML_int[1][15] ), .B(\ML_int[1][17] ), .S(n50), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 U55 ( .A(\ML_int[3][16] ), .B(\ML_int[3][24] ), .S(n29), .Z(n19) );
  MUX2_X1 U56 ( .A(\ML_int[1][10] ), .B(\ML_int[1][12] ), .S(n50), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 U57 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n54), .Z(n20) );
  INV_X1 U58 ( .A(n40), .ZN(n21) );
  INV_X1 U59 ( .A(n50), .ZN(n22) );
  INV_X1 U60 ( .A(n40), .ZN(n48) );
  INV_X1 U61 ( .A(SH[0]), .ZN(n23) );
  MUX2_X1 U62 ( .A(\ML_int[3][16] ), .B(\ML_int[3][24] ), .S(n29), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 U63 ( .A(A[18]), .B(A[17]), .S(n16), .Z(n24) );
  BUF_X1 U64 ( .A(n43), .Z(n25) );
  BUF_X1 U65 ( .A(n42), .Z(n26) );
  MUX2_X1 U66 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n57), .Z(n27) );
  MUX2_X1 U67 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n57), .Z(n28) );
  MUX2_X1 U68 ( .A(\ML_int[2][16] ), .B(\ML_int[2][20] ), .S(n10), .Z(
        \ML_int[3][20] ) );
  NAND2_X1 U69 ( .A1(\ML_int[3][27] ), .A2(n29), .ZN(n30) );
  NAND2_X1 U70 ( .A1(\ML_int[3][19] ), .A2(n57), .ZN(n31) );
  NAND2_X1 U71 ( .A1(n30), .A2(n31), .ZN(\ML_int[4][27] ) );
  INV_X1 U72 ( .A(n57), .ZN(n29) );
  BUF_X1 U73 ( .A(n42), .Z(n32) );
  BUF_X1 U74 ( .A(n43), .Z(n33) );
  BUF_X1 U75 ( .A(n43), .Z(n34) );
  BUF_X1 U76 ( .A(n43), .Z(n35) );
  BUF_X1 U77 ( .A(n43), .Z(n37) );
  INV_X1 U78 ( .A(n23), .ZN(n41) );
  INV_X1 U79 ( .A(n45), .ZN(n42) );
  INV_X1 U80 ( .A(n45), .ZN(n43) );
  BUF_X1 U81 ( .A(SH[4]), .Z(n61) );
  BUF_X1 U82 ( .A(SH[3]), .Z(n56) );
  BUF_X1 U83 ( .A(SH[3]), .Z(n58) );
  INV_X1 U84 ( .A(SH[0]), .ZN(n45) );
  INV_X1 U85 ( .A(n65), .ZN(n62) );
  INV_X1 U86 ( .A(\ML_int[1][1] ), .ZN(n63) );
  INV_X1 U87 ( .A(SH[1]), .ZN(n40) );
  INV_X1 U88 ( .A(n55), .ZN(n54) );
  BUF_X1 U89 ( .A(SH[3]), .Z(n59) );
  AND2_X1 U90 ( .A1(\ML_int[2][3] ), .A2(n10), .ZN(\ML_int[3][3] ) );
  AND2_X1 U91 ( .A1(\ML_int[2][2] ), .A2(n10), .ZN(\ML_int[3][2] ) );
  NOR2_X1 U92 ( .A1(n64), .A2(n63), .ZN(\ML_int[3][1] ) );
  NOR2_X1 U93 ( .A1(n64), .A2(n65), .ZN(\ML_int[3][0] ) );
  NAND2_X1 U94 ( .A1(n50), .A2(n10), .ZN(n64) );
  NOR2_X1 U95 ( .A1(n11), .A2(n63), .ZN(\ML_int[2][1] ) );
  NOR2_X1 U96 ( .A1(n11), .A2(n65), .ZN(\ML_int[2][0] ) );
  NAND2_X1 U97 ( .A1(A[0]), .A2(n17), .ZN(n65) );
endmodule


module FP_MULTIPLIER_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module FP_MULTIPLIER_DW01_add_1 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , \A[15] ,
         \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] ,
         \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132;
  assign SUM[22] = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  OR2_X1 U2 ( .A1(B[24]), .A2(A[24]), .ZN(n17) );
  INV_X1 U3 ( .A(n17), .ZN(n130) );
  XOR2_X1 U4 ( .A(n27), .B(n78), .Z(SUM[38]) );
  AND2_X1 U5 ( .A1(n30), .A2(n132), .ZN(SUM[23]) );
  XOR2_X1 U6 ( .A(n25), .B(n101), .Z(SUM[32]) );
  CLKBUF_X1 U7 ( .A(n75), .Z(n3) );
  OAI21_X1 U8 ( .B1(n110), .B2(n109), .A(n111), .ZN(n4) );
  AOI21_X1 U9 ( .B1(n75), .B2(n38), .A(n76), .ZN(n5) );
  CLKBUF_X1 U10 ( .A(n83), .Z(n6) );
  CLKBUF_X1 U11 ( .A(n96), .Z(n7) );
  AOI21_X1 U12 ( .B1(n3), .B2(n38), .A(n76), .ZN(n16) );
  CLKBUF_X1 U13 ( .A(A[23]), .Z(n8) );
  AND2_X1 U14 ( .A1(n8), .A2(B[23]), .ZN(n9) );
  CLKBUF_X1 U15 ( .A(n121), .Z(n10) );
  CLKBUF_X1 U16 ( .A(n88), .Z(n11) );
  CLKBUF_X1 U17 ( .A(n126), .Z(n12) );
  OAI21_X1 U18 ( .B1(n5), .B2(n72), .A(n73), .ZN(n13) );
  OAI21_X1 U19 ( .B1(n72), .B2(n16), .A(n73), .ZN(n14) );
  OAI21_X1 U20 ( .B1(n103), .B2(n102), .A(n104), .ZN(n15) );
  AND2_X1 U21 ( .A1(A[23]), .A2(B[23]), .ZN(n24) );
  INV_X1 U22 ( .A(n9), .ZN(n132) );
  CLKBUF_X1 U23 ( .A(n113), .Z(n18) );
  CLKBUF_X1 U24 ( .A(n4), .Z(n19) );
  CLKBUF_X1 U25 ( .A(n110), .Z(n20) );
  AOI21_X1 U26 ( .B1(n13), .B2(n36), .A(n69), .ZN(n21) );
  OAI21_X1 U27 ( .B1(n21), .B2(n65), .A(n67), .ZN(n22) );
  AOI21_X1 U28 ( .B1(n40), .B2(n6), .A(n84), .ZN(n23) );
  CLKBUF_X1 U29 ( .A(n15), .Z(n25) );
  CLKBUF_X1 U30 ( .A(n91), .Z(n26) );
  OAI21_X1 U31 ( .B1(n79), .B2(n23), .A(n81), .ZN(n27) );
  XNOR2_X1 U32 ( .A(n52), .B(B[45]), .ZN(SUM[45]) );
  AOI21_X1 U33 ( .B1(n34), .B2(n22), .A(n62), .ZN(n28) );
  CLKBUF_X1 U34 ( .A(n103), .Z(n29) );
  XOR2_X1 U35 ( .A(n9), .B(n131), .Z(SUM[24]) );
  INV_X1 U36 ( .A(n87), .ZN(n41) );
  INV_X1 U37 ( .A(n109), .ZN(n47) );
  INV_X1 U38 ( .A(n102), .ZN(n45) );
  INV_X1 U39 ( .A(n79), .ZN(n39) );
  INV_X1 U40 ( .A(n95), .ZN(n43) );
  INV_X1 U41 ( .A(n57), .ZN(n33) );
  INV_X1 U42 ( .A(n125), .ZN(n51) );
  INV_X1 U43 ( .A(n117), .ZN(n49) );
  INV_X1 U44 ( .A(n72), .ZN(n37) );
  INV_X1 U45 ( .A(n65), .ZN(n35) );
  INV_X1 U46 ( .A(n77), .ZN(n38) );
  INV_X1 U47 ( .A(n107), .ZN(n46) );
  INV_X1 U48 ( .A(n100), .ZN(n44) );
  INV_X1 U49 ( .A(n70), .ZN(n36) );
  INV_X1 U50 ( .A(n85), .ZN(n40) );
  INV_X1 U51 ( .A(n93), .ZN(n42) );
  INV_X1 U52 ( .A(n63), .ZN(n34) );
  INV_X1 U53 ( .A(n115), .ZN(n48) );
  INV_X1 U54 ( .A(n123), .ZN(n50) );
  INV_X1 U55 ( .A(n55), .ZN(n32) );
  OR2_X1 U56 ( .A1(B[23]), .A2(n8), .ZN(n30) );
  CLKBUF_X1 U57 ( .A(n118), .Z(n31) );
  AOI21_X1 U58 ( .B1(n53), .B2(n32), .A(n54), .ZN(n52) );
  XOR2_X1 U59 ( .A(n53), .B(n56), .Z(SUM[44]) );
  NOR2_X1 U60 ( .A1(n54), .A2(n55), .ZN(n56) );
  NOR2_X1 U61 ( .A1(B[44]), .A2(A[44]), .ZN(n55) );
  AND2_X1 U62 ( .A1(B[44]), .A2(A[44]), .ZN(n54) );
  OAI21_X1 U63 ( .B1(n58), .B2(n57), .A(n59), .ZN(n53) );
  XOR2_X1 U64 ( .A(n60), .B(n28), .Z(SUM[43]) );
  AOI21_X1 U65 ( .B1(n61), .B2(n34), .A(n62), .ZN(n58) );
  NAND2_X1 U66 ( .A1(n33), .A2(n59), .ZN(n60) );
  NAND2_X1 U67 ( .A1(B[43]), .A2(A[43]), .ZN(n59) );
  NOR2_X1 U68 ( .A1(B[43]), .A2(A[43]), .ZN(n57) );
  XOR2_X1 U69 ( .A(n61), .B(n64), .Z(SUM[42]) );
  NOR2_X1 U70 ( .A1(n62), .A2(n63), .ZN(n64) );
  NOR2_X1 U71 ( .A1(B[42]), .A2(A[42]), .ZN(n63) );
  AND2_X1 U72 ( .A1(B[42]), .A2(A[42]), .ZN(n62) );
  OAI21_X1 U73 ( .B1(n66), .B2(n65), .A(n67), .ZN(n61) );
  XOR2_X1 U74 ( .A(n68), .B(n21), .Z(SUM[41]) );
  AOI21_X1 U75 ( .B1(n13), .B2(n36), .A(n69), .ZN(n66) );
  NAND2_X1 U76 ( .A1(n35), .A2(n67), .ZN(n68) );
  NAND2_X1 U77 ( .A1(B[41]), .A2(A[41]), .ZN(n67) );
  NOR2_X1 U78 ( .A1(B[41]), .A2(A[41]), .ZN(n65) );
  XOR2_X1 U79 ( .A(n14), .B(n71), .Z(SUM[40]) );
  NOR2_X1 U80 ( .A1(n69), .A2(n70), .ZN(n71) );
  NOR2_X1 U81 ( .A1(B[40]), .A2(A[40]), .ZN(n70) );
  AND2_X1 U82 ( .A1(B[40]), .A2(A[40]), .ZN(n69) );
  XOR2_X1 U83 ( .A(n74), .B(n16), .Z(SUM[39]) );
  NAND2_X1 U84 ( .A1(n37), .A2(n73), .ZN(n74) );
  NAND2_X1 U85 ( .A1(B[39]), .A2(A[39]), .ZN(n73) );
  NOR2_X1 U86 ( .A1(B[39]), .A2(A[39]), .ZN(n72) );
  NOR2_X1 U87 ( .A1(n76), .A2(n77), .ZN(n78) );
  NOR2_X1 U88 ( .A1(B[38]), .A2(A[38]), .ZN(n77) );
  AND2_X1 U89 ( .A1(B[38]), .A2(A[38]), .ZN(n76) );
  OAI21_X1 U90 ( .B1(n80), .B2(n79), .A(n81), .ZN(n75) );
  XOR2_X1 U91 ( .A(n82), .B(n23), .Z(SUM[37]) );
  AOI21_X1 U92 ( .B1(n83), .B2(n40), .A(n84), .ZN(n80) );
  NAND2_X1 U93 ( .A1(n39), .A2(n81), .ZN(n82) );
  NAND2_X1 U94 ( .A1(B[37]), .A2(A[37]), .ZN(n81) );
  NOR2_X1 U95 ( .A1(B[37]), .A2(A[37]), .ZN(n79) );
  XOR2_X1 U96 ( .A(n6), .B(n86), .Z(SUM[36]) );
  NOR2_X1 U97 ( .A1(n84), .A2(n85), .ZN(n86) );
  NOR2_X1 U98 ( .A1(B[36]), .A2(A[36]), .ZN(n85) );
  AND2_X1 U99 ( .A1(B[36]), .A2(A[36]), .ZN(n84) );
  OAI21_X1 U100 ( .B1(n88), .B2(n87), .A(n89), .ZN(n83) );
  XOR2_X1 U101 ( .A(n90), .B(n11), .Z(SUM[35]) );
  AOI21_X1 U102 ( .B1(n91), .B2(n42), .A(n92), .ZN(n88) );
  NAND2_X1 U103 ( .A1(n41), .A2(n89), .ZN(n90) );
  NAND2_X1 U104 ( .A1(B[35]), .A2(A[35]), .ZN(n89) );
  NOR2_X1 U105 ( .A1(B[35]), .A2(A[35]), .ZN(n87) );
  XOR2_X1 U106 ( .A(n26), .B(n94), .Z(SUM[34]) );
  NOR2_X1 U107 ( .A1(n92), .A2(n93), .ZN(n94) );
  NOR2_X1 U108 ( .A1(B[34]), .A2(A[34]), .ZN(n93) );
  AND2_X1 U109 ( .A1(B[34]), .A2(A[34]), .ZN(n92) );
  OAI21_X1 U110 ( .B1(n96), .B2(n95), .A(n97), .ZN(n91) );
  XOR2_X1 U111 ( .A(n98), .B(n7), .Z(SUM[33]) );
  AOI21_X1 U112 ( .B1(n15), .B2(n44), .A(n99), .ZN(n96) );
  NAND2_X1 U113 ( .A1(n43), .A2(n97), .ZN(n98) );
  NAND2_X1 U114 ( .A1(B[33]), .A2(A[33]), .ZN(n97) );
  NOR2_X1 U115 ( .A1(B[33]), .A2(A[33]), .ZN(n95) );
  NOR2_X1 U116 ( .A1(n99), .A2(n100), .ZN(n101) );
  NOR2_X1 U117 ( .A1(B[32]), .A2(A[32]), .ZN(n100) );
  AND2_X1 U118 ( .A1(B[32]), .A2(A[32]), .ZN(n99) );
  XOR2_X1 U119 ( .A(n105), .B(n29), .Z(SUM[31]) );
  AOI21_X1 U120 ( .B1(n4), .B2(n46), .A(n106), .ZN(n103) );
  NAND2_X1 U121 ( .A1(n45), .A2(n104), .ZN(n105) );
  NAND2_X1 U122 ( .A1(B[31]), .A2(A[31]), .ZN(n104) );
  NOR2_X1 U123 ( .A1(B[31]), .A2(A[31]), .ZN(n102) );
  XOR2_X1 U124 ( .A(n19), .B(n108), .Z(SUM[30]) );
  NOR2_X1 U125 ( .A1(n106), .A2(n107), .ZN(n108) );
  NOR2_X1 U126 ( .A1(B[30]), .A2(A[30]), .ZN(n107) );
  AND2_X1 U127 ( .A1(B[30]), .A2(A[30]), .ZN(n106) );
  XOR2_X1 U128 ( .A(n112), .B(n20), .Z(SUM[29]) );
  AOI21_X1 U129 ( .B1(n113), .B2(n48), .A(n114), .ZN(n110) );
  NAND2_X1 U130 ( .A1(n47), .A2(n111), .ZN(n112) );
  NAND2_X1 U131 ( .A1(B[29]), .A2(A[29]), .ZN(n111) );
  NOR2_X1 U132 ( .A1(B[29]), .A2(A[29]), .ZN(n109) );
  XOR2_X1 U133 ( .A(n18), .B(n116), .Z(SUM[28]) );
  NOR2_X1 U134 ( .A1(n114), .A2(n115), .ZN(n116) );
  NOR2_X1 U135 ( .A1(B[28]), .A2(A[28]), .ZN(n115) );
  AND2_X1 U136 ( .A1(B[28]), .A2(A[28]), .ZN(n114) );
  OAI21_X1 U137 ( .B1(n118), .B2(n117), .A(n119), .ZN(n113) );
  XOR2_X1 U138 ( .A(n120), .B(n31), .Z(SUM[27]) );
  AOI21_X1 U139 ( .B1(n121), .B2(n50), .A(n122), .ZN(n118) );
  NAND2_X1 U140 ( .A1(n49), .A2(n119), .ZN(n120) );
  NAND2_X1 U141 ( .A1(B[27]), .A2(A[27]), .ZN(n119) );
  NOR2_X1 U142 ( .A1(B[27]), .A2(A[27]), .ZN(n117) );
  XOR2_X1 U143 ( .A(n10), .B(n124), .Z(SUM[26]) );
  NOR2_X1 U144 ( .A1(n122), .A2(n123), .ZN(n124) );
  NOR2_X1 U145 ( .A1(B[26]), .A2(A[26]), .ZN(n123) );
  AND2_X1 U146 ( .A1(B[26]), .A2(A[26]), .ZN(n122) );
  OAI21_X1 U147 ( .B1(n126), .B2(n125), .A(n127), .ZN(n121) );
  XOR2_X1 U148 ( .A(n128), .B(n12), .Z(SUM[25]) );
  AOI21_X1 U149 ( .B1(n24), .B2(n17), .A(n129), .ZN(n126) );
  NAND2_X1 U150 ( .A1(n51), .A2(n127), .ZN(n128) );
  NAND2_X1 U151 ( .A1(B[25]), .A2(A[25]), .ZN(n127) );
  NOR2_X1 U152 ( .A1(B[25]), .A2(A[25]), .ZN(n125) );
  NOR2_X1 U153 ( .A1(n129), .A2(n130), .ZN(n131) );
  AND2_X1 U154 ( .A1(B[24]), .A2(A[24]), .ZN(n129) );
endmodule


module FP_MULTIPLIER_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   \ab[23][22] , \ab[23][21] , \ab[23][20] , \ab[23][19] , \ab[23][18] ,
         \ab[23][17] , \ab[23][16] , \ab[23][15] , \ab[23][14] , \ab[23][13] ,
         \ab[23][12] , \ab[23][11] , \ab[23][10] , \ab[23][9] , \ab[23][8] ,
         \ab[23][7] , \ab[23][6] , \ab[23][5] , \ab[23][4] , \ab[23][3] ,
         \ab[23][2] , \ab[23][1] , \ab[23][0] , \ab[22][23] , \ab[22][22] ,
         \ab[22][21] , \ab[22][20] , \ab[22][19] , \ab[22][18] , \ab[22][17] ,
         \ab[22][16] , \ab[22][15] , \ab[22][14] , \ab[22][13] , \ab[22][12] ,
         \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] , \ab[22][7] ,
         \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] , \ab[22][2] ,
         \ab[22][1] , \ab[22][0] , \ab[21][23] , \ab[21][22] , \ab[21][21] ,
         \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] , \ab[21][16] ,
         \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] , \ab[21][11] ,
         \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] , \ab[21][6] ,
         \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] , \ab[21][1] ,
         \ab[21][0] , \ab[20][23] , \ab[20][22] , \ab[20][21] , \ab[20][20] ,
         \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] , \ab[20][15] ,
         \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] , \ab[20][10] ,
         \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][5] ,
         \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] ,
         \ab[19][23] , \ab[19][22] , \ab[19][21] , \ab[19][20] , \ab[19][19] ,
         \ab[19][18] , \ab[19][17] , \ab[19][16] , \ab[19][15] , \ab[19][14] ,
         \ab[19][13] , \ab[19][12] , \ab[19][11] , \ab[19][10] , \ab[19][9] ,
         \ab[19][8] , \ab[19][7] , \ab[19][6] , \ab[19][5] , \ab[19][4] ,
         \ab[19][3] , \ab[19][2] , \ab[19][1] , \ab[19][0] , \ab[18][23] ,
         \ab[18][22] , \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] ,
         \ab[18][17] , \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] ,
         \ab[18][12] , \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] ,
         \ab[18][7] , \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] ,
         \ab[18][2] , \ab[18][1] , \ab[18][0] , \ab[17][23] , \ab[17][22] ,
         \ab[17][21] , \ab[17][20] , \ab[17][19] , \ab[17][18] , \ab[17][17] ,
         \ab[17][16] , \ab[17][15] , \ab[17][14] , \ab[17][13] , \ab[17][12] ,
         \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] , \ab[17][7] ,
         \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] , \ab[17][2] ,
         \ab[17][1] , \ab[17][0] , \ab[16][23] , \ab[16][22] , \ab[16][21] ,
         \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] , \ab[16][16] ,
         \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] , \ab[16][11] ,
         \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] , \ab[16][6] ,
         \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] , \ab[16][1] ,
         \ab[16][0] , \ab[15][23] , \ab[15][22] , \ab[15][21] , \ab[15][20] ,
         \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] , \ab[15][15] ,
         \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] , \ab[15][10] ,
         \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] , \ab[15][5] ,
         \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] , \ab[15][0] ,
         \ab[14][23] , \ab[14][22] , \ab[14][21] , \ab[14][20] , \ab[14][19] ,
         \ab[14][18] , \ab[14][17] , \ab[14][16] , \ab[14][15] , \ab[14][14] ,
         \ab[14][13] , \ab[14][12] , \ab[14][11] , \ab[14][10] , \ab[14][9] ,
         \ab[14][8] , \ab[14][7] , \ab[14][6] , \ab[14][5] , \ab[14][4] ,
         \ab[14][3] , \ab[14][2] , \ab[14][1] , \ab[14][0] , \ab[13][23] ,
         \ab[13][22] , \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] ,
         \ab[13][17] , \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][23] , \ab[12][22] ,
         \ab[12][21] , \ab[12][20] , \ab[12][19] , \ab[12][18] , \ab[12][17] ,
         \ab[12][16] , \ab[12][15] , \ab[12][14] , \ab[12][13] , \ab[12][12] ,
         \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] , \ab[12][7] ,
         \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] , \ab[12][2] ,
         \ab[12][1] , \ab[12][0] , \ab[11][23] , \ab[11][22] , \ab[11][21] ,
         \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] , \ab[11][16] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][23] , \ab[10][22] , \ab[10][21] , \ab[10][20] ,
         \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] , \ab[10][15] ,
         \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] ,
         \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] ,
         \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] ,
         \ab[9][23] , \ab[9][22] , \ab[9][21] , \ab[9][20] , \ab[9][19] ,
         \ab[9][18] , \ab[9][17] , \ab[9][16] , \ab[9][15] , \ab[9][14] ,
         \ab[9][13] , \ab[9][12] , \ab[9][11] , \ab[9][10] , \ab[9][9] ,
         \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] , \ab[9][4] ,
         \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] , \ab[8][23] ,
         \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] ,
         \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][23] , \ab[7][22] ,
         \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] , \ab[7][17] ,
         \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] , \ab[7][12] ,
         \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] , \ab[7][7] ,
         \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] , \ab[7][2] ,
         \ab[7][1] , \ab[7][0] , \ab[6][23] , \ab[6][22] , \ab[6][21] ,
         \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] , \ab[6][16] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][23] , \ab[5][22] , \ab[5][21] , \ab[5][20] ,
         \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][15] ,
         \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] ,
         \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][23] , \ab[4][22] , \ab[4][21] , \ab[4][20] , \ab[4][19] ,
         \ab[4][18] , \ab[4][17] , \ab[4][16] , \ab[4][15] , \ab[4][14] ,
         \ab[4][13] , \ab[4][12] , \ab[4][11] , \ab[4][10] , \ab[4][9] ,
         \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] ,
         \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][23] ,
         \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] ,
         \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][23] , \ab[2][22] ,
         \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] , \ab[2][17] ,
         \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] , \ab[2][12] ,
         \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] , \ab[2][7] ,
         \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] , \ab[2][2] ,
         \ab[2][1] , \ab[2][0] , \ab[1][23] , \ab[1][22] , \ab[1][21] ,
         \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] , \ab[1][16] ,
         \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] ,
         \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[1][0] , \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] ,
         \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] ,
         \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][22] , \CARRYB[22][21] , \CARRYB[22][20] ,
         \CARRYB[22][19] , \CARRYB[22][18] , \CARRYB[22][17] ,
         \CARRYB[22][16] , \CARRYB[22][15] , \CARRYB[22][14] ,
         \CARRYB[22][13] , \CARRYB[22][12] , \CARRYB[22][11] ,
         \CARRYB[22][10] , \CARRYB[22][9] , \CARRYB[22][8] , \CARRYB[22][7] ,
         \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] ,
         \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][22] , \CARRYB[20][21] , \CARRYB[20][20] ,
         \CARRYB[20][19] , \CARRYB[20][18] , \CARRYB[20][17] ,
         \CARRYB[20][16] , \CARRYB[20][15] , \CARRYB[20][14] ,
         \CARRYB[20][13] , \CARRYB[20][12] , \CARRYB[20][11] ,
         \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] , \CARRYB[20][7] ,
         \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] , \CARRYB[20][3] ,
         \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] , \CARRYB[19][22] ,
         \CARRYB[19][21] , \CARRYB[19][20] , \CARRYB[19][19] ,
         \CARRYB[19][18] , \CARRYB[19][17] , \CARRYB[19][16] ,
         \CARRYB[19][15] , \CARRYB[19][14] , \CARRYB[19][13] ,
         \CARRYB[19][12] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] ,
         \CARRYB[19][8] , \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] ,
         \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] ,
         \CARRYB[19][0] , \CARRYB[18][22] , \CARRYB[18][21] , \CARRYB[18][20] ,
         \CARRYB[18][19] , \CARRYB[18][18] , \CARRYB[18][17] ,
         \CARRYB[18][16] , \CARRYB[18][15] , \CARRYB[18][14] ,
         \CARRYB[18][13] , \CARRYB[18][12] , \CARRYB[18][11] ,
         \CARRYB[18][10] , \CARRYB[18][9] , \CARRYB[18][8] , \CARRYB[18][7] ,
         \CARRYB[18][6] , \CARRYB[18][5] , \CARRYB[18][4] , \CARRYB[18][3] ,
         \CARRYB[18][2] , \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][22] ,
         \CARRYB[17][21] , \CARRYB[17][20] , \CARRYB[17][19] ,
         \CARRYB[17][18] , \CARRYB[17][17] , \CARRYB[17][16] ,
         \CARRYB[17][15] , \CARRYB[17][14] , \CARRYB[17][13] ,
         \CARRYB[17][12] , \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] ,
         \CARRYB[17][8] , \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][22] , \CARRYB[16][21] , \CARRYB[16][20] ,
         \CARRYB[16][19] , \CARRYB[16][18] , \CARRYB[16][17] ,
         \CARRYB[16][16] , \CARRYB[16][15] , \CARRYB[16][14] ,
         \CARRYB[16][13] , \CARRYB[16][12] , \CARRYB[16][11] ,
         \CARRYB[16][10] , \CARRYB[16][9] , \CARRYB[16][8] , \CARRYB[16][7] ,
         \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] , \CARRYB[16][3] ,
         \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] , \CARRYB[15][22] ,
         \CARRYB[15][21] , \CARRYB[15][20] , \CARRYB[15][19] ,
         \CARRYB[15][18] , \CARRYB[15][17] , \CARRYB[15][16] ,
         \CARRYB[15][15] , \CARRYB[15][14] , \CARRYB[15][13] ,
         \CARRYB[15][12] , \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] ,
         \CARRYB[15][8] , \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] ,
         \CARRYB[15][4] , \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] ,
         \CARRYB[15][0] , \CARRYB[14][22] , \CARRYB[14][21] , \CARRYB[14][20] ,
         \CARRYB[14][19] , \CARRYB[14][18] , \CARRYB[14][17] ,
         \CARRYB[14][16] , \CARRYB[14][15] , \CARRYB[14][14] ,
         \CARRYB[14][13] , \CARRYB[14][12] , \CARRYB[14][11] ,
         \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] , \CARRYB[14][7] ,
         \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] ,
         \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][22] , \CARRYB[12][21] , \CARRYB[12][20] ,
         \CARRYB[12][19] , \CARRYB[12][18] , \CARRYB[12][17] ,
         \CARRYB[12][16] , \CARRYB[12][15] , \CARRYB[12][14] ,
         \CARRYB[12][13] , \CARRYB[12][12] , \CARRYB[12][11] ,
         \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] , \CARRYB[12][7] ,
         \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] ,
         \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][22] , \CARRYB[10][21] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][22] ,
         \CARRYB[9][21] , \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] ,
         \CARRYB[9][17] , \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][22] , \CARRYB[8][21] ,
         \CARRYB[8][20] , \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] ,
         \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][22] ,
         \CARRYB[1][20] , \SUMB[23][22] , \SUMB[23][21] , \SUMB[23][20] ,
         \SUMB[23][19] , \SUMB[23][18] , \SUMB[23][17] , \SUMB[23][16] ,
         \SUMB[23][15] , \SUMB[23][14] , \SUMB[23][13] , \SUMB[23][12] ,
         \SUMB[23][11] , \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] ,
         \SUMB[23][7] , \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] ,
         \SUMB[23][3] , \SUMB[23][2] , \SUMB[23][1] , \SUMB[23][0] ,
         \SUMB[22][22] , \SUMB[22][21] , \SUMB[22][20] , \SUMB[22][19] ,
         \SUMB[22][18] , \SUMB[22][17] , \SUMB[22][16] , \SUMB[22][15] ,
         \SUMB[22][14] , \SUMB[22][13] , \SUMB[22][12] , \SUMB[22][11] ,
         \SUMB[22][10] , \SUMB[22][9] , \SUMB[22][8] , \SUMB[22][7] ,
         \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] , \SUMB[22][3] ,
         \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][22] , \SUMB[21][21] ,
         \SUMB[21][20] , \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] ,
         \SUMB[21][16] , \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] ,
         \SUMB[21][12] , \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] ,
         \SUMB[21][8] , \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] ,
         \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] ,
         \SUMB[20][22] , \SUMB[20][21] , \SUMB[20][20] , \SUMB[20][19] ,
         \SUMB[20][18] , \SUMB[20][17] , \SUMB[20][16] , \SUMB[20][15] ,
         \SUMB[20][14] , \SUMB[20][13] , \SUMB[20][12] , \SUMB[20][11] ,
         \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] ,
         \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] ,
         \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][22] , \SUMB[19][21] ,
         \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] ,
         \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] , \SUMB[19][13] ,
         \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] , \SUMB[19][9] ,
         \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] , \SUMB[19][5] ,
         \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] , \SUMB[19][1] ,
         \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] , \SUMB[18][19] ,
         \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] , \SUMB[18][15] ,
         \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] ,
         \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] ,
         \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] ,
         \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][22] , \SUMB[17][21] ,
         \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] ,
         \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] ,
         \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] ,
         \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] ,
         \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] , \SUMB[16][19] ,
         \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] , \SUMB[16][15] ,
         \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] , \SUMB[16][11] ,
         \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] , \SUMB[16][7] ,
         \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] ,
         \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][22] , \SUMB[15][21] ,
         \SUMB[15][20] , \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] ,
         \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] ,
         \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] ,
         \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] ,
         \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[14][22] , \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] ,
         \SUMB[14][18] , \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] ,
         \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] ,
         \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] ,
         \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] ,
         \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][22] , \SUMB[13][21] ,
         \SUMB[13][20] , \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] ,
         \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][22] , \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] ,
         \SUMB[12][18] , \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] ,
         \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] ,
         \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] ,
         \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] ,
         \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][22] , \SUMB[11][21] ,
         \SUMB[11][20] , \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] ,
         \SUMB[11][16] , \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] ,
         \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] ,
         \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] ,
         \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] ,
         \SUMB[10][22] , \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] ,
         \SUMB[10][18] , \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] ,
         \SUMB[10][14] , \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] ,
         \SUMB[10][10] , \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] ,
         \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] ,
         \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][22] , \SUMB[9][21] ,
         \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] ,
         \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][22] ,
         \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] ,
         \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] ,
         \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][22] ,
         \SUMB[1][20] , \A1[23] , \A1[20] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[24] , n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174;
  assign \ab[23][22]  = B[22];
  assign \ab[23][21]  = B[21];
  assign \ab[23][20]  = B[20];
  assign \ab[23][19]  = B[19];
  assign \ab[23][18]  = B[18];
  assign \ab[23][17]  = B[17];
  assign \ab[23][16]  = B[16];
  assign \ab[23][15]  = B[15];
  assign \ab[23][14]  = B[14];
  assign \ab[23][13]  = B[13];
  assign \ab[23][12]  = B[12];
  assign \ab[23][11]  = B[11];
  assign \ab[23][10]  = B[10];
  assign \ab[23][9]  = B[9];
  assign \ab[23][8]  = B[8];
  assign \ab[23][7]  = B[7];
  assign \ab[23][6]  = B[6];
  assign \ab[23][5]  = B[5];
  assign \ab[23][4]  = B[4];
  assign \ab[23][3]  = B[3];
  assign \ab[23][2]  = B[2];
  assign \ab[23][1]  = B[1];
  assign \ab[23][0]  = B[0];
  assign \ab[22][23]  = A[22];
  assign \ab[21][23]  = A[21];
  assign \ab[20][23]  = A[20];
  assign \ab[19][23]  = A[19];
  assign \ab[18][23]  = A[18];
  assign \ab[17][23]  = A[17];
  assign \ab[16][23]  = A[16];
  assign \ab[15][23]  = A[15];
  assign \ab[14][23]  = A[14];
  assign \ab[13][23]  = A[13];
  assign \ab[12][23]  = A[12];
  assign \ab[11][23]  = A[11];
  assign \ab[10][23]  = A[10];
  assign \ab[9][23]  = A[9];
  assign \ab[8][23]  = A[8];
  assign \ab[7][23]  = A[7];
  assign \ab[6][23]  = A[6];
  assign \ab[5][23]  = A[5];
  assign \ab[4][23]  = A[4];
  assign \ab[3][23]  = A[3];
  assign \ab[2][23]  = A[2];
  assign \ab[1][23]  = A[1];
  assign \ab[0][23]  = A[0];

  FA_X1 S4_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), .CO(
        \CARRYB[23][0] ), .S(\SUMB[23][0] ) );
  FA_X1 S4_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), .CO(
        \CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA_X1 S4_2 ( .A(\CARRYB[22][2] ), .B(\ab[23][2] ), .CI(\SUMB[22][3] ), .CO(
        \CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA_X1 S4_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), .CO(
        \CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA_X1 S4_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), .CO(
        \CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA_X1 S4_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), .CO(
        \CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA_X1 S4_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), .CO(
        \CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA_X1 S4_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), .CO(
        \CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA_X1 S4_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), .CO(
        \CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA_X1 S4_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), .CO(
        \CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA_X1 S4_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA_X1 S4_11 ( .A(\ab[23][11] ), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA_X1 S4_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA_X1 S4_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA_X1 S4_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA_X1 S4_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA_X1 S4_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA_X1 S4_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA_X1 S4_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA_X1 S4_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA_X1 S4_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA_X1 S4_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA_X1 S5_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\ab[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA_X1 S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FA_X1 S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA_X1 S2_22_2 ( .A(\CARRYB[21][2] ), .B(\ab[22][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA_X1 S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA_X1 S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA_X1 S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA_X1 S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA_X1 S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA_X1 S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA_X1 S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA_X1 S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA_X1 S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), 
        .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA_X1 S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), 
        .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA_X1 S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(\SUMB[21][14] ), 
        .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FA_X1 S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), 
        .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA_X1 S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA_X1 S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA_X1 S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA_X1 S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA_X1 S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA_X1 S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA_X1 S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA_X1 S3_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\ab[21][23] ), 
        .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA_X1 S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FA_X1 S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA_X1 S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA_X1 S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA_X1 S2_21_4 ( .A(\CARRYB[20][4] ), .B(\ab[21][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA_X1 S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA_X1 S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA_X1 S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA_X1 S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA_X1 S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA_X1 S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA_X1 S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA_X1 S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA_X1 S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA_X1 S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA_X1 S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA_X1 S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA_X1 S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA_X1 S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA_X1 S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA_X1 S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA_X1 S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA_X1 S3_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\ab[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA_X1 S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA_X1 S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA_X1 S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA_X1 S2_20_3 ( .A(\CARRYB[19][3] ), .B(\ab[20][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA_X1 S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA_X1 S2_20_5 ( .A(\CARRYB[19][5] ), .B(\ab[20][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA_X1 S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA_X1 S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA_X1 S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA_X1 S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA_X1 S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA_X1 S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA_X1 S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA_X1 S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA_X1 S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA_X1 S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA_X1 S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA_X1 S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA_X1 S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA_X1 S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA_X1 S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA_X1 S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA_X1 S3_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\ab[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA_X1 S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA_X1 S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA_X1 S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA_X1 S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA_X1 S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA_X1 S2_19_5 ( .A(\CARRYB[18][5] ), .B(\ab[19][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA_X1 S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA_X1 S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA_X1 S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA_X1 S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA_X1 S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA_X1 S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA_X1 S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA_X1 S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA_X1 S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA_X1 S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA_X1 S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA_X1 S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA_X1 S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA_X1 S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA_X1 S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA_X1 S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA_X1 S3_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\ab[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA_X1 S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA_X1 S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA_X1 S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA_X1 S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA_X1 S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA_X1 S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA_X1 S2_18_6 ( .A(\CARRYB[17][6] ), .B(\ab[18][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA_X1 S2_18_7 ( .A(\CARRYB[17][7] ), .B(\ab[18][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA_X1 S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA_X1 S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA_X1 S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA_X1 S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA_X1 S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA_X1 S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA_X1 S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA_X1 S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA_X1 S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA_X1 S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA_X1 S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA_X1 S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA_X1 S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA_X1 S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA_X1 S3_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\ab[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA_X1 S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA_X1 S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA_X1 S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA_X1 S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA_X1 S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA_X1 S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA_X1 S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA_X1 S2_17_7 ( .A(\CARRYB[16][7] ), .B(\ab[17][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA_X1 S2_17_8 ( .A(\CARRYB[16][8] ), .B(\ab[17][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA_X1 S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA_X1 S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA_X1 S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA_X1 S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA_X1 S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA_X1 S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA_X1 S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA_X1 S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA_X1 S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA_X1 S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA_X1 S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA_X1 S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA_X1 S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA_X1 S3_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\ab[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA_X1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA_X1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA_X1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA_X1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA_X1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA_X1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA_X1 S2_16_6 ( .A(\CARRYB[15][6] ), .B(\ab[16][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA_X1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA_X1 S2_16_8 ( .A(\CARRYB[15][8] ), .B(\ab[16][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA_X1 S2_16_9 ( .A(\CARRYB[15][9] ), .B(\ab[16][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA_X1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA_X1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA_X1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA_X1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA_X1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA_X1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA_X1 S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA_X1 S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA_X1 S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA_X1 S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA_X1 S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA_X1 S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA_X1 S3_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\ab[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA_X1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA_X1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S2_15_9 ( .A(\CARRYB[14][9] ), .B(\ab[15][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S2_15_10 ( .A(\CARRYB[14][10] ), .B(\ab[15][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA_X1 S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA_X1 S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA_X1 S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA_X1 S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA_X1 S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA_X1 S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA_X1 S3_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\ab[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\CARRYB[13][10] ), .B(\ab[14][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\CARRYB[13][11] ), .B(\ab[14][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA_X1 S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA_X1 S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA_X1 S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA_X1 S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA_X1 S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA_X1 S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA_X1 S3_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\ab[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\CARRYB[12][8] ), .B(\ab[13][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\CARRYB[12][9] ), .B(\ab[13][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\CARRYB[12][10] ), .B(\ab[13][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA_X1 S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA_X1 S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA_X1 S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA_X1 S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA_X1 S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA_X1 S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA_X1 S3_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\ab[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\CARRYB[11][9] ), .B(\ab[12][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\CARRYB[11][13] ), .B(\ab[12][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA_X1 S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA_X1 S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA_X1 S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA_X1 S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA_X1 S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA_X1 S3_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\ab[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\CARRYB[10][9] ), .B(\ab[11][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\CARRYB[10][10] ), .B(\ab[11][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\CARRYB[10][13] ), .B(\ab[11][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA_X1 S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA_X1 S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA_X1 S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA_X1 S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA_X1 S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA_X1 S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA_X1 S3_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\ab[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\CARRYB[9][10] ), .B(\ab[10][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\CARRYB[9][13] ), .B(\ab[10][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S2_10_14 ( .A(\CARRYB[9][14] ), .B(\ab[10][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S2_10_15 ( .A(\CARRYB[9][15] ), .B(\ab[10][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA_X1 S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA_X1 S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA_X1 S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA_X1 S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA_X1 S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA_X1 S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA_X1 S3_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\ab[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\CARRYB[8][11] ), .B(\ab[9][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\CARRYB[8][13] ), .B(\ab[9][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S2_9_15 ( .A(\CARRYB[8][15] ), .B(\ab[9][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA_X1 S2_9_16 ( .A(\CARRYB[8][16] ), .B(\ab[9][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA_X1 S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA_X1 S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA_X1 S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA_X1 S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA_X1 S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA_X1 S3_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\ab[8][23] ), .CO(
        \CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\CARRYB[7][12] ), .B(\ab[8][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\CARRYB[7][13] ), .B(\ab[8][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA_X1 S2_8_16 ( .A(\CARRYB[7][16] ), .B(\ab[8][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA_X1 S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA_X1 S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA_X1 S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA_X1 S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA_X1 S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA_X1 S3_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\ab[7][23] ), .CO(
        \CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\CARRYB[6][13] ), .B(\ab[7][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA_X1 S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA_X1 S2_7_17 ( .A(\CARRYB[6][17] ), .B(\ab[7][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA_X1 S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA_X1 S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA_X1 S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA_X1 S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA_X1 S3_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\ab[6][23] ), .CO(
        \CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\CARRYB[5][13] ), .B(\ab[6][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S2_6_14 ( .A(\CARRYB[5][14] ), .B(\ab[6][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_6_15 ( .A(\CARRYB[5][15] ), .B(\ab[6][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA_X1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA_X1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA_X1 S2_6_19 ( .A(\CARRYB[5][19] ), .B(\ab[6][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA_X1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA_X1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA_X1 S3_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\ab[5][23] ), .CO(
        \CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S2_5_15 ( .A(\CARRYB[4][15] ), .B(\ab[5][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA_X1 S2_5_16 ( .A(\CARRYB[4][16] ), .B(\ab[5][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA_X1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA_X1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA_X1 S2_5_19 ( .A(\CARRYB[4][19] ), .B(\ab[5][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA_X1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA_X1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA_X1 S3_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\ab[4][23] ), .CO(
        \CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA_X1 S2_4_16 ( .A(\CARRYB[3][16] ), .B(\ab[4][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA_X1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA_X1 S2_4_19 ( .A(\SUMB[3][20] ), .B(\ab[4][19] ), .CI(\CARRYB[3][19] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA_X1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA_X1 S2_4_21 ( .A(\SUMB[3][22] ), .B(\ab[4][21] ), .CI(\CARRYB[3][21] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA_X1 S3_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\ab[3][23] ), .CO(
        \CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA_X1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA_X1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA_X1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA_X1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA_X1 S2_3_20 ( .A(\CARRYB[2][20] ), .B(\ab[3][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n17), .CI(n26), .CO(\CARRYB[2][0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n9), .CI(n34), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n16), .CI(n25), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n8), .CI(n33), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n15), .CI(n24), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n7), .CI(n32), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n14), .CI(n23), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n6), .CI(n31), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n13), .CI(n22), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n5), .CI(n30), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n12), .CI(n21), .CO(\CARRYB[2][10] ), 
        .S(\SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n4), .CI(n29), .CO(\CARRYB[2][11] ), .S(
        \SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n11), .CI(n20), .CO(\CARRYB[2][12] ), 
        .S(\SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n3), .CI(n28), .CO(\CARRYB[2][13] ), .S(
        \SUMB[2][13] ) );
  FA_X1 S2_2_14 ( .A(\ab[2][14] ), .B(n10), .CI(n27), .CO(\CARRYB[2][14] ), 
        .S(\SUMB[2][14] ) );
  FA_X1 S2_2_15 ( .A(\ab[2][15] ), .B(n18), .CI(n42), .CO(\CARRYB[2][15] ), 
        .S(\SUMB[2][15] ) );
  FA_X1 S2_2_16 ( .A(\ab[2][16] ), .B(n39), .CI(n62), .CO(\CARRYB[2][16] ), 
        .S(\SUMB[2][16] ) );
  FA_X1 S2_2_17 ( .A(\ab[2][17] ), .B(n40), .CI(n79), .CO(\CARRYB[2][17] ), 
        .S(\SUMB[2][17] ) );
  FA_X1 S2_2_18 ( .A(\ab[2][18] ), .B(n19), .CI(n69), .CO(\CARRYB[2][18] ), 
        .S(\SUMB[2][18] ) );
  FA_X1 S2_2_20 ( .A(n86), .B(\ab[2][20] ), .CI(\CARRYB[1][20] ), .CO(
        \CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA_X1 S2_2_21 ( .A(\ab[2][21] ), .B(n88), .CI(\SUMB[1][22] ), .CO(
        \CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FP_MULTIPLIER_DW01_add_1 FS_1 ( .A({1'b0, n132, n90, n120, n99, n119, n98, 
        n112, n93, n111, n96, n118, n91, n113, n94, n114, n95, n115, n92, n116, 
        n97, n117, \A1[23] , n89, \SUMB[23][0] , \A1[20] , \A1[19] , \A1[18] , 
        \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , 
        \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , 
        \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\CARRYB[23][22] , n130, n110, 
        n129, n109, n128, n108, n122, n104, n121, n100, n127, n101, n123, n106, 
        n124, n105, n125, n102, n126, n107, \A2[24] , n103, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(
        PRODUCT[47:2]) );
  FA_X1 S0_20 ( .A(\ab[0][21] ), .B(1'b0), .CI(\ab[1][20] ), .CO(
        \CARRYB[1][20] ), .S(\SUMB[1][20] ) );
  FA_X1 S14_25 ( .A(1'b0), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), .CO(
        \A2[24] ), .S(\A1[23] ) );
  INV_X2 U2 ( .A(n83), .ZN(\CARRYB[1][22] ) );
  INV_X2 U3 ( .A(\ab[0][23] ), .ZN(n45) );
  NOR2_X1 U4 ( .A1(n154), .A2(n153), .ZN(\ab[2][22] ) );
  INV_X1 U5 ( .A(\ab[8][23] ), .ZN(n147) );
  INV_X1 U6 ( .A(\ab[9][23] ), .ZN(n146) );
  AND2_X1 U7 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n3) );
  AND2_X1 U8 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n4) );
  AND2_X1 U9 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n5) );
  AND2_X1 U10 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n6) );
  AND2_X1 U11 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n7) );
  AND2_X1 U12 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n8) );
  AND2_X1 U13 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n9) );
  AND2_X1 U14 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n10) );
  AND2_X1 U15 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n11) );
  AND2_X1 U16 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n12) );
  AND2_X1 U17 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n13) );
  AND2_X1 U18 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n14) );
  AND2_X1 U19 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n15) );
  AND2_X1 U20 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n16) );
  AND2_X1 U21 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n17) );
  AND2_X1 U22 ( .A1(\ab[0][16] ), .A2(\ab[1][15] ), .ZN(n18) );
  AND2_X1 U23 ( .A1(\ab[0][19] ), .A2(\ab[1][18] ), .ZN(n19) );
  XOR2_X1 U24 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n20) );
  XOR2_X1 U25 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n21) );
  XOR2_X1 U26 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n22) );
  XOR2_X1 U27 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n23) );
  XOR2_X1 U28 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n24) );
  XOR2_X1 U29 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n25) );
  XOR2_X1 U30 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n26) );
  XOR2_X1 U31 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(n27) );
  XOR2_X1 U32 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n28) );
  XOR2_X1 U33 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n29) );
  XOR2_X1 U34 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n30) );
  XOR2_X1 U35 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n31) );
  XOR2_X1 U36 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n32) );
  XOR2_X1 U37 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n33) );
  XOR2_X1 U38 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n34) );
  BUF_X1 U39 ( .A(n156), .Z(n65) );
  XOR2_X1 U40 ( .A(\ab[3][22] ), .B(\ab[2][23] ), .Z(n35) );
  XOR2_X1 U41 ( .A(\CARRYB[2][22] ), .B(n35), .Z(\SUMB[3][22] ) );
  NAND2_X1 U42 ( .A1(\CARRYB[2][22] ), .A2(\ab[3][22] ), .ZN(n36) );
  NAND2_X1 U43 ( .A1(\CARRYB[2][22] ), .A2(\ab[2][23] ), .ZN(n37) );
  NAND2_X1 U44 ( .A1(\ab[3][22] ), .A2(\ab[2][23] ), .ZN(n38) );
  NAND3_X1 U45 ( .A1(n36), .A2(n37), .A3(n38), .ZN(\CARRYB[3][22] ) );
  BUF_X1 U46 ( .A(n131), .Z(n73) );
  INV_X2 U47 ( .A(\ab[23][20] ), .ZN(n61) );
  AND2_X1 U48 ( .A1(\ab[1][23] ), .A2(\ab[23][20] ), .ZN(\ab[1][20] ) );
  AND2_X1 U49 ( .A1(\ab[1][23] ), .A2(\ab[23][21] ), .ZN(\ab[1][21] ) );
  AND2_X2 U50 ( .A1(\ab[1][23] ), .A2(\ab[23][22] ), .ZN(\ab[1][22] ) );
  AND2_X1 U51 ( .A1(\ab[0][17] ), .A2(\ab[1][16] ), .ZN(n39) );
  AND2_X1 U52 ( .A1(\ab[23][19] ), .A2(\ab[1][23] ), .ZN(\ab[1][19] ) );
  INV_X2 U53 ( .A(\ab[23][22] ), .ZN(n72) );
  INV_X1 U54 ( .A(\ab[1][23] ), .ZN(n68) );
  AND2_X1 U55 ( .A1(\ab[0][18] ), .A2(\ab[1][17] ), .ZN(n40) );
  INV_X4 U56 ( .A(\ab[23][16] ), .ZN(n158) );
  XNOR2_X1 U57 ( .A(n41), .B(\ab[0][18] ), .ZN(n62) );
  OR2_X1 U58 ( .A1(n46), .A2(n44), .ZN(n41) );
  AND2_X1 U59 ( .A1(\ab[0][23] ), .A2(\ab[23][21] ), .ZN(\ab[0][21] ) );
  CLKBUF_X1 U60 ( .A(n61), .Z(n84) );
  XOR2_X1 U61 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(n42) );
  XNOR2_X1 U62 ( .A(\SUMB[5][18] ), .B(n43), .ZN(\SUMB[6][17] ) );
  XNOR2_X1 U63 ( .A(\CARRYB[5][17] ), .B(\ab[6][17] ), .ZN(n43) );
  INV_X1 U64 ( .A(\ab[1][23] ), .ZN(n44) );
  XNOR2_X1 U65 ( .A(\ab[1][22] ), .B(n45), .ZN(\SUMB[1][22] ) );
  INV_X2 U66 ( .A(\ab[23][17] ), .ZN(n46) );
  INV_X2 U67 ( .A(\ab[23][17] ), .ZN(n47) );
  NAND2_X1 U68 ( .A1(\SUMB[5][18] ), .A2(\CARRYB[5][17] ), .ZN(n48) );
  NAND2_X1 U69 ( .A1(\SUMB[5][18] ), .A2(\ab[6][17] ), .ZN(n49) );
  NAND2_X1 U70 ( .A1(\CARRYB[5][17] ), .A2(\ab[6][17] ), .ZN(n50) );
  NAND3_X1 U71 ( .A1(n48), .A2(n49), .A3(n50), .ZN(\CARRYB[6][17] ) );
  XNOR2_X1 U72 ( .A(n51), .B(\SUMB[1][20] ), .ZN(\SUMB[2][19] ) );
  XNOR2_X1 U73 ( .A(n87), .B(\ab[2][19] ), .ZN(n51) );
  XNOR2_X1 U74 ( .A(\SUMB[3][19] ), .B(n52), .ZN(\SUMB[4][18] ) );
  XNOR2_X1 U75 ( .A(\CARRYB[3][18] ), .B(\ab[4][18] ), .ZN(n52) );
  NAND2_X1 U76 ( .A1(\SUMB[3][19] ), .A2(\CARRYB[3][18] ), .ZN(n53) );
  NAND2_X1 U77 ( .A1(\SUMB[3][19] ), .A2(\ab[4][18] ), .ZN(n54) );
  NAND2_X1 U78 ( .A1(\CARRYB[3][18] ), .A2(\ab[4][18] ), .ZN(n55) );
  NAND3_X1 U79 ( .A1(n53), .A2(n54), .A3(n55), .ZN(\CARRYB[4][18] ) );
  XOR2_X1 U80 ( .A(\ab[2][22] ), .B(\ab[1][23] ), .Z(n56) );
  XOR2_X1 U81 ( .A(\CARRYB[1][22] ), .B(n56), .Z(\SUMB[2][22] ) );
  NAND2_X1 U82 ( .A1(\CARRYB[1][22] ), .A2(\ab[2][22] ), .ZN(n57) );
  NAND2_X1 U83 ( .A1(\CARRYB[1][22] ), .A2(\ab[1][23] ), .ZN(n58) );
  NAND2_X1 U84 ( .A1(\ab[2][22] ), .A2(\ab[1][23] ), .ZN(n59) );
  NAND3_X1 U85 ( .A1(n57), .A2(n58), .A3(n59), .ZN(\CARRYB[2][22] ) );
  INV_X1 U86 ( .A(\ab[23][21] ), .ZN(n60) );
  CLKBUF_X1 U87 ( .A(n157), .Z(n63) );
  INV_X1 U88 ( .A(\ab[23][18] ), .ZN(n157) );
  INV_X2 U89 ( .A(\ab[2][23] ), .ZN(n64) );
  INV_X1 U90 ( .A(\ab[2][23] ), .ZN(n153) );
  AND2_X1 U91 ( .A1(\ab[23][19] ), .A2(\ab[0][23] ), .ZN(\ab[0][19] ) );
  INV_X1 U92 ( .A(\ab[23][19] ), .ZN(n156) );
  INV_X1 U93 ( .A(\ab[0][23] ), .ZN(n66) );
  INV_X1 U94 ( .A(\ab[0][23] ), .ZN(n67) );
  AND2_X1 U95 ( .A1(\ab[0][23] ), .A2(\ab[23][22] ), .ZN(\ab[0][22] ) );
  XOR2_X1 U96 ( .A(\ab[0][20] ), .B(\ab[1][19] ), .Z(n69) );
  BUF_X1 U97 ( .A(n87), .Z(n70) );
  AND2_X1 U98 ( .A1(\ab[0][20] ), .A2(\ab[1][19] ), .ZN(n87) );
  XNOR2_X1 U99 ( .A(\SUMB[2][22] ), .B(n71), .ZN(\SUMB[3][21] ) );
  XNOR2_X1 U100 ( .A(\CARRYB[2][21] ), .B(\ab[3][21] ), .ZN(n71) );
  BUF_X1 U101 ( .A(n60), .Z(n131) );
  NAND2_X1 U102 ( .A1(\SUMB[2][22] ), .A2(\CARRYB[2][21] ), .ZN(n74) );
  NAND2_X1 U103 ( .A1(\SUMB[2][22] ), .A2(\ab[3][21] ), .ZN(n75) );
  NAND2_X1 U104 ( .A1(\CARRYB[2][21] ), .A2(\ab[3][21] ), .ZN(n76) );
  NAND3_X1 U105 ( .A1(n74), .A2(n75), .A3(n76), .ZN(\CARRYB[3][21] ) );
  INV_X1 U106 ( .A(\ab[0][23] ), .ZN(n77) );
  INV_X1 U107 ( .A(\ab[0][23] ), .ZN(n78) );
  XOR2_X1 U108 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(n79) );
  NAND2_X1 U109 ( .A1(\SUMB[1][20] ), .A2(n70), .ZN(n80) );
  NAND2_X1 U110 ( .A1(\SUMB[1][20] ), .A2(\ab[2][19] ), .ZN(n81) );
  NAND2_X1 U111 ( .A1(n70), .A2(\ab[2][19] ), .ZN(n82) );
  NAND3_X1 U112 ( .A1(n80), .A2(n81), .A3(n82), .ZN(\CARRYB[2][19] ) );
  NAND2_X1 U113 ( .A1(\ab[1][22] ), .A2(\ab[0][23] ), .ZN(n83) );
  INV_X1 U114 ( .A(\ab[23][20] ), .ZN(n155) );
  INV_X4 U115 ( .A(\ab[23][11] ), .ZN(n163) );
  INV_X4 U116 ( .A(\ab[23][13] ), .ZN(n161) );
  INV_X4 U117 ( .A(\ab[23][9] ), .ZN(n165) );
  INV_X4 U118 ( .A(\ab[23][7] ), .ZN(n167) );
  INV_X4 U119 ( .A(\ab[23][5] ), .ZN(n169) );
  INV_X4 U120 ( .A(\ab[23][15] ), .ZN(n159) );
  INV_X4 U121 ( .A(\ab[23][3] ), .ZN(n171) );
  XOR2_X1 U122 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  XOR2_X1 U123 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(n86) );
  AND2_X1 U124 ( .A1(\ab[1][21] ), .A2(\ab[0][22] ), .ZN(n88) );
  XOR2_X1 U125 ( .A(\CARRYB[23][0] ), .B(\SUMB[23][1] ), .Z(n89) );
  INV_X1 U126 ( .A(\CARRYB[23][22] ), .ZN(n132) );
  XOR2_X1 U127 ( .A(\CARRYB[23][21] ), .B(\SUMB[23][22] ), .Z(n90) );
  XOR2_X1 U128 ( .A(\CARRYB[23][11] ), .B(\SUMB[23][12] ), .Z(n91) );
  XOR2_X1 U129 ( .A(\CARRYB[23][5] ), .B(\SUMB[23][6] ), .Z(n92) );
  XOR2_X1 U130 ( .A(\CARRYB[23][15] ), .B(\SUMB[23][16] ), .Z(n93) );
  XOR2_X1 U131 ( .A(\CARRYB[23][9] ), .B(\SUMB[23][10] ), .Z(n94) );
  XOR2_X1 U132 ( .A(\CARRYB[23][7] ), .B(\SUMB[23][8] ), .Z(n95) );
  XOR2_X1 U133 ( .A(\CARRYB[23][13] ), .B(\SUMB[23][14] ), .Z(n96) );
  XOR2_X1 U134 ( .A(\CARRYB[23][3] ), .B(\SUMB[23][4] ), .Z(n97) );
  XOR2_X1 U135 ( .A(\CARRYB[23][17] ), .B(\SUMB[23][18] ), .Z(n98) );
  XOR2_X1 U136 ( .A(\CARRYB[23][19] ), .B(\SUMB[23][20] ), .Z(n99) );
  AND2_X1 U137 ( .A1(\CARRYB[23][12] ), .A2(\SUMB[23][13] ), .ZN(n100) );
  AND2_X1 U138 ( .A1(\CARRYB[23][10] ), .A2(\SUMB[23][11] ), .ZN(n101) );
  AND2_X1 U139 ( .A1(\CARRYB[23][4] ), .A2(\SUMB[23][5] ), .ZN(n102) );
  AND2_X1 U140 ( .A1(\CARRYB[23][0] ), .A2(\SUMB[23][1] ), .ZN(n103) );
  AND2_X1 U141 ( .A1(\CARRYB[23][14] ), .A2(\SUMB[23][15] ), .ZN(n104) );
  AND2_X1 U142 ( .A1(\CARRYB[23][6] ), .A2(\SUMB[23][7] ), .ZN(n105) );
  AND2_X1 U143 ( .A1(\CARRYB[23][8] ), .A2(\SUMB[23][9] ), .ZN(n106) );
  AND2_X1 U144 ( .A1(\CARRYB[23][2] ), .A2(\SUMB[23][3] ), .ZN(n107) );
  AND2_X1 U145 ( .A1(\CARRYB[23][16] ), .A2(\SUMB[23][17] ), .ZN(n108) );
  AND2_X1 U146 ( .A1(\CARRYB[23][18] ), .A2(\SUMB[23][19] ), .ZN(n109) );
  AND2_X1 U147 ( .A1(\CARRYB[23][20] ), .A2(\SUMB[23][21] ), .ZN(n110) );
  XOR2_X1 U148 ( .A(\CARRYB[23][14] ), .B(\SUMB[23][15] ), .Z(n111) );
  XOR2_X1 U149 ( .A(\CARRYB[23][16] ), .B(\SUMB[23][17] ), .Z(n112) );
  XOR2_X1 U150 ( .A(\CARRYB[23][10] ), .B(\SUMB[23][11] ), .Z(n113) );
  XOR2_X1 U151 ( .A(\CARRYB[23][8] ), .B(\SUMB[23][9] ), .Z(n114) );
  XOR2_X1 U152 ( .A(\CARRYB[23][6] ), .B(\SUMB[23][7] ), .Z(n115) );
  XOR2_X1 U153 ( .A(\CARRYB[23][4] ), .B(\SUMB[23][5] ), .Z(n116) );
  XOR2_X1 U154 ( .A(\CARRYB[23][2] ), .B(\SUMB[23][3] ), .Z(n117) );
  XOR2_X1 U155 ( .A(\CARRYB[23][12] ), .B(\SUMB[23][13] ), .Z(n118) );
  XOR2_X1 U156 ( .A(\CARRYB[23][18] ), .B(\SUMB[23][19] ), .Z(n119) );
  XOR2_X1 U157 ( .A(\CARRYB[23][20] ), .B(\SUMB[23][21] ), .Z(n120) );
  AND2_X1 U158 ( .A1(\CARRYB[23][13] ), .A2(\SUMB[23][14] ), .ZN(n121) );
  AND2_X1 U159 ( .A1(\CARRYB[23][15] ), .A2(\SUMB[23][16] ), .ZN(n122) );
  AND2_X1 U160 ( .A1(\CARRYB[23][9] ), .A2(\SUMB[23][10] ), .ZN(n123) );
  AND2_X1 U161 ( .A1(\CARRYB[23][7] ), .A2(\SUMB[23][8] ), .ZN(n124) );
  AND2_X1 U162 ( .A1(\CARRYB[23][5] ), .A2(\SUMB[23][6] ), .ZN(n125) );
  AND2_X1 U163 ( .A1(\CARRYB[23][3] ), .A2(\SUMB[23][4] ), .ZN(n126) );
  AND2_X1 U164 ( .A1(\CARRYB[23][11] ), .A2(\SUMB[23][12] ), .ZN(n127) );
  AND2_X1 U165 ( .A1(\CARRYB[23][17] ), .A2(\SUMB[23][18] ), .ZN(n128) );
  AND2_X1 U166 ( .A1(\CARRYB[23][19] ), .A2(\SUMB[23][20] ), .ZN(n129) );
  AND2_X1 U167 ( .A1(\CARRYB[23][21] ), .A2(\SUMB[23][22] ), .ZN(n130) );
  INV_X2 U168 ( .A(\ab[23][10] ), .ZN(n164) );
  INV_X2 U169 ( .A(\ab[23][12] ), .ZN(n162) );
  INV_X2 U170 ( .A(\ab[23][8] ), .ZN(n166) );
  INV_X2 U171 ( .A(\ab[23][6] ), .ZN(n168) );
  INV_X2 U172 ( .A(\ab[23][4] ), .ZN(n170) );
  INV_X2 U173 ( .A(\ab[23][14] ), .ZN(n160) );
  INV_X2 U174 ( .A(\ab[23][2] ), .ZN(n172) );
  INV_X2 U175 ( .A(\ab[23][0] ), .ZN(n174) );
  INV_X2 U176 ( .A(\ab[3][23] ), .ZN(n152) );
  INV_X2 U177 ( .A(\ab[4][23] ), .ZN(n151) );
  INV_X2 U178 ( .A(\ab[5][23] ), .ZN(n150) );
  INV_X2 U179 ( .A(\ab[6][23] ), .ZN(n149) );
  INV_X2 U180 ( .A(\ab[7][23] ), .ZN(n148) );
  INV_X1 U181 ( .A(\ab[10][23] ), .ZN(n145) );
  INV_X1 U182 ( .A(\ab[11][23] ), .ZN(n144) );
  INV_X1 U183 ( .A(\ab[12][23] ), .ZN(n143) );
  INV_X1 U184 ( .A(\ab[13][23] ), .ZN(n142) );
  INV_X1 U185 ( .A(\ab[14][23] ), .ZN(n141) );
  INV_X1 U186 ( .A(\ab[15][23] ), .ZN(n140) );
  INV_X1 U187 ( .A(\ab[16][23] ), .ZN(n139) );
  INV_X1 U188 ( .A(\ab[17][23] ), .ZN(n138) );
  INV_X1 U189 ( .A(\ab[18][23] ), .ZN(n137) );
  INV_X1 U190 ( .A(\ab[19][23] ), .ZN(n136) );
  INV_X1 U191 ( .A(\ab[20][23] ), .ZN(n135) );
  INV_X1 U192 ( .A(\ab[21][23] ), .ZN(n134) );
  INV_X1 U193 ( .A(\ab[22][23] ), .ZN(n133) );
  INV_X1 U194 ( .A(\ab[23][22] ), .ZN(n154) );
  INV_X4 U195 ( .A(\ab[23][1] ), .ZN(n173) );
  NOR2_X1 U197 ( .A1(n146), .A2(n165), .ZN(\ab[9][9] ) );
  NOR2_X1 U198 ( .A1(n146), .A2(n166), .ZN(\ab[9][8] ) );
  NOR2_X1 U199 ( .A1(n146), .A2(n167), .ZN(\ab[9][7] ) );
  NOR2_X1 U200 ( .A1(n146), .A2(n168), .ZN(\ab[9][6] ) );
  NOR2_X1 U201 ( .A1(n146), .A2(n169), .ZN(\ab[9][5] ) );
  NOR2_X1 U202 ( .A1(n146), .A2(n170), .ZN(\ab[9][4] ) );
  NOR2_X1 U203 ( .A1(n146), .A2(n171), .ZN(\ab[9][3] ) );
  NOR2_X1 U204 ( .A1(n146), .A2(n172), .ZN(\ab[9][2] ) );
  NOR2_X1 U205 ( .A1(n146), .A2(n72), .ZN(\ab[9][22] ) );
  NOR2_X1 U206 ( .A1(n146), .A2(n73), .ZN(\ab[9][21] ) );
  NOR2_X1 U207 ( .A1(n146), .A2(n61), .ZN(\ab[9][20] ) );
  NOR2_X1 U208 ( .A1(n146), .A2(n173), .ZN(\ab[9][1] ) );
  NOR2_X1 U209 ( .A1(n146), .A2(n65), .ZN(\ab[9][19] ) );
  NOR2_X1 U210 ( .A1(n146), .A2(n63), .ZN(\ab[9][18] ) );
  NOR2_X1 U211 ( .A1(n146), .A2(n47), .ZN(\ab[9][17] ) );
  NOR2_X1 U212 ( .A1(n146), .A2(n158), .ZN(\ab[9][16] ) );
  NOR2_X1 U213 ( .A1(n146), .A2(n159), .ZN(\ab[9][15] ) );
  NOR2_X1 U214 ( .A1(n146), .A2(n160), .ZN(\ab[9][14] ) );
  NOR2_X1 U215 ( .A1(n146), .A2(n161), .ZN(\ab[9][13] ) );
  NOR2_X1 U216 ( .A1(n146), .A2(n162), .ZN(\ab[9][12] ) );
  NOR2_X1 U217 ( .A1(n146), .A2(n163), .ZN(\ab[9][11] ) );
  NOR2_X1 U218 ( .A1(n146), .A2(n164), .ZN(\ab[9][10] ) );
  NOR2_X1 U219 ( .A1(n146), .A2(n174), .ZN(\ab[9][0] ) );
  NOR2_X1 U220 ( .A1(n165), .A2(n147), .ZN(\ab[8][9] ) );
  NOR2_X1 U221 ( .A1(n166), .A2(n147), .ZN(\ab[8][8] ) );
  NOR2_X1 U222 ( .A1(n167), .A2(n147), .ZN(\ab[8][7] ) );
  NOR2_X1 U223 ( .A1(n168), .A2(n147), .ZN(\ab[8][6] ) );
  NOR2_X1 U224 ( .A1(n169), .A2(n147), .ZN(\ab[8][5] ) );
  NOR2_X1 U225 ( .A1(n170), .A2(n147), .ZN(\ab[8][4] ) );
  NOR2_X1 U226 ( .A1(n171), .A2(n147), .ZN(\ab[8][3] ) );
  NOR2_X1 U227 ( .A1(n172), .A2(n147), .ZN(\ab[8][2] ) );
  NOR2_X1 U228 ( .A1(n147), .A2(n72), .ZN(\ab[8][22] ) );
  NOR2_X1 U229 ( .A1(n73), .A2(n147), .ZN(\ab[8][21] ) );
  NOR2_X1 U230 ( .A1(n61), .A2(n147), .ZN(\ab[8][20] ) );
  NOR2_X1 U231 ( .A1(n173), .A2(n147), .ZN(\ab[8][1] ) );
  NOR2_X1 U232 ( .A1(n65), .A2(n147), .ZN(\ab[8][19] ) );
  NOR2_X1 U233 ( .A1(n63), .A2(n147), .ZN(\ab[8][18] ) );
  NOR2_X1 U234 ( .A1(n47), .A2(n147), .ZN(\ab[8][17] ) );
  NOR2_X1 U235 ( .A1(n158), .A2(n147), .ZN(\ab[8][16] ) );
  NOR2_X1 U236 ( .A1(n159), .A2(n147), .ZN(\ab[8][15] ) );
  NOR2_X1 U237 ( .A1(n160), .A2(n147), .ZN(\ab[8][14] ) );
  NOR2_X1 U238 ( .A1(n161), .A2(n147), .ZN(\ab[8][13] ) );
  NOR2_X1 U239 ( .A1(n162), .A2(n147), .ZN(\ab[8][12] ) );
  NOR2_X1 U240 ( .A1(n163), .A2(n147), .ZN(\ab[8][11] ) );
  NOR2_X1 U241 ( .A1(n164), .A2(n147), .ZN(\ab[8][10] ) );
  NOR2_X1 U242 ( .A1(n174), .A2(n147), .ZN(\ab[8][0] ) );
  NOR2_X1 U243 ( .A1(n165), .A2(n148), .ZN(\ab[7][9] ) );
  NOR2_X1 U244 ( .A1(n166), .A2(n148), .ZN(\ab[7][8] ) );
  NOR2_X1 U245 ( .A1(n167), .A2(n148), .ZN(\ab[7][7] ) );
  NOR2_X1 U246 ( .A1(n168), .A2(n148), .ZN(\ab[7][6] ) );
  NOR2_X1 U247 ( .A1(n169), .A2(n148), .ZN(\ab[7][5] ) );
  NOR2_X1 U248 ( .A1(n170), .A2(n148), .ZN(\ab[7][4] ) );
  NOR2_X1 U249 ( .A1(n171), .A2(n148), .ZN(\ab[7][3] ) );
  NOR2_X1 U250 ( .A1(n172), .A2(n148), .ZN(\ab[7][2] ) );
  NOR2_X1 U251 ( .A1(n72), .A2(n148), .ZN(\ab[7][22] ) );
  NOR2_X1 U252 ( .A1(n73), .A2(n148), .ZN(\ab[7][21] ) );
  NOR2_X1 U253 ( .A1(n61), .A2(n148), .ZN(\ab[7][20] ) );
  NOR2_X1 U254 ( .A1(n173), .A2(n148), .ZN(\ab[7][1] ) );
  NOR2_X1 U255 ( .A1(n65), .A2(n148), .ZN(\ab[7][19] ) );
  NOR2_X1 U256 ( .A1(n63), .A2(n148), .ZN(\ab[7][18] ) );
  NOR2_X1 U257 ( .A1(n46), .A2(n148), .ZN(\ab[7][17] ) );
  NOR2_X1 U258 ( .A1(n158), .A2(n148), .ZN(\ab[7][16] ) );
  NOR2_X1 U259 ( .A1(n159), .A2(n148), .ZN(\ab[7][15] ) );
  NOR2_X1 U260 ( .A1(n160), .A2(n148), .ZN(\ab[7][14] ) );
  NOR2_X1 U261 ( .A1(n161), .A2(n148), .ZN(\ab[7][13] ) );
  NOR2_X1 U262 ( .A1(n162), .A2(n148), .ZN(\ab[7][12] ) );
  NOR2_X1 U263 ( .A1(n163), .A2(n148), .ZN(\ab[7][11] ) );
  NOR2_X1 U264 ( .A1(n164), .A2(n148), .ZN(\ab[7][10] ) );
  NOR2_X1 U265 ( .A1(n174), .A2(n148), .ZN(\ab[7][0] ) );
  NOR2_X1 U266 ( .A1(n165), .A2(n149), .ZN(\ab[6][9] ) );
  NOR2_X1 U267 ( .A1(n166), .A2(n149), .ZN(\ab[6][8] ) );
  NOR2_X1 U268 ( .A1(n167), .A2(n149), .ZN(\ab[6][7] ) );
  NOR2_X1 U269 ( .A1(n168), .A2(n149), .ZN(\ab[6][6] ) );
  NOR2_X1 U270 ( .A1(n169), .A2(n149), .ZN(\ab[6][5] ) );
  NOR2_X1 U271 ( .A1(n170), .A2(n149), .ZN(\ab[6][4] ) );
  NOR2_X1 U272 ( .A1(n171), .A2(n149), .ZN(\ab[6][3] ) );
  NOR2_X1 U273 ( .A1(n172), .A2(n149), .ZN(\ab[6][2] ) );
  NOR2_X1 U274 ( .A1(n72), .A2(n149), .ZN(\ab[6][22] ) );
  NOR2_X1 U275 ( .A1(n73), .A2(n149), .ZN(\ab[6][21] ) );
  NOR2_X1 U276 ( .A1(n61), .A2(n149), .ZN(\ab[6][20] ) );
  NOR2_X1 U277 ( .A1(n173), .A2(n149), .ZN(\ab[6][1] ) );
  NOR2_X1 U278 ( .A1(n65), .A2(n149), .ZN(\ab[6][19] ) );
  NOR2_X1 U279 ( .A1(n63), .A2(n149), .ZN(\ab[6][18] ) );
  NOR2_X1 U280 ( .A1(n47), .A2(n149), .ZN(\ab[6][17] ) );
  NOR2_X1 U281 ( .A1(n158), .A2(n149), .ZN(\ab[6][16] ) );
  NOR2_X1 U282 ( .A1(n159), .A2(n149), .ZN(\ab[6][15] ) );
  NOR2_X1 U283 ( .A1(n160), .A2(n149), .ZN(\ab[6][14] ) );
  NOR2_X1 U284 ( .A1(n161), .A2(n149), .ZN(\ab[6][13] ) );
  NOR2_X1 U285 ( .A1(n162), .A2(n149), .ZN(\ab[6][12] ) );
  NOR2_X1 U286 ( .A1(n163), .A2(n149), .ZN(\ab[6][11] ) );
  NOR2_X1 U287 ( .A1(n164), .A2(n149), .ZN(\ab[6][10] ) );
  NOR2_X1 U288 ( .A1(n174), .A2(n149), .ZN(\ab[6][0] ) );
  NOR2_X1 U289 ( .A1(n165), .A2(n150), .ZN(\ab[5][9] ) );
  NOR2_X1 U290 ( .A1(n166), .A2(n150), .ZN(\ab[5][8] ) );
  NOR2_X1 U291 ( .A1(n167), .A2(n150), .ZN(\ab[5][7] ) );
  NOR2_X1 U292 ( .A1(n168), .A2(n150), .ZN(\ab[5][6] ) );
  NOR2_X1 U293 ( .A1(n169), .A2(n150), .ZN(\ab[5][5] ) );
  NOR2_X1 U294 ( .A1(n170), .A2(n150), .ZN(\ab[5][4] ) );
  NOR2_X1 U295 ( .A1(n171), .A2(n150), .ZN(\ab[5][3] ) );
  NOR2_X1 U296 ( .A1(n172), .A2(n150), .ZN(\ab[5][2] ) );
  NOR2_X1 U297 ( .A1(n72), .A2(n150), .ZN(\ab[5][22] ) );
  NOR2_X1 U298 ( .A1(n131), .A2(n150), .ZN(\ab[5][21] ) );
  NOR2_X1 U299 ( .A1(n61), .A2(n150), .ZN(\ab[5][20] ) );
  NOR2_X1 U300 ( .A1(n173), .A2(n150), .ZN(\ab[5][1] ) );
  NOR2_X1 U301 ( .A1(n156), .A2(n150), .ZN(\ab[5][19] ) );
  NOR2_X1 U302 ( .A1(n157), .A2(n150), .ZN(\ab[5][18] ) );
  NOR2_X1 U303 ( .A1(n47), .A2(n150), .ZN(\ab[5][17] ) );
  NOR2_X1 U304 ( .A1(n158), .A2(n150), .ZN(\ab[5][16] ) );
  NOR2_X1 U305 ( .A1(n159), .A2(n150), .ZN(\ab[5][15] ) );
  NOR2_X1 U306 ( .A1(n160), .A2(n150), .ZN(\ab[5][14] ) );
  NOR2_X1 U307 ( .A1(n161), .A2(n150), .ZN(\ab[5][13] ) );
  NOR2_X1 U308 ( .A1(n162), .A2(n150), .ZN(\ab[5][12] ) );
  NOR2_X1 U309 ( .A1(n163), .A2(n150), .ZN(\ab[5][11] ) );
  NOR2_X1 U310 ( .A1(n164), .A2(n150), .ZN(\ab[5][10] ) );
  NOR2_X1 U311 ( .A1(n174), .A2(n150), .ZN(\ab[5][0] ) );
  NOR2_X1 U312 ( .A1(n165), .A2(n151), .ZN(\ab[4][9] ) );
  NOR2_X1 U313 ( .A1(n166), .A2(n151), .ZN(\ab[4][8] ) );
  NOR2_X1 U314 ( .A1(n167), .A2(n151), .ZN(\ab[4][7] ) );
  NOR2_X1 U315 ( .A1(n168), .A2(n151), .ZN(\ab[4][6] ) );
  NOR2_X1 U316 ( .A1(n169), .A2(n151), .ZN(\ab[4][5] ) );
  NOR2_X1 U317 ( .A1(n170), .A2(n151), .ZN(\ab[4][4] ) );
  NOR2_X1 U318 ( .A1(n171), .A2(n151), .ZN(\ab[4][3] ) );
  NOR2_X1 U319 ( .A1(n172), .A2(n151), .ZN(\ab[4][2] ) );
  NOR2_X1 U320 ( .A1(n72), .A2(n151), .ZN(\ab[4][22] ) );
  NOR2_X1 U321 ( .A1(n131), .A2(n151), .ZN(\ab[4][21] ) );
  NOR2_X1 U322 ( .A1(n61), .A2(n151), .ZN(\ab[4][20] ) );
  NOR2_X1 U323 ( .A1(n173), .A2(n151), .ZN(\ab[4][1] ) );
  NOR2_X1 U324 ( .A1(n156), .A2(n151), .ZN(\ab[4][19] ) );
  NOR2_X1 U325 ( .A1(n157), .A2(n151), .ZN(\ab[4][18] ) );
  NOR2_X1 U326 ( .A1(n47), .A2(n151), .ZN(\ab[4][17] ) );
  NOR2_X1 U327 ( .A1(n158), .A2(n151), .ZN(\ab[4][16] ) );
  NOR2_X1 U328 ( .A1(n159), .A2(n151), .ZN(\ab[4][15] ) );
  NOR2_X1 U329 ( .A1(n160), .A2(n151), .ZN(\ab[4][14] ) );
  NOR2_X1 U330 ( .A1(n161), .A2(n151), .ZN(\ab[4][13] ) );
  NOR2_X1 U331 ( .A1(n162), .A2(n151), .ZN(\ab[4][12] ) );
  NOR2_X1 U332 ( .A1(n163), .A2(n151), .ZN(\ab[4][11] ) );
  NOR2_X1 U333 ( .A1(n164), .A2(n151), .ZN(\ab[4][10] ) );
  NOR2_X1 U334 ( .A1(n174), .A2(n151), .ZN(\ab[4][0] ) );
  NOR2_X1 U335 ( .A1(n165), .A2(n152), .ZN(\ab[3][9] ) );
  NOR2_X1 U336 ( .A1(n166), .A2(n152), .ZN(\ab[3][8] ) );
  NOR2_X1 U337 ( .A1(n167), .A2(n152), .ZN(\ab[3][7] ) );
  NOR2_X1 U338 ( .A1(n168), .A2(n152), .ZN(\ab[3][6] ) );
  NOR2_X1 U339 ( .A1(n169), .A2(n152), .ZN(\ab[3][5] ) );
  NOR2_X1 U340 ( .A1(n170), .A2(n152), .ZN(\ab[3][4] ) );
  NOR2_X1 U341 ( .A1(n171), .A2(n152), .ZN(\ab[3][3] ) );
  NOR2_X1 U342 ( .A1(n172), .A2(n152), .ZN(\ab[3][2] ) );
  NOR2_X1 U343 ( .A1(n72), .A2(n152), .ZN(\ab[3][22] ) );
  NOR2_X1 U344 ( .A1(n131), .A2(n152), .ZN(\ab[3][21] ) );
  NOR2_X1 U345 ( .A1(n61), .A2(n152), .ZN(\ab[3][20] ) );
  NOR2_X1 U346 ( .A1(n173), .A2(n152), .ZN(\ab[3][1] ) );
  NOR2_X1 U347 ( .A1(n156), .A2(n152), .ZN(\ab[3][19] ) );
  NOR2_X1 U348 ( .A1(n157), .A2(n152), .ZN(\ab[3][18] ) );
  NOR2_X1 U349 ( .A1(n46), .A2(n152), .ZN(\ab[3][17] ) );
  NOR2_X1 U350 ( .A1(n158), .A2(n152), .ZN(\ab[3][16] ) );
  NOR2_X1 U351 ( .A1(n159), .A2(n152), .ZN(\ab[3][15] ) );
  NOR2_X1 U352 ( .A1(n160), .A2(n152), .ZN(\ab[3][14] ) );
  NOR2_X1 U353 ( .A1(n161), .A2(n152), .ZN(\ab[3][13] ) );
  NOR2_X1 U354 ( .A1(n162), .A2(n152), .ZN(\ab[3][12] ) );
  NOR2_X1 U355 ( .A1(n163), .A2(n152), .ZN(\ab[3][11] ) );
  NOR2_X1 U356 ( .A1(n164), .A2(n152), .ZN(\ab[3][10] ) );
  NOR2_X1 U357 ( .A1(n174), .A2(n152), .ZN(\ab[3][0] ) );
  NOR2_X1 U358 ( .A1(n165), .A2(n64), .ZN(\ab[2][9] ) );
  NOR2_X1 U359 ( .A1(n166), .A2(n64), .ZN(\ab[2][8] ) );
  NOR2_X1 U360 ( .A1(n167), .A2(n64), .ZN(\ab[2][7] ) );
  NOR2_X1 U361 ( .A1(n168), .A2(n64), .ZN(\ab[2][6] ) );
  NOR2_X1 U362 ( .A1(n169), .A2(n64), .ZN(\ab[2][5] ) );
  NOR2_X1 U363 ( .A1(n170), .A2(n64), .ZN(\ab[2][4] ) );
  NOR2_X1 U364 ( .A1(n171), .A2(n64), .ZN(\ab[2][3] ) );
  NOR2_X1 U365 ( .A1(n172), .A2(n64), .ZN(\ab[2][2] ) );
  NOR2_X1 U366 ( .A1(n60), .A2(n153), .ZN(\ab[2][21] ) );
  NOR2_X1 U367 ( .A1(n155), .A2(n153), .ZN(\ab[2][20] ) );
  NOR2_X1 U368 ( .A1(n173), .A2(n64), .ZN(\ab[2][1] ) );
  NOR2_X1 U369 ( .A1(n156), .A2(n153), .ZN(\ab[2][19] ) );
  NOR2_X1 U370 ( .A1(n157), .A2(n64), .ZN(\ab[2][18] ) );
  NOR2_X1 U371 ( .A1(n46), .A2(n64), .ZN(\ab[2][17] ) );
  NOR2_X1 U372 ( .A1(n158), .A2(n64), .ZN(\ab[2][16] ) );
  NOR2_X1 U373 ( .A1(n159), .A2(n64), .ZN(\ab[2][15] ) );
  NOR2_X1 U374 ( .A1(n160), .A2(n64), .ZN(\ab[2][14] ) );
  NOR2_X1 U375 ( .A1(n161), .A2(n64), .ZN(\ab[2][13] ) );
  NOR2_X1 U376 ( .A1(n162), .A2(n64), .ZN(\ab[2][12] ) );
  NOR2_X1 U377 ( .A1(n163), .A2(n64), .ZN(\ab[2][11] ) );
  NOR2_X1 U378 ( .A1(n164), .A2(n64), .ZN(\ab[2][10] ) );
  NOR2_X1 U379 ( .A1(n174), .A2(n64), .ZN(\ab[2][0] ) );
  NOR2_X1 U380 ( .A1(n165), .A2(n133), .ZN(\ab[22][9] ) );
  NOR2_X1 U381 ( .A1(n166), .A2(n133), .ZN(\ab[22][8] ) );
  NOR2_X1 U382 ( .A1(n167), .A2(n133), .ZN(\ab[22][7] ) );
  NOR2_X1 U383 ( .A1(n168), .A2(n133), .ZN(\ab[22][6] ) );
  NOR2_X1 U384 ( .A1(n169), .A2(n133), .ZN(\ab[22][5] ) );
  NOR2_X1 U385 ( .A1(n170), .A2(n133), .ZN(\ab[22][4] ) );
  NOR2_X1 U386 ( .A1(n171), .A2(n133), .ZN(\ab[22][3] ) );
  NOR2_X1 U387 ( .A1(n172), .A2(n133), .ZN(\ab[22][2] ) );
  NOR2_X1 U388 ( .A1(n72), .A2(n133), .ZN(\ab[22][22] ) );
  NOR2_X1 U389 ( .A1(n73), .A2(n133), .ZN(\ab[22][21] ) );
  NOR2_X1 U390 ( .A1(n84), .A2(n133), .ZN(\ab[22][20] ) );
  NOR2_X1 U391 ( .A1(n173), .A2(n133), .ZN(\ab[22][1] ) );
  NOR2_X1 U392 ( .A1(n65), .A2(n133), .ZN(\ab[22][19] ) );
  NOR2_X1 U393 ( .A1(n63), .A2(n133), .ZN(\ab[22][18] ) );
  NOR2_X1 U394 ( .A1(n46), .A2(n133), .ZN(\ab[22][17] ) );
  NOR2_X1 U395 ( .A1(n158), .A2(n133), .ZN(\ab[22][16] ) );
  NOR2_X1 U396 ( .A1(n159), .A2(n133), .ZN(\ab[22][15] ) );
  NOR2_X1 U397 ( .A1(n160), .A2(n133), .ZN(\ab[22][14] ) );
  NOR2_X1 U398 ( .A1(n161), .A2(n133), .ZN(\ab[22][13] ) );
  NOR2_X1 U399 ( .A1(n162), .A2(n133), .ZN(\ab[22][12] ) );
  NOR2_X1 U400 ( .A1(n163), .A2(n133), .ZN(\ab[22][11] ) );
  NOR2_X1 U401 ( .A1(n164), .A2(n133), .ZN(\ab[22][10] ) );
  NOR2_X1 U402 ( .A1(n174), .A2(n133), .ZN(\ab[22][0] ) );
  NOR2_X1 U403 ( .A1(n165), .A2(n134), .ZN(\ab[21][9] ) );
  NOR2_X1 U404 ( .A1(n166), .A2(n134), .ZN(\ab[21][8] ) );
  NOR2_X1 U405 ( .A1(n167), .A2(n134), .ZN(\ab[21][7] ) );
  NOR2_X1 U406 ( .A1(n168), .A2(n134), .ZN(\ab[21][6] ) );
  NOR2_X1 U407 ( .A1(n169), .A2(n134), .ZN(\ab[21][5] ) );
  NOR2_X1 U408 ( .A1(n170), .A2(n134), .ZN(\ab[21][4] ) );
  NOR2_X1 U409 ( .A1(n171), .A2(n134), .ZN(\ab[21][3] ) );
  NOR2_X1 U410 ( .A1(n172), .A2(n134), .ZN(\ab[21][2] ) );
  NOR2_X1 U411 ( .A1(n72), .A2(n134), .ZN(\ab[21][22] ) );
  NOR2_X1 U412 ( .A1(n73), .A2(n134), .ZN(\ab[21][21] ) );
  NOR2_X1 U413 ( .A1(n84), .A2(n134), .ZN(\ab[21][20] ) );
  NOR2_X1 U414 ( .A1(n173), .A2(n134), .ZN(\ab[21][1] ) );
  NOR2_X1 U415 ( .A1(n65), .A2(n134), .ZN(\ab[21][19] ) );
  NOR2_X1 U416 ( .A1(n63), .A2(n134), .ZN(\ab[21][18] ) );
  NOR2_X1 U417 ( .A1(n47), .A2(n134), .ZN(\ab[21][17] ) );
  NOR2_X1 U418 ( .A1(n158), .A2(n134), .ZN(\ab[21][16] ) );
  NOR2_X1 U419 ( .A1(n159), .A2(n134), .ZN(\ab[21][15] ) );
  NOR2_X1 U420 ( .A1(n160), .A2(n134), .ZN(\ab[21][14] ) );
  NOR2_X1 U421 ( .A1(n161), .A2(n134), .ZN(\ab[21][13] ) );
  NOR2_X1 U422 ( .A1(n162), .A2(n134), .ZN(\ab[21][12] ) );
  NOR2_X1 U423 ( .A1(n163), .A2(n134), .ZN(\ab[21][11] ) );
  NOR2_X1 U424 ( .A1(n164), .A2(n134), .ZN(\ab[21][10] ) );
  NOR2_X1 U425 ( .A1(n174), .A2(n134), .ZN(\ab[21][0] ) );
  NOR2_X1 U426 ( .A1(n165), .A2(n135), .ZN(\ab[20][9] ) );
  NOR2_X1 U427 ( .A1(n166), .A2(n135), .ZN(\ab[20][8] ) );
  NOR2_X1 U428 ( .A1(n167), .A2(n135), .ZN(\ab[20][7] ) );
  NOR2_X1 U429 ( .A1(n168), .A2(n135), .ZN(\ab[20][6] ) );
  NOR2_X1 U430 ( .A1(n169), .A2(n135), .ZN(\ab[20][5] ) );
  NOR2_X1 U431 ( .A1(n170), .A2(n135), .ZN(\ab[20][4] ) );
  NOR2_X1 U432 ( .A1(n171), .A2(n135), .ZN(\ab[20][3] ) );
  NOR2_X1 U433 ( .A1(n172), .A2(n135), .ZN(\ab[20][2] ) );
  NOR2_X1 U434 ( .A1(n72), .A2(n135), .ZN(\ab[20][22] ) );
  NOR2_X1 U435 ( .A1(n73), .A2(n135), .ZN(\ab[20][21] ) );
  NOR2_X1 U436 ( .A1(n84), .A2(n135), .ZN(\ab[20][20] ) );
  NOR2_X1 U437 ( .A1(n173), .A2(n135), .ZN(\ab[20][1] ) );
  NOR2_X1 U438 ( .A1(n65), .A2(n135), .ZN(\ab[20][19] ) );
  NOR2_X1 U439 ( .A1(n63), .A2(n135), .ZN(\ab[20][18] ) );
  NOR2_X1 U440 ( .A1(n46), .A2(n135), .ZN(\ab[20][17] ) );
  NOR2_X1 U441 ( .A1(n158), .A2(n135), .ZN(\ab[20][16] ) );
  NOR2_X1 U442 ( .A1(n159), .A2(n135), .ZN(\ab[20][15] ) );
  NOR2_X1 U443 ( .A1(n160), .A2(n135), .ZN(\ab[20][14] ) );
  NOR2_X1 U444 ( .A1(n161), .A2(n135), .ZN(\ab[20][13] ) );
  NOR2_X1 U445 ( .A1(n162), .A2(n135), .ZN(\ab[20][12] ) );
  NOR2_X1 U446 ( .A1(n163), .A2(n135), .ZN(\ab[20][11] ) );
  NOR2_X1 U447 ( .A1(n164), .A2(n135), .ZN(\ab[20][10] ) );
  NOR2_X1 U448 ( .A1(n174), .A2(n135), .ZN(\ab[20][0] ) );
  NOR2_X1 U449 ( .A1(n165), .A2(n68), .ZN(\ab[1][9] ) );
  NOR2_X1 U450 ( .A1(n166), .A2(n44), .ZN(\ab[1][8] ) );
  NOR2_X1 U451 ( .A1(n167), .A2(n44), .ZN(\ab[1][7] ) );
  NOR2_X1 U452 ( .A1(n168), .A2(n44), .ZN(\ab[1][6] ) );
  NOR2_X1 U453 ( .A1(n169), .A2(n68), .ZN(\ab[1][5] ) );
  NOR2_X1 U454 ( .A1(n170), .A2(n44), .ZN(\ab[1][4] ) );
  NOR2_X1 U455 ( .A1(n171), .A2(n68), .ZN(\ab[1][3] ) );
  NOR2_X1 U456 ( .A1(n172), .A2(n44), .ZN(\ab[1][2] ) );
  NOR2_X1 U457 ( .A1(n173), .A2(n68), .ZN(\ab[1][1] ) );
  NOR2_X1 U458 ( .A1(n157), .A2(n68), .ZN(\ab[1][18] ) );
  NOR2_X1 U459 ( .A1(n47), .A2(n68), .ZN(\ab[1][17] ) );
  NOR2_X1 U460 ( .A1(n158), .A2(n44), .ZN(\ab[1][16] ) );
  NOR2_X1 U461 ( .A1(n159), .A2(n44), .ZN(\ab[1][15] ) );
  NOR2_X1 U462 ( .A1(n160), .A2(n44), .ZN(\ab[1][14] ) );
  NOR2_X1 U463 ( .A1(n161), .A2(n68), .ZN(\ab[1][13] ) );
  NOR2_X1 U464 ( .A1(n162), .A2(n44), .ZN(\ab[1][12] ) );
  NOR2_X1 U465 ( .A1(n163), .A2(n68), .ZN(\ab[1][11] ) );
  NOR2_X1 U466 ( .A1(n164), .A2(n44), .ZN(\ab[1][10] ) );
  NOR2_X1 U467 ( .A1(n174), .A2(n44), .ZN(\ab[1][0] ) );
  NOR2_X1 U468 ( .A1(n165), .A2(n136), .ZN(\ab[19][9] ) );
  NOR2_X1 U469 ( .A1(n166), .A2(n136), .ZN(\ab[19][8] ) );
  NOR2_X1 U470 ( .A1(n167), .A2(n136), .ZN(\ab[19][7] ) );
  NOR2_X1 U471 ( .A1(n168), .A2(n136), .ZN(\ab[19][6] ) );
  NOR2_X1 U472 ( .A1(n169), .A2(n136), .ZN(\ab[19][5] ) );
  NOR2_X1 U473 ( .A1(n170), .A2(n136), .ZN(\ab[19][4] ) );
  NOR2_X1 U474 ( .A1(n171), .A2(n136), .ZN(\ab[19][3] ) );
  NOR2_X1 U475 ( .A1(n172), .A2(n136), .ZN(\ab[19][2] ) );
  NOR2_X1 U476 ( .A1(n72), .A2(n136), .ZN(\ab[19][22] ) );
  NOR2_X1 U477 ( .A1(n73), .A2(n136), .ZN(\ab[19][21] ) );
  NOR2_X1 U478 ( .A1(n61), .A2(n136), .ZN(\ab[19][20] ) );
  NOR2_X1 U479 ( .A1(n173), .A2(n136), .ZN(\ab[19][1] ) );
  NOR2_X1 U480 ( .A1(n65), .A2(n136), .ZN(\ab[19][19] ) );
  NOR2_X1 U481 ( .A1(n63), .A2(n136), .ZN(\ab[19][18] ) );
  NOR2_X1 U482 ( .A1(n47), .A2(n136), .ZN(\ab[19][17] ) );
  NOR2_X1 U483 ( .A1(n158), .A2(n136), .ZN(\ab[19][16] ) );
  NOR2_X1 U484 ( .A1(n159), .A2(n136), .ZN(\ab[19][15] ) );
  NOR2_X1 U485 ( .A1(n160), .A2(n136), .ZN(\ab[19][14] ) );
  NOR2_X1 U486 ( .A1(n161), .A2(n136), .ZN(\ab[19][13] ) );
  NOR2_X1 U487 ( .A1(n162), .A2(n136), .ZN(\ab[19][12] ) );
  NOR2_X1 U488 ( .A1(n163), .A2(n136), .ZN(\ab[19][11] ) );
  NOR2_X1 U489 ( .A1(n164), .A2(n136), .ZN(\ab[19][10] ) );
  NOR2_X1 U490 ( .A1(n174), .A2(n136), .ZN(\ab[19][0] ) );
  NOR2_X1 U491 ( .A1(n165), .A2(n137), .ZN(\ab[18][9] ) );
  NOR2_X1 U492 ( .A1(n166), .A2(n137), .ZN(\ab[18][8] ) );
  NOR2_X1 U493 ( .A1(n167), .A2(n137), .ZN(\ab[18][7] ) );
  NOR2_X1 U494 ( .A1(n168), .A2(n137), .ZN(\ab[18][6] ) );
  NOR2_X1 U495 ( .A1(n169), .A2(n137), .ZN(\ab[18][5] ) );
  NOR2_X1 U496 ( .A1(n170), .A2(n137), .ZN(\ab[18][4] ) );
  NOR2_X1 U497 ( .A1(n171), .A2(n137), .ZN(\ab[18][3] ) );
  NOR2_X1 U498 ( .A1(n172), .A2(n137), .ZN(\ab[18][2] ) );
  NOR2_X1 U499 ( .A1(n72), .A2(n137), .ZN(\ab[18][22] ) );
  NOR2_X1 U500 ( .A1(n73), .A2(n137), .ZN(\ab[18][21] ) );
  NOR2_X1 U501 ( .A1(n61), .A2(n137), .ZN(\ab[18][20] ) );
  NOR2_X1 U502 ( .A1(n173), .A2(n137), .ZN(\ab[18][1] ) );
  NOR2_X1 U503 ( .A1(n65), .A2(n137), .ZN(\ab[18][19] ) );
  NOR2_X1 U504 ( .A1(n63), .A2(n137), .ZN(\ab[18][18] ) );
  NOR2_X1 U505 ( .A1(n46), .A2(n137), .ZN(\ab[18][17] ) );
  NOR2_X1 U506 ( .A1(n158), .A2(n137), .ZN(\ab[18][16] ) );
  NOR2_X1 U507 ( .A1(n159), .A2(n137), .ZN(\ab[18][15] ) );
  NOR2_X1 U508 ( .A1(n160), .A2(n137), .ZN(\ab[18][14] ) );
  NOR2_X1 U509 ( .A1(n161), .A2(n137), .ZN(\ab[18][13] ) );
  NOR2_X1 U510 ( .A1(n162), .A2(n137), .ZN(\ab[18][12] ) );
  NOR2_X1 U511 ( .A1(n163), .A2(n137), .ZN(\ab[18][11] ) );
  NOR2_X1 U512 ( .A1(n164), .A2(n137), .ZN(\ab[18][10] ) );
  NOR2_X1 U513 ( .A1(n174), .A2(n137), .ZN(\ab[18][0] ) );
  NOR2_X1 U514 ( .A1(n165), .A2(n138), .ZN(\ab[17][9] ) );
  NOR2_X1 U515 ( .A1(n166), .A2(n138), .ZN(\ab[17][8] ) );
  NOR2_X1 U516 ( .A1(n167), .A2(n138), .ZN(\ab[17][7] ) );
  NOR2_X1 U517 ( .A1(n168), .A2(n138), .ZN(\ab[17][6] ) );
  NOR2_X1 U518 ( .A1(n169), .A2(n138), .ZN(\ab[17][5] ) );
  NOR2_X1 U519 ( .A1(n170), .A2(n138), .ZN(\ab[17][4] ) );
  NOR2_X1 U520 ( .A1(n171), .A2(n138), .ZN(\ab[17][3] ) );
  NOR2_X1 U521 ( .A1(n172), .A2(n138), .ZN(\ab[17][2] ) );
  NOR2_X1 U522 ( .A1(n72), .A2(n138), .ZN(\ab[17][22] ) );
  NOR2_X1 U523 ( .A1(n73), .A2(n138), .ZN(\ab[17][21] ) );
  NOR2_X1 U524 ( .A1(n61), .A2(n138), .ZN(\ab[17][20] ) );
  NOR2_X1 U525 ( .A1(n173), .A2(n138), .ZN(\ab[17][1] ) );
  NOR2_X1 U526 ( .A1(n65), .A2(n138), .ZN(\ab[17][19] ) );
  NOR2_X1 U527 ( .A1(n63), .A2(n138), .ZN(\ab[17][18] ) );
  NOR2_X1 U528 ( .A1(n47), .A2(n138), .ZN(\ab[17][17] ) );
  NOR2_X1 U529 ( .A1(n158), .A2(n138), .ZN(\ab[17][16] ) );
  NOR2_X1 U530 ( .A1(n159), .A2(n138), .ZN(\ab[17][15] ) );
  NOR2_X1 U531 ( .A1(n160), .A2(n138), .ZN(\ab[17][14] ) );
  NOR2_X1 U532 ( .A1(n161), .A2(n138), .ZN(\ab[17][13] ) );
  NOR2_X1 U533 ( .A1(n162), .A2(n138), .ZN(\ab[17][12] ) );
  NOR2_X1 U534 ( .A1(n163), .A2(n138), .ZN(\ab[17][11] ) );
  NOR2_X1 U535 ( .A1(n164), .A2(n138), .ZN(\ab[17][10] ) );
  NOR2_X1 U536 ( .A1(n174), .A2(n138), .ZN(\ab[17][0] ) );
  NOR2_X1 U537 ( .A1(n165), .A2(n139), .ZN(\ab[16][9] ) );
  NOR2_X1 U538 ( .A1(n166), .A2(n139), .ZN(\ab[16][8] ) );
  NOR2_X1 U539 ( .A1(n167), .A2(n139), .ZN(\ab[16][7] ) );
  NOR2_X1 U540 ( .A1(n168), .A2(n139), .ZN(\ab[16][6] ) );
  NOR2_X1 U541 ( .A1(n169), .A2(n139), .ZN(\ab[16][5] ) );
  NOR2_X1 U542 ( .A1(n170), .A2(n139), .ZN(\ab[16][4] ) );
  NOR2_X1 U543 ( .A1(n171), .A2(n139), .ZN(\ab[16][3] ) );
  NOR2_X1 U544 ( .A1(n172), .A2(n139), .ZN(\ab[16][2] ) );
  NOR2_X1 U545 ( .A1(n72), .A2(n139), .ZN(\ab[16][22] ) );
  NOR2_X1 U546 ( .A1(n73), .A2(n139), .ZN(\ab[16][21] ) );
  NOR2_X1 U547 ( .A1(n61), .A2(n139), .ZN(\ab[16][20] ) );
  NOR2_X1 U548 ( .A1(n173), .A2(n139), .ZN(\ab[16][1] ) );
  NOR2_X1 U549 ( .A1(n65), .A2(n139), .ZN(\ab[16][19] ) );
  NOR2_X1 U550 ( .A1(n63), .A2(n139), .ZN(\ab[16][18] ) );
  NOR2_X1 U551 ( .A1(n46), .A2(n139), .ZN(\ab[16][17] ) );
  NOR2_X1 U552 ( .A1(n158), .A2(n139), .ZN(\ab[16][16] ) );
  NOR2_X1 U553 ( .A1(n159), .A2(n139), .ZN(\ab[16][15] ) );
  NOR2_X1 U554 ( .A1(n160), .A2(n139), .ZN(\ab[16][14] ) );
  NOR2_X1 U555 ( .A1(n161), .A2(n139), .ZN(\ab[16][13] ) );
  NOR2_X1 U556 ( .A1(n162), .A2(n139), .ZN(\ab[16][12] ) );
  NOR2_X1 U557 ( .A1(n163), .A2(n139), .ZN(\ab[16][11] ) );
  NOR2_X1 U558 ( .A1(n164), .A2(n139), .ZN(\ab[16][10] ) );
  NOR2_X1 U559 ( .A1(n174), .A2(n139), .ZN(\ab[16][0] ) );
  NOR2_X1 U560 ( .A1(n165), .A2(n140), .ZN(\ab[15][9] ) );
  NOR2_X1 U561 ( .A1(n166), .A2(n140), .ZN(\ab[15][8] ) );
  NOR2_X1 U562 ( .A1(n167), .A2(n140), .ZN(\ab[15][7] ) );
  NOR2_X1 U563 ( .A1(n168), .A2(n140), .ZN(\ab[15][6] ) );
  NOR2_X1 U564 ( .A1(n169), .A2(n140), .ZN(\ab[15][5] ) );
  NOR2_X1 U565 ( .A1(n170), .A2(n140), .ZN(\ab[15][4] ) );
  NOR2_X1 U566 ( .A1(n171), .A2(n140), .ZN(\ab[15][3] ) );
  NOR2_X1 U567 ( .A1(n172), .A2(n140), .ZN(\ab[15][2] ) );
  NOR2_X1 U568 ( .A1(n72), .A2(n140), .ZN(\ab[15][22] ) );
  NOR2_X1 U569 ( .A1(n73), .A2(n140), .ZN(\ab[15][21] ) );
  NOR2_X1 U570 ( .A1(n61), .A2(n140), .ZN(\ab[15][20] ) );
  NOR2_X1 U571 ( .A1(n173), .A2(n140), .ZN(\ab[15][1] ) );
  NOR2_X1 U572 ( .A1(n65), .A2(n140), .ZN(\ab[15][19] ) );
  NOR2_X1 U573 ( .A1(n63), .A2(n140), .ZN(\ab[15][18] ) );
  NOR2_X1 U574 ( .A1(n47), .A2(n140), .ZN(\ab[15][17] ) );
  NOR2_X1 U575 ( .A1(n158), .A2(n140), .ZN(\ab[15][16] ) );
  NOR2_X1 U576 ( .A1(n159), .A2(n140), .ZN(\ab[15][15] ) );
  NOR2_X1 U577 ( .A1(n160), .A2(n140), .ZN(\ab[15][14] ) );
  NOR2_X1 U578 ( .A1(n161), .A2(n140), .ZN(\ab[15][13] ) );
  NOR2_X1 U579 ( .A1(n162), .A2(n140), .ZN(\ab[15][12] ) );
  NOR2_X1 U580 ( .A1(n163), .A2(n140), .ZN(\ab[15][11] ) );
  NOR2_X1 U581 ( .A1(n164), .A2(n140), .ZN(\ab[15][10] ) );
  NOR2_X1 U582 ( .A1(n174), .A2(n140), .ZN(\ab[15][0] ) );
  NOR2_X1 U583 ( .A1(n165), .A2(n141), .ZN(\ab[14][9] ) );
  NOR2_X1 U584 ( .A1(n166), .A2(n141), .ZN(\ab[14][8] ) );
  NOR2_X1 U585 ( .A1(n167), .A2(n141), .ZN(\ab[14][7] ) );
  NOR2_X1 U586 ( .A1(n168), .A2(n141), .ZN(\ab[14][6] ) );
  NOR2_X1 U587 ( .A1(n169), .A2(n141), .ZN(\ab[14][5] ) );
  NOR2_X1 U588 ( .A1(n170), .A2(n141), .ZN(\ab[14][4] ) );
  NOR2_X1 U589 ( .A1(n171), .A2(n141), .ZN(\ab[14][3] ) );
  NOR2_X1 U590 ( .A1(n172), .A2(n141), .ZN(\ab[14][2] ) );
  NOR2_X1 U591 ( .A1(n72), .A2(n141), .ZN(\ab[14][22] ) );
  NOR2_X1 U592 ( .A1(n73), .A2(n141), .ZN(\ab[14][21] ) );
  NOR2_X1 U593 ( .A1(n61), .A2(n141), .ZN(\ab[14][20] ) );
  NOR2_X1 U594 ( .A1(n173), .A2(n141), .ZN(\ab[14][1] ) );
  NOR2_X1 U595 ( .A1(n65), .A2(n141), .ZN(\ab[14][19] ) );
  NOR2_X1 U596 ( .A1(n63), .A2(n141), .ZN(\ab[14][18] ) );
  NOR2_X1 U597 ( .A1(n46), .A2(n141), .ZN(\ab[14][17] ) );
  NOR2_X1 U598 ( .A1(n158), .A2(n141), .ZN(\ab[14][16] ) );
  NOR2_X1 U599 ( .A1(n159), .A2(n141), .ZN(\ab[14][15] ) );
  NOR2_X1 U600 ( .A1(n160), .A2(n141), .ZN(\ab[14][14] ) );
  NOR2_X1 U601 ( .A1(n161), .A2(n141), .ZN(\ab[14][13] ) );
  NOR2_X1 U602 ( .A1(n162), .A2(n141), .ZN(\ab[14][12] ) );
  NOR2_X1 U603 ( .A1(n163), .A2(n141), .ZN(\ab[14][11] ) );
  NOR2_X1 U604 ( .A1(n164), .A2(n141), .ZN(\ab[14][10] ) );
  NOR2_X1 U605 ( .A1(n174), .A2(n141), .ZN(\ab[14][0] ) );
  NOR2_X1 U606 ( .A1(n165), .A2(n142), .ZN(\ab[13][9] ) );
  NOR2_X1 U607 ( .A1(n166), .A2(n142), .ZN(\ab[13][8] ) );
  NOR2_X1 U608 ( .A1(n167), .A2(n142), .ZN(\ab[13][7] ) );
  NOR2_X1 U609 ( .A1(n168), .A2(n142), .ZN(\ab[13][6] ) );
  NOR2_X1 U610 ( .A1(n169), .A2(n142), .ZN(\ab[13][5] ) );
  NOR2_X1 U611 ( .A1(n170), .A2(n142), .ZN(\ab[13][4] ) );
  NOR2_X1 U612 ( .A1(n171), .A2(n142), .ZN(\ab[13][3] ) );
  NOR2_X1 U613 ( .A1(n172), .A2(n142), .ZN(\ab[13][2] ) );
  NOR2_X1 U614 ( .A1(n72), .A2(n142), .ZN(\ab[13][22] ) );
  NOR2_X1 U615 ( .A1(n73), .A2(n142), .ZN(\ab[13][21] ) );
  NOR2_X1 U616 ( .A1(n61), .A2(n142), .ZN(\ab[13][20] ) );
  NOR2_X1 U617 ( .A1(n173), .A2(n142), .ZN(\ab[13][1] ) );
  NOR2_X1 U618 ( .A1(n65), .A2(n142), .ZN(\ab[13][19] ) );
  NOR2_X1 U619 ( .A1(n63), .A2(n142), .ZN(\ab[13][18] ) );
  NOR2_X1 U620 ( .A1(n47), .A2(n142), .ZN(\ab[13][17] ) );
  NOR2_X1 U621 ( .A1(n158), .A2(n142), .ZN(\ab[13][16] ) );
  NOR2_X1 U622 ( .A1(n159), .A2(n142), .ZN(\ab[13][15] ) );
  NOR2_X1 U623 ( .A1(n160), .A2(n142), .ZN(\ab[13][14] ) );
  NOR2_X1 U624 ( .A1(n161), .A2(n142), .ZN(\ab[13][13] ) );
  NOR2_X1 U625 ( .A1(n162), .A2(n142), .ZN(\ab[13][12] ) );
  NOR2_X1 U626 ( .A1(n163), .A2(n142), .ZN(\ab[13][11] ) );
  NOR2_X1 U627 ( .A1(n164), .A2(n142), .ZN(\ab[13][10] ) );
  NOR2_X1 U628 ( .A1(n174), .A2(n142), .ZN(\ab[13][0] ) );
  NOR2_X1 U629 ( .A1(n165), .A2(n143), .ZN(\ab[12][9] ) );
  NOR2_X1 U630 ( .A1(n166), .A2(n143), .ZN(\ab[12][8] ) );
  NOR2_X1 U631 ( .A1(n167), .A2(n143), .ZN(\ab[12][7] ) );
  NOR2_X1 U632 ( .A1(n168), .A2(n143), .ZN(\ab[12][6] ) );
  NOR2_X1 U633 ( .A1(n169), .A2(n143), .ZN(\ab[12][5] ) );
  NOR2_X1 U634 ( .A1(n170), .A2(n143), .ZN(\ab[12][4] ) );
  NOR2_X1 U635 ( .A1(n171), .A2(n143), .ZN(\ab[12][3] ) );
  NOR2_X1 U636 ( .A1(n172), .A2(n143), .ZN(\ab[12][2] ) );
  NOR2_X1 U637 ( .A1(n72), .A2(n143), .ZN(\ab[12][22] ) );
  NOR2_X1 U638 ( .A1(n73), .A2(n143), .ZN(\ab[12][21] ) );
  NOR2_X1 U639 ( .A1(n61), .A2(n143), .ZN(\ab[12][20] ) );
  NOR2_X1 U640 ( .A1(n173), .A2(n143), .ZN(\ab[12][1] ) );
  NOR2_X1 U641 ( .A1(n65), .A2(n143), .ZN(\ab[12][19] ) );
  NOR2_X1 U642 ( .A1(n63), .A2(n143), .ZN(\ab[12][18] ) );
  NOR2_X1 U643 ( .A1(n46), .A2(n143), .ZN(\ab[12][17] ) );
  NOR2_X1 U644 ( .A1(n158), .A2(n143), .ZN(\ab[12][16] ) );
  NOR2_X1 U645 ( .A1(n159), .A2(n143), .ZN(\ab[12][15] ) );
  NOR2_X1 U646 ( .A1(n160), .A2(n143), .ZN(\ab[12][14] ) );
  NOR2_X1 U647 ( .A1(n161), .A2(n143), .ZN(\ab[12][13] ) );
  NOR2_X1 U648 ( .A1(n162), .A2(n143), .ZN(\ab[12][12] ) );
  NOR2_X1 U649 ( .A1(n163), .A2(n143), .ZN(\ab[12][11] ) );
  NOR2_X1 U650 ( .A1(n164), .A2(n143), .ZN(\ab[12][10] ) );
  NOR2_X1 U651 ( .A1(n174), .A2(n143), .ZN(\ab[12][0] ) );
  NOR2_X1 U652 ( .A1(n165), .A2(n144), .ZN(\ab[11][9] ) );
  NOR2_X1 U653 ( .A1(n166), .A2(n144), .ZN(\ab[11][8] ) );
  NOR2_X1 U654 ( .A1(n167), .A2(n144), .ZN(\ab[11][7] ) );
  NOR2_X1 U655 ( .A1(n168), .A2(n144), .ZN(\ab[11][6] ) );
  NOR2_X1 U656 ( .A1(n169), .A2(n144), .ZN(\ab[11][5] ) );
  NOR2_X1 U657 ( .A1(n170), .A2(n144), .ZN(\ab[11][4] ) );
  NOR2_X1 U658 ( .A1(n171), .A2(n144), .ZN(\ab[11][3] ) );
  NOR2_X1 U659 ( .A1(n172), .A2(n144), .ZN(\ab[11][2] ) );
  NOR2_X1 U660 ( .A1(n72), .A2(n144), .ZN(\ab[11][22] ) );
  NOR2_X1 U661 ( .A1(n73), .A2(n144), .ZN(\ab[11][21] ) );
  NOR2_X1 U662 ( .A1(n61), .A2(n144), .ZN(\ab[11][20] ) );
  NOR2_X1 U663 ( .A1(n173), .A2(n144), .ZN(\ab[11][1] ) );
  NOR2_X1 U664 ( .A1(n65), .A2(n144), .ZN(\ab[11][19] ) );
  NOR2_X1 U665 ( .A1(n63), .A2(n144), .ZN(\ab[11][18] ) );
  NOR2_X1 U666 ( .A1(n47), .A2(n144), .ZN(\ab[11][17] ) );
  NOR2_X1 U667 ( .A1(n158), .A2(n144), .ZN(\ab[11][16] ) );
  NOR2_X1 U668 ( .A1(n159), .A2(n144), .ZN(\ab[11][15] ) );
  NOR2_X1 U669 ( .A1(n160), .A2(n144), .ZN(\ab[11][14] ) );
  NOR2_X1 U670 ( .A1(n161), .A2(n144), .ZN(\ab[11][13] ) );
  NOR2_X1 U671 ( .A1(n162), .A2(n144), .ZN(\ab[11][12] ) );
  NOR2_X1 U672 ( .A1(n163), .A2(n144), .ZN(\ab[11][11] ) );
  NOR2_X1 U673 ( .A1(n164), .A2(n144), .ZN(\ab[11][10] ) );
  NOR2_X1 U674 ( .A1(n174), .A2(n144), .ZN(\ab[11][0] ) );
  NOR2_X1 U675 ( .A1(n165), .A2(n145), .ZN(\ab[10][9] ) );
  NOR2_X1 U676 ( .A1(n166), .A2(n145), .ZN(\ab[10][8] ) );
  NOR2_X1 U677 ( .A1(n167), .A2(n145), .ZN(\ab[10][7] ) );
  NOR2_X1 U678 ( .A1(n168), .A2(n145), .ZN(\ab[10][6] ) );
  NOR2_X1 U679 ( .A1(n169), .A2(n145), .ZN(\ab[10][5] ) );
  NOR2_X1 U680 ( .A1(n170), .A2(n145), .ZN(\ab[10][4] ) );
  NOR2_X1 U681 ( .A1(n171), .A2(n145), .ZN(\ab[10][3] ) );
  NOR2_X1 U682 ( .A1(n172), .A2(n145), .ZN(\ab[10][2] ) );
  NOR2_X1 U683 ( .A1(n72), .A2(n145), .ZN(\ab[10][22] ) );
  NOR2_X1 U684 ( .A1(n73), .A2(n145), .ZN(\ab[10][21] ) );
  NOR2_X1 U685 ( .A1(n61), .A2(n145), .ZN(\ab[10][20] ) );
  NOR2_X1 U686 ( .A1(n173), .A2(n145), .ZN(\ab[10][1] ) );
  NOR2_X1 U687 ( .A1(n65), .A2(n145), .ZN(\ab[10][19] ) );
  NOR2_X1 U688 ( .A1(n63), .A2(n145), .ZN(\ab[10][18] ) );
  NOR2_X1 U689 ( .A1(n46), .A2(n145), .ZN(\ab[10][17] ) );
  NOR2_X1 U690 ( .A1(n158), .A2(n145), .ZN(\ab[10][16] ) );
  NOR2_X1 U691 ( .A1(n159), .A2(n145), .ZN(\ab[10][15] ) );
  NOR2_X1 U692 ( .A1(n160), .A2(n145), .ZN(\ab[10][14] ) );
  NOR2_X1 U693 ( .A1(n161), .A2(n145), .ZN(\ab[10][13] ) );
  NOR2_X1 U694 ( .A1(n162), .A2(n145), .ZN(\ab[10][12] ) );
  NOR2_X1 U695 ( .A1(n163), .A2(n145), .ZN(\ab[10][11] ) );
  NOR2_X1 U696 ( .A1(n164), .A2(n145), .ZN(\ab[10][10] ) );
  NOR2_X1 U697 ( .A1(n174), .A2(n145), .ZN(\ab[10][0] ) );
  NOR2_X1 U698 ( .A1(n165), .A2(n78), .ZN(\ab[0][9] ) );
  NOR2_X1 U699 ( .A1(n166), .A2(n78), .ZN(\ab[0][8] ) );
  NOR2_X1 U700 ( .A1(n167), .A2(n67), .ZN(\ab[0][7] ) );
  NOR2_X1 U701 ( .A1(n168), .A2(n66), .ZN(\ab[0][6] ) );
  NOR2_X1 U702 ( .A1(n169), .A2(n66), .ZN(\ab[0][5] ) );
  NOR2_X1 U703 ( .A1(n170), .A2(n77), .ZN(\ab[0][4] ) );
  NOR2_X1 U704 ( .A1(n171), .A2(n77), .ZN(\ab[0][3] ) );
  NOR2_X1 U705 ( .A1(n172), .A2(n78), .ZN(\ab[0][2] ) );
  NOR2_X1 U706 ( .A1(n155), .A2(n67), .ZN(\ab[0][20] ) );
  NOR2_X1 U707 ( .A1(n173), .A2(n78), .ZN(\ab[0][1] ) );
  NOR2_X1 U708 ( .A1(n157), .A2(n77), .ZN(\ab[0][18] ) );
  NOR2_X1 U709 ( .A1(n47), .A2(n66), .ZN(\ab[0][17] ) );
  NOR2_X1 U710 ( .A1(n158), .A2(n77), .ZN(\ab[0][16] ) );
  NOR2_X1 U711 ( .A1(n159), .A2(n78), .ZN(\ab[0][15] ) );
  NOR2_X1 U712 ( .A1(n160), .A2(n78), .ZN(\ab[0][14] ) );
  NOR2_X1 U713 ( .A1(n161), .A2(n66), .ZN(\ab[0][13] ) );
  NOR2_X1 U714 ( .A1(n162), .A2(n66), .ZN(\ab[0][12] ) );
  NOR2_X1 U715 ( .A1(n163), .A2(n77), .ZN(\ab[0][11] ) );
  NOR2_X1 U716 ( .A1(n164), .A2(n77), .ZN(\ab[0][10] ) );
  NOR2_X1 U717 ( .A1(n174), .A2(n66), .ZN(PRODUCT[0]) );
endmodule


module FP_MULTIPLIER ( clk, rst, A, B, P_reg );
  input [31:0] A;
  input [31:0] B;
  output [31:0] P_reg;
  input clk, rst;
  wire   N105, N106, N107, N108, N109, N110, N111, N112, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n113, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, N96, N103, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234;
  wire   [31:0] P;
  wire   [47:0] mantissa_product;
  wire   [4:0] count;
  wire   [46:24] shifted_mantissa_product;
  wire   [7:0] exponent_sum;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  DFFR_X1 \P_reg_reg[31]  ( .D(P[31]), .CK(clk), .RN(n207), .Q(P_reg[31]) );
  DFFR_X1 \P_reg_reg[30]  ( .D(n219), .CK(clk), .RN(n207), .Q(P_reg[30]) );
  DFFR_X1 \P_reg_reg[29]  ( .D(n218), .CK(clk), .RN(n207), .Q(P_reg[29]) );
  DFFR_X1 \P_reg_reg[28]  ( .D(n217), .CK(clk), .RN(n207), .Q(P_reg[28]) );
  DFFR_X1 \P_reg_reg[27]  ( .D(n216), .CK(clk), .RN(n207), .Q(P_reg[27]) );
  DFFR_X1 \P_reg_reg[26]  ( .D(n215), .CK(clk), .RN(n207), .Q(P_reg[26]) );
  DFFR_X1 \P_reg_reg[25]  ( .D(n214), .CK(clk), .RN(n207), .Q(P_reg[25]) );
  DFFR_X1 \P_reg_reg[24]  ( .D(n213), .CK(clk), .RN(n207), .Q(P_reg[24]) );
  DFFR_X1 \P_reg_reg[23]  ( .D(n212), .CK(clk), .RN(n207), .Q(P_reg[23]) );
  DFFR_X1 \P_reg_reg[22]  ( .D(P[22]), .CK(clk), .RN(n207), .Q(P_reg[22]) );
  DFFR_X1 \P_reg_reg[21]  ( .D(P[21]), .CK(clk), .RN(n207), .Q(P_reg[21]) );
  DFFR_X1 \P_reg_reg[20]  ( .D(P[20]), .CK(clk), .RN(n207), .Q(P_reg[20]) );
  DFFR_X1 \P_reg_reg[19]  ( .D(P[19]), .CK(clk), .RN(n208), .Q(P_reg[19]) );
  DFFR_X1 \P_reg_reg[18]  ( .D(P[18]), .CK(clk), .RN(n208), .Q(P_reg[18]) );
  DFFR_X1 \P_reg_reg[17]  ( .D(P[17]), .CK(clk), .RN(n208), .Q(P_reg[17]) );
  DFFR_X1 \P_reg_reg[16]  ( .D(P[16]), .CK(clk), .RN(n208), .Q(P_reg[16]) );
  DFFR_X1 \P_reg_reg[15]  ( .D(P[15]), .CK(clk), .RN(n208), .Q(P_reg[15]) );
  DFFR_X1 \P_reg_reg[14]  ( .D(P[14]), .CK(clk), .RN(n208), .Q(P_reg[14]) );
  DFFR_X1 \P_reg_reg[13]  ( .D(P[13]), .CK(clk), .RN(n208), .Q(P_reg[13]) );
  DFFR_X1 \P_reg_reg[12]  ( .D(P[12]), .CK(clk), .RN(n208), .Q(P_reg[12]) );
  DFFR_X1 \P_reg_reg[11]  ( .D(P[11]), .CK(clk), .RN(n208), .Q(P_reg[11]) );
  DFFR_X1 \P_reg_reg[10]  ( .D(P[10]), .CK(clk), .RN(n208), .Q(P_reg[10]) );
  DFFR_X1 \P_reg_reg[9]  ( .D(P[9]), .CK(clk), .RN(n208), .Q(P_reg[9]) );
  DFFR_X1 \P_reg_reg[8]  ( .D(P[8]), .CK(clk), .RN(n208), .Q(P_reg[8]) );
  DFFR_X1 \P_reg_reg[7]  ( .D(P[7]), .CK(clk), .RN(n209), .Q(P_reg[7]) );
  DFFR_X1 \P_reg_reg[6]  ( .D(P[6]), .CK(clk), .RN(n209), .Q(P_reg[6]) );
  DFFR_X1 \P_reg_reg[5]  ( .D(P[5]), .CK(clk), .RN(n209), .Q(P_reg[5]) );
  DFFR_X1 \P_reg_reg[4]  ( .D(P[4]), .CK(clk), .RN(n209), .Q(P_reg[4]) );
  DFFR_X1 \P_reg_reg[3]  ( .D(P[3]), .CK(clk), .RN(n209), .Q(P_reg[3]) );
  DFFR_X1 \P_reg_reg[2]  ( .D(P[2]), .CK(clk), .RN(n209), .Q(P_reg[2]) );
  DFFR_X1 \P_reg_reg[1]  ( .D(P[1]), .CK(clk), .RN(n209), .Q(P_reg[1]) );
  DFFR_X1 \P_reg_reg[0]  ( .D(P[0]), .CK(clk), .RN(n209), .Q(P_reg[0]) );
  XOR2_X1 U122 ( .A(B[31]), .B(A[31]), .Z(P[31]) );
  FP_MULTIPLIER_DW01_inc_0 add_46 ( .A(exponent_sum), .SUM({N112, N111, N110, 
        N109, N108, N107, N106, N105}) );
  FP_MULTIPLIER_DW01_ash_0 sll_40 ( .A({n157, n168, mantissa_product[44:0]}), 
        .DATA_TC(1'b0), .SH({n211, count[3:0]}), .SH_TC(1'b0), .B({
        shifted_mantissa_product, SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23}) );
  FP_MULTIPLIER_DW01_add_0 add_0_root_sub_0_root_sub_44 ( .A(B[30:23]), .B({
        N103, n192, n191, n190, n189, n188, n134, N96}), .CI(1'b0), .SUM(
        exponent_sum) );
  FP_MULTIPLIER_DW02_mult_0 mult_36 ( .A({1'b1, A[22:0]}), .B({1'b1, B[22:0]}), 
        .TC(1'b0), .PRODUCT(mantissa_product) );
  NOR2_X1 U123 ( .A1(mantissa_product[40]), .A2(mantissa_product[39]), .ZN(
        n180) );
  CLKBUF_X1 U124 ( .A(n113), .Z(n124) );
  CLKBUF_X1 U125 ( .A(count[0]), .Z(n125) );
  OR3_X1 U126 ( .A1(mantissa_product[33]), .A2(mantissa_product[34]), .A3(n186), .ZN(n126) );
  AND3_X1 U127 ( .A1(n86), .A2(n87), .A3(n88), .ZN(n127) );
  AND2_X1 U128 ( .A1(n233), .A2(mantissa_product[24]), .ZN(n128) );
  NOR2_X1 U129 ( .A1(n187), .A2(n136), .ZN(n129) );
  AND2_X1 U130 ( .A1(n185), .A2(n181), .ZN(n130) );
  NAND2_X1 U131 ( .A1(n173), .A2(n176), .ZN(n131) );
  NAND2_X1 U132 ( .A1(n232), .A2(n201), .ZN(n132) );
  AND4_X1 U133 ( .A1(n115), .A2(n116), .A3(n117), .A4(n118), .ZN(n133) );
  XOR2_X1 U134 ( .A(A[24]), .B(A[23]), .Z(n134) );
  INV_X1 U135 ( .A(mantissa_product[34]), .ZN(n163) );
  CLKBUF_X1 U136 ( .A(n164), .Z(n135) );
  NAND2_X1 U137 ( .A1(n206), .A2(n150), .ZN(n136) );
  CLKBUF_X1 U138 ( .A(n87), .Z(n137) );
  OR2_X1 U139 ( .A1(n223), .A2(n138), .ZN(n102) );
  NAND2_X1 U140 ( .A1(mantissa_product[38]), .A2(n148), .ZN(n138) );
  NOR2_X1 U141 ( .A1(mantissa_product[40]), .A2(mantissa_product[39]), .ZN(
        n148) );
  AND2_X1 U142 ( .A1(n140), .A2(n139), .ZN(n105) );
  NOR2_X1 U143 ( .A1(n158), .A2(n178), .ZN(n139) );
  AND2_X1 U144 ( .A1(n97), .A2(n148), .ZN(n202) );
  NOR3_X1 U145 ( .A1(mantissa_product[47]), .A2(mantissa_product[46]), .A3(n93), .ZN(n140) );
  AND2_X1 U146 ( .A1(n182), .A2(n109), .ZN(n141) );
  AND2_X1 U147 ( .A1(mantissa_product[27]), .A2(n156), .ZN(n142) );
  NOR3_X1 U148 ( .A1(n141), .A2(n142), .A3(n92), .ZN(n107) );
  OR2_X1 U149 ( .A1(n187), .A2(n143), .ZN(n103) );
  NAND2_X1 U150 ( .A1(mantissa_product[32]), .A2(n150), .ZN(n143) );
  NAND2_X1 U151 ( .A1(n101), .A2(n183), .ZN(n144) );
  NOR2_X1 U152 ( .A1(n144), .A2(n145), .ZN(n172) );
  OR2_X1 U153 ( .A1(n132), .A2(n171), .ZN(n145) );
  AND2_X1 U154 ( .A1(n90), .A2(mantissa_product[37]), .ZN(n146) );
  AND2_X1 U155 ( .A1(mantissa_product[29]), .A2(n91), .ZN(n147) );
  NOR3_X1 U156 ( .A1(n92), .A2(n147), .A3(n146), .ZN(n89) );
  AND2_X1 U157 ( .A1(n164), .A2(n149), .ZN(n91) );
  NOR2_X1 U158 ( .A1(n174), .A2(n161), .ZN(n149) );
  NOR2_X1 U159 ( .A1(mantissa_product[34]), .A2(mantissa_product[33]), .ZN(
        n150) );
  AND2_X1 U160 ( .A1(n97), .A2(n180), .ZN(n151) );
  AND2_X1 U161 ( .A1(n151), .A2(n152), .ZN(n110) );
  AND2_X1 U162 ( .A1(n153), .A2(n183), .ZN(n152) );
  INV_X1 U163 ( .A(n171), .ZN(n153) );
  INV_X1 U164 ( .A(n223), .ZN(n154) );
  AND2_X1 U165 ( .A1(n108), .A2(n166), .ZN(n97) );
  OR2_X1 U166 ( .A1(n113), .A2(n155), .ZN(n187) );
  OR2_X1 U167 ( .A1(mantissa_product[41]), .A2(n131), .ZN(n155) );
  NOR2_X1 U168 ( .A1(n170), .A2(n171), .ZN(n156) );
  CLKBUF_X1 U169 ( .A(mantissa_product[46]), .Z(n157) );
  OR2_X1 U170 ( .A1(mantissa_product[41]), .A2(n159), .ZN(n158) );
  INV_X1 U171 ( .A(n173), .ZN(n159) );
  CLKBUF_X1 U172 ( .A(mantissa_product[47]), .Z(n160) );
  NAND2_X1 U173 ( .A1(n205), .A2(n181), .ZN(n161) );
  CLKBUF_X1 U174 ( .A(n104), .Z(n162) );
  OR2_X1 U175 ( .A1(n163), .A2(n186), .ZN(n104) );
  NOR2_X1 U176 ( .A1(n113), .A2(n165), .ZN(n164) );
  OR2_X1 U177 ( .A1(mantissa_product[41]), .A2(n159), .ZN(n165) );
  NOR2_X1 U178 ( .A1(n178), .A2(mantissa_product[41]), .ZN(n166) );
  CLKBUF_X1 U179 ( .A(n103), .Z(n167) );
  CLKBUF_X1 U180 ( .A(mantissa_product[45]), .Z(n168) );
  AND4_X1 U181 ( .A1(n102), .A2(n167), .A3(n162), .A4(n137), .ZN(n169) );
  NAND2_X1 U182 ( .A1(n101), .A2(n183), .ZN(n170) );
  NAND2_X1 U183 ( .A1(n130), .A2(n176), .ZN(n171) );
  AND3_X1 U184 ( .A1(n110), .A2(n232), .A3(n201), .ZN(n99) );
  AND2_X1 U185 ( .A1(n183), .A2(n180), .ZN(n173) );
  NAND2_X1 U186 ( .A1(n228), .A2(n229), .ZN(n174) );
  AND2_X1 U187 ( .A1(n97), .A2(n180), .ZN(n101) );
  NAND2_X1 U188 ( .A1(n228), .A2(n229), .ZN(n175) );
  INV_X1 U189 ( .A(n175), .ZN(n176) );
  CLKBUF_X1 U190 ( .A(n93), .Z(n177) );
  OR2_X1 U191 ( .A1(mantissa_product[45]), .A2(mantissa_product[44]), .ZN(n93)
         );
  NAND2_X1 U192 ( .A1(n172), .A2(n128), .ZN(n77) );
  NAND2_X1 U193 ( .A1(n89), .A2(n127), .ZN(count[1]) );
  NAND2_X1 U194 ( .A1(n225), .A2(n226), .ZN(n178) );
  NAND2_X1 U195 ( .A1(n140), .A2(n179), .ZN(n113) );
  INV_X1 U196 ( .A(n178), .ZN(n179) );
  NOR2_X1 U197 ( .A1(mantissa_product[34]), .A2(mantissa_product[33]), .ZN(
        n181) );
  NOR3_X1 U198 ( .A1(n177), .A2(n157), .A3(n160), .ZN(n182) );
  AND2_X1 U199 ( .A1(n204), .A2(n203), .ZN(n183) );
  AND2_X1 U200 ( .A1(n231), .A2(n199), .ZN(n184) );
  AND2_X1 U201 ( .A1(n205), .A2(n184), .ZN(n185) );
  NAND3_X1 U202 ( .A1(n105), .A2(n228), .A3(n229), .ZN(n186) );
  NOR4_X1 U203 ( .A1(count[2]), .A2(count[3]), .A3(n200), .A4(n76), .ZN(n75)
         );
  OR2_X1 U204 ( .A1(n125), .A2(n211), .ZN(n76) );
  INV_X1 U205 ( .A(mantissa_product[33]), .ZN(n230) );
  INV_X1 U206 ( .A(mantissa_product[37]), .ZN(n203) );
  INV_X1 U207 ( .A(mantissa_product[38]), .ZN(n204) );
  NAND4_X1 U208 ( .A1(n103), .A2(n87), .A3(n104), .A4(n102), .ZN(n83) );
  INV_X1 U209 ( .A(mantissa_product[35]), .ZN(n229) );
  AOI21_X1 U210 ( .B1(mantissa_product[42]), .B2(n225), .A(
        mantissa_product[44]), .ZN(n84) );
  INV_X1 U211 ( .A(mantissa_product[28]), .ZN(n199) );
  INV_X1 U212 ( .A(mantissa_product[42]), .ZN(n226) );
  INV_X1 U213 ( .A(mantissa_product[40]), .ZN(n227) );
  NAND3_X1 U214 ( .A1(n224), .A2(n220), .A3(n177), .ZN(n88) );
  INV_X1 U215 ( .A(mantissa_product[43]), .ZN(n225) );
  INV_X1 U216 ( .A(mantissa_product[36]), .ZN(n228) );
  INV_X1 U217 ( .A(n157), .ZN(n224) );
  BUF_X1 U218 ( .A(count[4]), .Z(n211) );
  INV_X1 U219 ( .A(mantissa_product[31]), .ZN(n206) );
  NAND3_X1 U220 ( .A1(n110), .A2(n232), .A3(mantissa_product[26]), .ZN(n78) );
  NAND4_X1 U221 ( .A1(n169), .A2(n94), .A3(n95), .A4(n96), .ZN(count[3]) );
  AND2_X1 U222 ( .A1(n86), .A2(n85), .ZN(n79) );
  OAI21_X1 U223 ( .B1(n168), .B2(n84), .A(n224), .ZN(n82) );
  NAND4_X1 U224 ( .A1(n78), .A2(n162), .A3(n106), .A4(n107), .ZN(count[2]) );
  NAND2_X1 U225 ( .A1(n225), .A2(n226), .ZN(n109) );
  INV_X1 U226 ( .A(mantissa_product[26]), .ZN(n201) );
  AND2_X1 U227 ( .A1(n75), .A2(n210), .ZN(n66) );
  NOR2_X1 U228 ( .A1(mantissa_product[25]), .A2(mantissa_product[24]), .ZN(n98) );
  INV_X1 U229 ( .A(mantissa_product[25]), .ZN(n233) );
  AND2_X1 U230 ( .A1(shifted_mantissa_product[32]), .A2(n210), .ZN(P[8]) );
  AND2_X1 U231 ( .A1(shifted_mantissa_product[33]), .A2(n210), .ZN(P[9]) );
  AND2_X1 U232 ( .A1(shifted_mantissa_product[31]), .A2(n210), .ZN(P[7]) );
  AND2_X1 U233 ( .A1(shifted_mantissa_product[39]), .A2(n210), .ZN(P[15]) );
  AND2_X1 U234 ( .A1(shifted_mantissa_product[34]), .A2(n210), .ZN(P[10]) );
  NOR2_X1 U235 ( .A1(n75), .A2(n133), .ZN(n67) );
  INV_X1 U236 ( .A(n74), .ZN(n212) );
  AOI22_X1 U237 ( .A1(N105), .A2(n66), .B1(exponent_sum[0]), .B2(n67), .ZN(n74) );
  INV_X1 U238 ( .A(n73), .ZN(n213) );
  AOI22_X1 U239 ( .A1(N106), .A2(n66), .B1(exponent_sum[1]), .B2(n67), .ZN(n73) );
  INV_X1 U240 ( .A(n72), .ZN(n214) );
  AOI22_X1 U241 ( .A1(N107), .A2(n66), .B1(exponent_sum[2]), .B2(n67), .ZN(n72) );
  INV_X1 U242 ( .A(n71), .ZN(n215) );
  AOI22_X1 U243 ( .A1(N108), .A2(n66), .B1(exponent_sum[3]), .B2(n67), .ZN(n71) );
  INV_X1 U244 ( .A(n70), .ZN(n216) );
  AOI22_X1 U245 ( .A1(N109), .A2(n66), .B1(exponent_sum[4]), .B2(n67), .ZN(n70) );
  INV_X1 U246 ( .A(n69), .ZN(n217) );
  AOI22_X1 U247 ( .A1(N110), .A2(n66), .B1(exponent_sum[5]), .B2(n67), .ZN(n69) );
  INV_X1 U248 ( .A(n68), .ZN(n218) );
  AOI22_X1 U249 ( .A1(N111), .A2(n66), .B1(exponent_sum[6]), .B2(n67), .ZN(n68) );
  INV_X1 U250 ( .A(n133), .ZN(n210) );
  BUF_X1 U251 ( .A(n234), .Z(n208) );
  BUF_X1 U252 ( .A(n234), .Z(n207) );
  BUF_X1 U253 ( .A(n234), .Z(n209) );
  INV_X1 U254 ( .A(n65), .ZN(n219) );
  AOI22_X1 U255 ( .A1(N112), .A2(n66), .B1(exponent_sum[7]), .B2(n67), .ZN(n65) );
  NOR4_X1 U256 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n122) );
  OR4_X1 U257 ( .A1(A[13]), .A2(A[12]), .A3(A[15]), .A4(A[14]), .ZN(n123) );
  NOR4_X1 U258 ( .A1(A[19]), .A2(A[18]), .A3(A[17]), .A4(A[16]), .ZN(n115) );
  XOR2_X1 U259 ( .A(A[30]), .B(n198), .Z(N103) );
  NAND2_X1 U260 ( .A1(A[29]), .A2(n197), .ZN(n198) );
  XOR2_X1 U261 ( .A(A[25]), .B(n195), .Z(n188) );
  XOR2_X1 U262 ( .A(A[26]), .B(n193), .Z(n189) );
  XOR2_X1 U263 ( .A(A[27]), .B(n194), .Z(n190) );
  XOR2_X1 U264 ( .A(A[28]), .B(n196), .Z(n191) );
  XOR2_X1 U265 ( .A(A[29]), .B(n197), .Z(n192) );
  AND2_X1 U266 ( .A1(A[25]), .A2(n195), .ZN(n193) );
  AND2_X1 U267 ( .A1(A[26]), .A2(n193), .ZN(n194) );
  AND2_X1 U268 ( .A1(A[24]), .A2(A[23]), .ZN(n195) );
  INV_X1 U269 ( .A(A[23]), .ZN(N96) );
  AND4_X1 U270 ( .A1(n119), .A2(n120), .A3(n121), .A4(n122), .ZN(n118) );
  NOR4_X1 U271 ( .A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n119) );
  NOR4_X1 U272 ( .A1(A[2]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n120) );
  NOR4_X1 U273 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[30]), .ZN(n121) );
  AND2_X1 U274 ( .A1(A[27]), .A2(n194), .ZN(n196) );
  AND2_X1 U275 ( .A1(A[28]), .A2(n196), .ZN(n197) );
  INV_X1 U276 ( .A(rst), .ZN(n234) );
  NOR4_X1 U277 ( .A1(n123), .A2(A[0]), .A3(A[11]), .A4(A[10]), .ZN(n117) );
  AND2_X1 U278 ( .A1(shifted_mantissa_product[38]), .A2(n210), .ZN(P[14]) );
  AND2_X1 U279 ( .A1(shifted_mantissa_product[37]), .A2(n210), .ZN(P[13]) );
  AND2_X1 U280 ( .A1(shifted_mantissa_product[36]), .A2(n210), .ZN(P[12]) );
  AND2_X1 U281 ( .A1(shifted_mantissa_product[35]), .A2(n210), .ZN(P[11]) );
  AOI21_X1 U282 ( .B1(n98), .B2(n172), .A(n100), .ZN(n95) );
  NAND2_X1 U283 ( .A1(n164), .A2(mantissa_product[36]), .ZN(n87) );
  NAND3_X1 U284 ( .A1(n135), .A2(n228), .A3(mantissa_product[35]), .ZN(n106)
         );
  NAND3_X1 U285 ( .A1(n154), .A2(n227), .A3(mantissa_product[39]), .ZN(n96) );
  NAND2_X1 U286 ( .A1(mantissa_product[40]), .A2(n154), .ZN(n85) );
  INV_X1 U287 ( .A(n124), .ZN(n221) );
  INV_X1 U288 ( .A(n160), .ZN(n220) );
  INV_X1 U289 ( .A(mantissa_product[29]), .ZN(n231) );
  NAND4_X1 U290 ( .A1(n89), .A2(n137), .A3(n88), .A4(n86), .ZN(n200) );
  INV_X1 U291 ( .A(mantissa_product[27]), .ZN(n232) );
  AND2_X1 U292 ( .A1(shifted_mantissa_product[30]), .A2(n210), .ZN(P[6]) );
  AND2_X1 U293 ( .A1(shifted_mantissa_product[29]), .A2(n210), .ZN(P[5]) );
  AND2_X1 U294 ( .A1(shifted_mantissa_product[28]), .A2(n210), .ZN(P[4]) );
  AND2_X1 U295 ( .A1(shifted_mantissa_product[27]), .A2(n210), .ZN(P[3]) );
  AND2_X1 U296 ( .A1(shifted_mantissa_product[26]), .A2(n210), .ZN(P[2]) );
  AND2_X1 U297 ( .A1(shifted_mantissa_product[25]), .A2(n210), .ZN(P[1]) );
  AND2_X1 U298 ( .A1(shifted_mantissa_product[24]), .A2(n210), .ZN(P[0]) );
  AND2_X1 U299 ( .A1(shifted_mantissa_product[43]), .A2(n210), .ZN(P[19]) );
  AND2_X1 U300 ( .A1(shifted_mantissa_product[46]), .A2(n210), .ZN(P[22]) );
  AND2_X1 U301 ( .A1(shifted_mantissa_product[45]), .A2(n210), .ZN(P[21]) );
  AND2_X1 U302 ( .A1(shifted_mantissa_product[44]), .A2(n210), .ZN(P[20]) );
  AND2_X1 U303 ( .A1(shifted_mantissa_product[42]), .A2(n210), .ZN(P[18]) );
  AND2_X1 U304 ( .A1(shifted_mantissa_product[41]), .A2(n210), .ZN(P[17]) );
  AND2_X1 U305 ( .A1(shifted_mantissa_product[40]), .A2(n210), .ZN(P[16]) );
  OAI21_X1 U306 ( .B1(mantissa_product[35]), .B2(mantissa_product[37]), .A(
        n202), .ZN(n94) );
  NOR2_X1 U307 ( .A1(mantissa_product[31]), .A2(mantissa_product[30]), .ZN(
        n205) );
  NOR4_X1 U308 ( .A1(A[22]), .A2(A[21]), .A3(A[20]), .A4(A[1]), .ZN(n116) );
  NAND3_X1 U309 ( .A1(n91), .A2(n231), .A3(mantissa_product[28]), .ZN(n86) );
  NOR2_X1 U310 ( .A1(n126), .A2(mantissa_product[32]), .ZN(count[4]) );
  NOR2_X1 U311 ( .A1(mantissa_product[38]), .A2(n222), .ZN(n90) );
  AOI221_X1 U312 ( .B1(mantissa_product[30]), .B2(n129), .C1(n82), .C2(n220), 
        .A(n83), .ZN(n80) );
  NAND4_X1 U313 ( .A1(n79), .A2(n80), .A3(n78), .A4(n77), .ZN(count[0]) );
  AOI221_X1 U314 ( .B1(mantissa_product[41]), .B2(n221), .C1(
        mantissa_product[25]), .C2(n99), .A(n100), .ZN(n111) );
  NOR3_X1 U315 ( .A1(mantissa_product[34]), .A2(n230), .A3(n187), .ZN(n100) );
  NAND4_X1 U316 ( .A1(n111), .A2(n85), .A3(n77), .A4(n167), .ZN(n92) );
  NOR3_X1 U317 ( .A1(mantissa_product[47]), .A2(mantissa_product[46]), .A3(n93), .ZN(n108) );
  INV_X1 U318 ( .A(n202), .ZN(n222) );
  INV_X1 U319 ( .A(n97), .ZN(n223) );
endmodule

