
module VerilogMultiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] ,
         \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173;
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2X2 U2 ( .IN1(n56), .IN2(n59), .Q(SUM[55]) );
  XOR2X2 U3 ( .IN1(n52), .IN2(n55), .Q(SUM[56]) );
  XOR2X2 U4 ( .IN1(n48), .IN2(n51), .Q(SUM[57]) );
  XOR3X2 U5 ( .IN1(B[60]), .IN2(A[60]), .IN3(n39), .Q(SUM[60]) );
  AND2X4 U6 ( .IN1(n105), .IN2(n104), .Q(n133) );
  NBUFFX2 U7 ( .INP(n152), .Z(n4) );
  NBUFFX2 U8 ( .INP(n137), .Z(n5) );
  XOR2X1 U9 ( .IN1(n3), .IN2(n71), .Q(SUM[52]) );
  NBUFFX4 U10 ( .INP(n68), .Z(n3) );
  XOR2X1 U11 ( .IN1(n60), .IN2(n63), .Q(SUM[54]) );
  OA21X1 U12 ( .IN1(n76), .IN2(n77), .IN3(n78), .Q(n1) );
  AO21X1 U13 ( .IN1(n68), .IN2(n16), .IN3(n69), .Q(n2) );
  AO21X1 U14 ( .IN1(n11), .IN2(n48), .IN3(n49), .Q(n6) );
  INVX0 U15 ( .INP(n42), .ZN(n9) );
  INVX0 U16 ( .INP(n46), .ZN(n10) );
  INVX0 U17 ( .INP(n62), .ZN(n14) );
  INVX0 U18 ( .INP(n58), .ZN(n13) );
  INVX0 U19 ( .INP(n54), .ZN(n12) );
  INVX0 U20 ( .INP(n50), .ZN(n11) );
  INVX0 U21 ( .INP(n66), .ZN(n15) );
  INVX0 U22 ( .INP(n70), .ZN(n16) );
  INVX0 U23 ( .INP(n168), .ZN(n36) );
  XOR2X1 U24 ( .IN1(n43), .IN2(n40), .Q(SUM[59]) );
  XOR2X1 U25 ( .IN1(n6), .IN2(n47), .Q(SUM[58]) );
  INVX0 U26 ( .INP(n73), .ZN(n17) );
  INVX0 U27 ( .INP(n77), .ZN(n18) );
  INVX0 U28 ( .INP(n81), .ZN(n19) );
  INVX0 U29 ( .INP(n116), .ZN(n25) );
  INVX0 U30 ( .INP(n88), .ZN(n21) );
  INVX0 U31 ( .INP(n85), .ZN(n20) );
  INVX0 U32 ( .INP(n123), .ZN(n28) );
  INVX0 U33 ( .INP(n141), .ZN(n32) );
  INVX0 U34 ( .INP(n93), .ZN(n22) );
  INVX0 U35 ( .INP(n121), .ZN(n26) );
  INVX0 U36 ( .INP(n96), .ZN(n23) );
  INVX0 U37 ( .INP(n139), .ZN(n30) );
  INVX0 U38 ( .INP(n124), .ZN(n27) );
  INVX0 U39 ( .INP(n99), .ZN(n24) );
  INVX0 U40 ( .INP(n142), .ZN(n31) );
  XOR2X1 U41 ( .IN1(n167), .IN2(n169), .Q(SUM[32]) );
  XOR3X1 U42 ( .IN1(B[61]), .IN2(A[61]), .IN3(n7), .Q(SUM[61]) );
  AO22X1 U43 ( .IN1(n38), .IN2(B[60]), .IN3(n39), .IN4(A[60]), .Q(n7) );
  INVX0 U44 ( .INP(n172), .ZN(n37) );
  INVX0 U45 ( .INP(n4), .ZN(n34) );
  INVX0 U46 ( .INP(n158), .ZN(n35) );
  OAI21X1 U47 ( .IN1(n170), .IN2(n171), .IN3(n172), .QN(n8) );
  OR4X1 U48 ( .IN1(n116), .IN2(n119), .IN3(n122), .IN4(n125), .Q(n101) );
  INVX0 U49 ( .INP(n134), .ZN(n29) );
  INVX0 U50 ( .INP(n153), .ZN(n33) );
  OR2X1 U51 ( .IN1(A[60]), .IN2(n39), .Q(n38) );
  AO21X1 U52 ( .IN1(n40), .IN2(n9), .IN3(n41), .Q(n39) );
  NOR2X0 U53 ( .IN1(n42), .IN2(n41), .QN(n43) );
  NOR2X0 U54 ( .IN1(B[59]), .IN2(A[59]), .QN(n42) );
  AND2X1 U55 ( .IN1(B[59]), .IN2(A[59]), .Q(n41) );
  AO21X1 U56 ( .IN1(n44), .IN2(n10), .IN3(n45), .Q(n40) );
  NOR2X0 U57 ( .IN1(n45), .IN2(n46), .QN(n47) );
  NOR2X0 U58 ( .IN1(B[58]), .IN2(A[58]), .QN(n46) );
  AND2X1 U59 ( .IN1(B[58]), .IN2(A[58]), .Q(n45) );
  AO21X1 U60 ( .IN1(n11), .IN2(n48), .IN3(n49), .Q(n44) );
  NOR2X0 U61 ( .IN1(n49), .IN2(n50), .QN(n51) );
  NOR2X0 U62 ( .IN1(A[57]), .IN2(B[57]), .QN(n50) );
  AND2X1 U63 ( .IN1(A[57]), .IN2(B[57]), .Q(n49) );
  AO21X1 U64 ( .IN1(n52), .IN2(n12), .IN3(n53), .Q(n48) );
  NOR2X0 U65 ( .IN1(n53), .IN2(n54), .QN(n55) );
  NOR2X0 U66 ( .IN1(B[56]), .IN2(A[56]), .QN(n54) );
  AND2X1 U67 ( .IN1(B[56]), .IN2(A[56]), .Q(n53) );
  AO21X1 U68 ( .IN1(n56), .IN2(n13), .IN3(n57), .Q(n52) );
  NOR2X0 U69 ( .IN1(n57), .IN2(n58), .QN(n59) );
  NOR2X0 U70 ( .IN1(A[55]), .IN2(B[55]), .QN(n58) );
  AND2X1 U71 ( .IN1(A[55]), .IN2(B[55]), .Q(n57) );
  AO21X1 U72 ( .IN1(n60), .IN2(n14), .IN3(n61), .Q(n56) );
  NOR2X0 U73 ( .IN1(n61), .IN2(n62), .QN(n63) );
  NOR2X0 U74 ( .IN1(B[54]), .IN2(A[54]), .QN(n62) );
  AND2X1 U75 ( .IN1(B[54]), .IN2(A[54]), .Q(n61) );
  AO21X1 U76 ( .IN1(n64), .IN2(n15), .IN3(n65), .Q(n60) );
  XOR2X1 U77 ( .IN1(n67), .IN2(n2), .Q(SUM[53]) );
  NOR2X0 U78 ( .IN1(n65), .IN2(n66), .QN(n67) );
  NOR2X0 U79 ( .IN1(B[53]), .IN2(A[53]), .QN(n66) );
  AND2X1 U80 ( .IN1(B[53]), .IN2(A[53]), .Q(n65) );
  AO21X1 U81 ( .IN1(n68), .IN2(n16), .IN3(n69), .Q(n64) );
  NOR2X0 U82 ( .IN1(n69), .IN2(n70), .QN(n71) );
  NOR2X0 U83 ( .IN1(B[52]), .IN2(A[52]), .QN(n70) );
  AND2X1 U84 ( .IN1(B[52]), .IN2(A[52]), .Q(n69) );
  OAI21X1 U85 ( .IN1(n73), .IN2(n72), .IN3(n74), .QN(n68) );
  XOR2X1 U86 ( .IN1(n75), .IN2(n1), .Q(SUM[51]) );
  OA21X1 U87 ( .IN1(n76), .IN2(n77), .IN3(n78), .Q(n72) );
  NAND2X0 U88 ( .IN1(n17), .IN2(n74), .QN(n75) );
  NAND2X0 U89 ( .IN1(B[51]), .IN2(A[51]), .QN(n74) );
  NOR2X0 U90 ( .IN1(B[51]), .IN2(A[51]), .QN(n73) );
  XOR2X1 U91 ( .IN1(n79), .IN2(n76), .Q(SUM[50]) );
  OA21X1 U92 ( .IN1(n81), .IN2(n80), .IN3(n82), .Q(n76) );
  NAND2X0 U93 ( .IN1(n18), .IN2(n78), .QN(n79) );
  NAND2X0 U94 ( .IN1(B[50]), .IN2(A[50]), .QN(n78) );
  NOR2X0 U95 ( .IN1(B[50]), .IN2(A[50]), .QN(n77) );
  XOR2X1 U96 ( .IN1(n83), .IN2(n80), .Q(SUM[49]) );
  OA21X1 U97 ( .IN1(n85), .IN2(n84), .IN3(n86), .Q(n80) );
  NAND2X0 U98 ( .IN1(n19), .IN2(n82), .QN(n83) );
  NAND2X0 U99 ( .IN1(B[49]), .IN2(A[49]), .QN(n82) );
  NOR2X0 U100 ( .IN1(B[49]), .IN2(A[49]), .QN(n81) );
  XOR2X1 U101 ( .IN1(n87), .IN2(n84), .Q(SUM[48]) );
  OA21X1 U102 ( .IN1(n88), .IN2(n89), .IN3(n90), .Q(n84) );
  OA21X1 U103 ( .IN1(n91), .IN2(n92), .IN3(n93), .Q(n89) );
  OA21X1 U104 ( .IN1(n94), .IN2(n95), .IN3(n96), .Q(n92) );
  OA21X1 U105 ( .IN1(n97), .IN2(n98), .IN3(n99), .Q(n95) );
  OA21X1 U106 ( .IN1(n101), .IN2(n100), .IN3(n102), .Q(n98) );
  OA221X1 U107 ( .IN1(n103), .IN2(n104), .IN3(n103), .IN4(n105), .IN5(n106), 
        .Q(n100) );
  NAND2X0 U108 ( .IN1(n20), .IN2(n86), .QN(n87) );
  NAND2X0 U109 ( .IN1(B[48]), .IN2(A[48]), .QN(n86) );
  NOR2X0 U110 ( .IN1(B[48]), .IN2(A[48]), .QN(n85) );
  XOR2X1 U111 ( .IN1(n107), .IN2(n108), .Q(SUM[47]) );
  OA21X1 U112 ( .IN1(n91), .IN2(n109), .IN3(n93), .Q(n108) );
  NAND2X0 U113 ( .IN1(n21), .IN2(n90), .QN(n107) );
  NAND2X0 U114 ( .IN1(B[47]), .IN2(A[47]), .QN(n90) );
  NOR2X0 U115 ( .IN1(B[47]), .IN2(A[47]), .QN(n88) );
  XNOR2X1 U116 ( .IN1(n109), .IN2(n110), .Q(SUM[46]) );
  NOR2X0 U117 ( .IN1(n22), .IN2(n91), .QN(n110) );
  NOR2X0 U118 ( .IN1(B[46]), .IN2(A[46]), .QN(n91) );
  NAND2X0 U119 ( .IN1(B[46]), .IN2(A[46]), .QN(n93) );
  OA21X1 U120 ( .IN1(n111), .IN2(n94), .IN3(n96), .Q(n109) );
  XNOR2X1 U121 ( .IN1(n111), .IN2(n112), .Q(SUM[45]) );
  NOR2X0 U122 ( .IN1(n23), .IN2(n94), .QN(n112) );
  NOR2X0 U123 ( .IN1(A[45]), .IN2(B[45]), .QN(n94) );
  NAND2X0 U124 ( .IN1(B[45]), .IN2(A[45]), .QN(n96) );
  OA21X1 U125 ( .IN1(n113), .IN2(n97), .IN3(n99), .Q(n111) );
  XNOR2X1 U126 ( .IN1(n113), .IN2(n114), .Q(SUM[44]) );
  NOR2X0 U127 ( .IN1(n24), .IN2(n97), .QN(n114) );
  NOR2X0 U128 ( .IN1(B[44]), .IN2(A[44]), .QN(n97) );
  NAND2X0 U129 ( .IN1(B[44]), .IN2(A[44]), .QN(n99) );
  OA21X1 U130 ( .IN1(n101), .IN2(n115), .IN3(n102), .Q(n113) );
  OA21X1 U131 ( .IN1(n116), .IN2(n117), .IN3(n118), .Q(n102) );
  OA21X1 U132 ( .IN1(n119), .IN2(n120), .IN3(n121), .Q(n117) );
  OA21X1 U133 ( .IN1(n122), .IN2(n123), .IN3(n124), .Q(n120) );
  XOR2X1 U134 ( .IN1(n126), .IN2(n127), .Q(SUM[43]) );
  OA21X1 U135 ( .IN1(n119), .IN2(n128), .IN3(n121), .Q(n127) );
  NAND2X0 U136 ( .IN1(n25), .IN2(n118), .QN(n126) );
  NAND2X0 U137 ( .IN1(B[43]), .IN2(A[43]), .QN(n118) );
  NOR2X0 U138 ( .IN1(B[43]), .IN2(A[43]), .QN(n116) );
  XNOR2X1 U139 ( .IN1(n128), .IN2(n129), .Q(SUM[42]) );
  NOR2X0 U140 ( .IN1(n26), .IN2(n119), .QN(n129) );
  NOR2X0 U141 ( .IN1(A[42]), .IN2(B[42]), .QN(n119) );
  NAND2X0 U142 ( .IN1(B[42]), .IN2(A[42]), .QN(n121) );
  OA21X1 U143 ( .IN1(n130), .IN2(n122), .IN3(n124), .Q(n128) );
  XNOR2X1 U144 ( .IN1(n130), .IN2(n131), .Q(SUM[41]) );
  NOR2X0 U145 ( .IN1(n27), .IN2(n122), .QN(n131) );
  NOR2X0 U146 ( .IN1(B[41]), .IN2(A[41]), .QN(n122) );
  NAND2X0 U147 ( .IN1(B[41]), .IN2(A[41]), .QN(n124) );
  OA21X1 U148 ( .IN1(n115), .IN2(n125), .IN3(n123), .Q(n130) );
  XNOR2X1 U149 ( .IN1(n115), .IN2(n132), .Q(SUM[40]) );
  NOR2X0 U150 ( .IN1(n28), .IN2(n125), .QN(n132) );
  NOR2X0 U151 ( .IN1(B[40]), .IN2(A[40]), .QN(n125) );
  NAND2X0 U152 ( .IN1(B[40]), .IN2(A[40]), .QN(n123) );
  OA21X1 U153 ( .IN1(n103), .IN2(n133), .IN3(n106), .Q(n115) );
  OA21X1 U154 ( .IN1(n134), .IN2(n135), .IN3(n136), .Q(n106) );
  OA21X1 U155 ( .IN1(n137), .IN2(n138), .IN3(n139), .Q(n135) );
  OA21X1 U156 ( .IN1(n140), .IN2(n141), .IN3(n142), .Q(n138) );
  OR4X1 U157 ( .IN1(n134), .IN2(n137), .IN3(n140), .IN4(n143), .Q(n103) );
  XOR2X1 U158 ( .IN1(n144), .IN2(n145), .Q(SUM[39]) );
  OA21X1 U159 ( .IN1(n5), .IN2(n146), .IN3(n139), .Q(n145) );
  NAND2X0 U160 ( .IN1(n29), .IN2(n136), .QN(n144) );
  NAND2X0 U161 ( .IN1(B[39]), .IN2(A[39]), .QN(n136) );
  NOR2X0 U162 ( .IN1(B[39]), .IN2(A[39]), .QN(n134) );
  XNOR2X1 U163 ( .IN1(n146), .IN2(n147), .Q(SUM[38]) );
  NOR2X0 U164 ( .IN1(n5), .IN2(n30), .QN(n147) );
  NOR2X0 U165 ( .IN1(B[38]), .IN2(A[38]), .QN(n137) );
  NAND2X0 U166 ( .IN1(B[38]), .IN2(A[38]), .QN(n139) );
  OA21X1 U167 ( .IN1(n148), .IN2(n140), .IN3(n142), .Q(n146) );
  XNOR2X1 U168 ( .IN1(n148), .IN2(n149), .Q(SUM[37]) );
  NOR2X0 U169 ( .IN1(n140), .IN2(n31), .QN(n149) );
  NOR2X0 U170 ( .IN1(B[37]), .IN2(A[37]), .QN(n140) );
  NAND2X0 U171 ( .IN1(B[37]), .IN2(A[37]), .QN(n142) );
  OA21X1 U172 ( .IN1(n133), .IN2(n143), .IN3(n141), .Q(n148) );
  XNOR2X1 U173 ( .IN1(n133), .IN2(n150), .Q(SUM[36]) );
  NOR2X0 U174 ( .IN1(n32), .IN2(n143), .QN(n150) );
  NOR2X0 U175 ( .IN1(B[36]), .IN2(A[36]), .QN(n143) );
  NAND2X0 U176 ( .IN1(B[36]), .IN2(A[36]), .QN(n141) );
  NAND4X0 U177 ( .IN1(n8), .IN2(n36), .IN3(n35), .IN4(n151), .QN(n104) );
  NOR2X0 U178 ( .IN1(n152), .IN2(n153), .QN(n151) );
  OA21X1 U179 ( .IN1(n153), .IN2(n154), .IN3(n155), .Q(n105) );
  OA21X1 U180 ( .IN1(n152), .IN2(n156), .IN3(n157), .Q(n154) );
  OA21X1 U181 ( .IN1(n158), .IN2(n159), .IN3(n160), .Q(n156) );
  XOR2X1 U182 ( .IN1(n161), .IN2(n162), .Q(SUM[35]) );
  OA21X1 U183 ( .IN1(n4), .IN2(n163), .IN3(n157), .Q(n162) );
  NAND2X0 U184 ( .IN1(n33), .IN2(n155), .QN(n161) );
  NAND2X0 U185 ( .IN1(B[35]), .IN2(A[35]), .QN(n155) );
  NOR2X0 U186 ( .IN1(B[35]), .IN2(A[35]), .QN(n153) );
  XOR2X1 U187 ( .IN1(n164), .IN2(n163), .Q(SUM[34]) );
  OA21X1 U188 ( .IN1(n158), .IN2(n165), .IN3(n160), .Q(n163) );
  NAND2X0 U189 ( .IN1(n34), .IN2(n157), .QN(n164) );
  NAND2X0 U190 ( .IN1(B[34]), .IN2(A[34]), .QN(n157) );
  NOR2X0 U191 ( .IN1(B[34]), .IN2(A[34]), .QN(n152) );
  XOR2X1 U192 ( .IN1(n166), .IN2(n165), .Q(SUM[33]) );
  OA21X1 U193 ( .IN1(n167), .IN2(n168), .IN3(n159), .Q(n165) );
  NAND2X0 U194 ( .IN1(n35), .IN2(n160), .QN(n166) );
  NAND2X0 U195 ( .IN1(A[33]), .IN2(B[33]), .QN(n160) );
  NOR2X0 U196 ( .IN1(B[33]), .IN2(A[33]), .QN(n158) );
  OA21X1 U197 ( .IN1(n170), .IN2(n171), .IN3(n172), .Q(n167) );
  NAND2X0 U198 ( .IN1(n36), .IN2(n159), .QN(n169) );
  NAND2X0 U199 ( .IN1(B[32]), .IN2(A[32]), .QN(n159) );
  NOR2X0 U200 ( .IN1(B[32]), .IN2(A[32]), .QN(n168) );
  XNOR2X1 U201 ( .IN1(n170), .IN2(n173), .Q(SUM[31]) );
  NOR2X0 U202 ( .IN1(n171), .IN2(n37), .QN(n173) );
  NOR2X0 U203 ( .IN1(A[31]), .IN2(B[31]), .QN(n171) );
  NAND2X0 U204 ( .IN1(B[31]), .IN2(A[31]), .QN(n172) );
  OA21X1 U205 ( .IN1(A[30]), .IN2(B[30]), .IN3(n170), .Q(SUM[30]) );
  NAND2X0 U206 ( .IN1(B[30]), .IN2(A[30]), .QN(n170) );
endmodule


module VerilogMultiplier_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \ab[31][31] , \ab[31][30] , \ab[31][29] , \ab[31][28] , \ab[31][27] ,
         \ab[31][26] , \ab[31][25] , \ab[31][24] , \ab[31][23] , \ab[31][22] ,
         \ab[31][21] , \ab[31][20] , \ab[31][19] , \ab[31][18] , \ab[31][17] ,
         \ab[31][16] , \ab[31][15] , \ab[31][14] , \ab[31][13] , \ab[31][12] ,
         \ab[31][11] , \ab[31][10] , \ab[31][9] , \ab[31][8] , \ab[31][7] ,
         \ab[31][6] , \ab[31][5] , \ab[31][4] , \ab[31][3] , \ab[31][2] ,
         \ab[31][1] , \ab[31][0] , \ab[30][31] , \ab[30][30] , \ab[30][29] ,
         \ab[30][28] , \ab[30][27] , \ab[30][26] , \ab[30][25] , \ab[30][24] ,
         \ab[30][23] , \ab[30][22] , \ab[30][21] , \ab[30][20] , \ab[30][19] ,
         \ab[30][18] , \ab[30][17] , \ab[30][16] , \ab[30][15] , \ab[30][14] ,
         \ab[30][13] , \ab[30][12] , \ab[30][11] , \ab[30][10] , \ab[30][9] ,
         \ab[30][8] , \ab[30][7] , \ab[30][6] , \ab[30][5] , \ab[30][4] ,
         \ab[30][3] , \ab[30][2] , \ab[30][1] , \ab[30][0] , \ab[29][31] ,
         \ab[29][30] , \ab[29][29] , \ab[29][28] , \ab[29][27] , \ab[29][26] ,
         \ab[29][25] , \ab[29][24] , \ab[29][23] , \ab[29][22] , \ab[29][21] ,
         \ab[29][20] , \ab[29][19] , \ab[29][18] , \ab[29][17] , \ab[29][16] ,
         \ab[29][15] , \ab[29][14] , \ab[29][13] , \ab[29][12] , \ab[29][11] ,
         \ab[29][10] , \ab[29][9] , \ab[29][8] , \ab[29][7] , \ab[29][6] ,
         \ab[29][5] , \ab[29][4] , \ab[29][3] , \ab[29][2] , \ab[29][1] ,
         \ab[29][0] , \ab[28][31] , \ab[28][30] , \ab[28][29] , \ab[28][28] ,
         \ab[28][27] , \ab[28][26] , \ab[28][25] , \ab[28][24] , \ab[28][23] ,
         \ab[28][22] , \ab[28][21] , \ab[28][20] , \ab[28][19] , \ab[28][18] ,
         \ab[28][17] , \ab[28][16] , \ab[28][15] , \ab[28][14] , \ab[28][13] ,
         \ab[28][12] , \ab[28][11] , \ab[28][10] , \ab[28][9] , \ab[28][8] ,
         \ab[28][7] , \ab[28][6] , \ab[28][5] , \ab[28][4] , \ab[28][3] ,
         \ab[28][2] , \ab[28][1] , \ab[28][0] , \ab[27][31] , \ab[27][30] ,
         \ab[27][29] , \ab[27][28] , \ab[27][27] , \ab[27][26] , \ab[27][25] ,
         \ab[27][24] , \ab[27][23] , \ab[27][22] , \ab[27][21] , \ab[27][20] ,
         \ab[27][19] , \ab[27][18] , \ab[27][17] , \ab[27][16] , \ab[27][15] ,
         \ab[27][14] , \ab[27][13] , \ab[27][12] , \ab[27][11] , \ab[27][10] ,
         \ab[27][9] , \ab[27][8] , \ab[27][7] , \ab[27][6] , \ab[27][5] ,
         \ab[27][4] , \ab[27][3] , \ab[27][2] , \ab[27][1] , \ab[27][0] ,
         \ab[26][31] , \ab[26][30] , \ab[26][29] , \ab[26][28] , \ab[26][27] ,
         \ab[26][26] , \ab[26][25] , \ab[26][24] , \ab[26][23] , \ab[26][22] ,
         \ab[26][21] , \ab[26][20] , \ab[26][19] , \ab[26][18] , \ab[26][17] ,
         \ab[26][16] , \ab[26][15] , \ab[26][14] , \ab[26][13] , \ab[26][12] ,
         \ab[26][11] , \ab[26][10] , \ab[26][9] , \ab[26][8] , \ab[26][7] ,
         \ab[26][6] , \ab[26][5] , \ab[26][4] , \ab[26][3] , \ab[26][2] ,
         \ab[26][1] , \ab[26][0] , \ab[25][31] , \ab[25][30] , \ab[25][29] ,
         \ab[25][28] , \ab[25][27] , \ab[25][26] , \ab[25][25] , \ab[25][24] ,
         \ab[25][23] , \ab[25][22] , \ab[25][21] , \ab[25][20] , \ab[25][19] ,
         \ab[25][18] , \ab[25][17] , \ab[25][16] , \ab[25][15] , \ab[25][14] ,
         \ab[25][13] , \ab[25][12] , \ab[25][11] , \ab[25][10] , \ab[25][9] ,
         \ab[25][8] , \ab[25][7] , \ab[25][6] , \ab[25][5] , \ab[25][4] ,
         \ab[25][3] , \ab[25][2] , \ab[25][1] , \ab[25][0] , \ab[24][31] ,
         \ab[24][30] , \ab[24][29] , \ab[24][28] , \ab[24][27] , \ab[24][26] ,
         \ab[24][25] , \ab[24][24] , \ab[24][23] , \ab[24][22] , \ab[24][21] ,
         \ab[24][20] , \ab[24][19] , \ab[24][18] , \ab[24][17] , \ab[24][16] ,
         \ab[24][15] , \ab[24][14] , \ab[24][13] , \ab[24][12] , \ab[24][11] ,
         \ab[24][10] , \ab[24][9] , \ab[24][8] , \ab[24][7] , \ab[24][6] ,
         \ab[24][5] , \ab[24][4] , \ab[24][3] , \ab[24][2] , \ab[24][1] ,
         \ab[24][0] , \ab[23][31] , \ab[23][30] , \ab[23][29] , \ab[23][28] ,
         \ab[23][27] , \ab[23][26] , \ab[23][25] , \ab[23][24] , \ab[23][23] ,
         \ab[23][22] , \ab[23][21] , \ab[23][20] , \ab[23][19] , \ab[23][18] ,
         \ab[23][17] , \ab[23][16] , \ab[23][15] , \ab[23][14] , \ab[23][13] ,
         \ab[23][12] , \ab[23][11] , \ab[23][10] , \ab[23][9] , \ab[23][8] ,
         \ab[23][7] , \ab[23][6] , \ab[23][5] , \ab[23][4] , \ab[23][3] ,
         \ab[23][2] , \ab[23][1] , \ab[23][0] , \ab[22][31] , \ab[22][30] ,
         \ab[22][29] , \ab[22][28] , \ab[22][27] , \ab[22][26] , \ab[22][25] ,
         \ab[22][24] , \ab[22][23] , \ab[22][22] , \ab[22][21] , \ab[22][20] ,
         \ab[22][19] , \ab[22][18] , \ab[22][17] , \ab[22][16] , \ab[22][15] ,
         \ab[22][14] , \ab[22][13] , \ab[22][12] , \ab[22][11] , \ab[22][10] ,
         \ab[22][9] , \ab[22][8] , \ab[22][7] , \ab[22][6] , \ab[22][5] ,
         \ab[22][4] , \ab[22][3] , \ab[22][2] , \ab[22][1] , \ab[22][0] ,
         \ab[21][31] , \ab[21][30] , \ab[21][29] , \ab[21][28] , \ab[21][27] ,
         \ab[21][26] , \ab[21][25] , \ab[21][24] , \ab[21][23] , \ab[21][22] ,
         \ab[21][21] , \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] ,
         \ab[21][16] , \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] ,
         \ab[21][11] , \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] ,
         \ab[21][6] , \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] ,
         \ab[21][1] , \ab[21][0] , \ab[20][31] , \ab[20][30] , \ab[20][29] ,
         \ab[20][28] , \ab[20][27] , \ab[20][26] , \ab[20][25] , \ab[20][24] ,
         \ab[20][23] , \ab[20][22] , \ab[20][21] , \ab[20][20] , \ab[20][19] ,
         \ab[20][18] , \ab[20][17] , \ab[20][16] , \ab[20][15] , \ab[20][14] ,
         \ab[20][13] , \ab[20][12] , \ab[20][11] , \ab[20][10] , \ab[20][9] ,
         \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][5] , \ab[20][4] ,
         \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] , \ab[19][31] ,
         \ab[19][30] , \ab[19][29] , \ab[19][28] , \ab[19][27] , \ab[19][26] ,
         \ab[19][25] , \ab[19][24] , \ab[19][23] , \ab[19][22] , \ab[19][21] ,
         \ab[19][20] , \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] ,
         \ab[19][15] , \ab[19][14] , \ab[19][13] , \ab[19][12] , \ab[19][11] ,
         \ab[19][10] , \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] ,
         \ab[19][5] , \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] ,
         \ab[19][0] , \ab[18][31] , \ab[18][30] , \ab[18][29] , \ab[18][28] ,
         \ab[18][27] , \ab[18][26] , \ab[18][25] , \ab[18][24] , \ab[18][23] ,
         \ab[18][22] , \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] ,
         \ab[18][17] , \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] ,
         \ab[18][12] , \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] ,
         \ab[18][7] , \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] ,
         \ab[18][2] , \ab[18][1] , \ab[18][0] , \ab[17][31] , \ab[17][30] ,
         \ab[17][29] , \ab[17][28] , \ab[17][27] , \ab[17][26] , \ab[17][25] ,
         \ab[17][24] , \ab[17][23] , \ab[17][22] , \ab[17][21] , \ab[17][20] ,
         \ab[17][19] , \ab[17][18] , \ab[17][17] , \ab[17][16] , \ab[17][15] ,
         \ab[17][14] , \ab[17][13] , \ab[17][12] , \ab[17][11] , \ab[17][10] ,
         \ab[17][9] , \ab[17][8] , \ab[17][7] , \ab[17][6] , \ab[17][5] ,
         \ab[17][4] , \ab[17][3] , \ab[17][2] , \ab[17][1] , \ab[17][0] ,
         \ab[16][31] , \ab[16][30] , \ab[16][29] , \ab[16][28] , \ab[16][27] ,
         \ab[16][26] , \ab[16][25] , \ab[16][24] , \ab[16][23] , \ab[16][22] ,
         \ab[16][21] , \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] ,
         \ab[16][16] , \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] ,
         \ab[16][11] , \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] ,
         \ab[16][6] , \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] ,
         \ab[16][1] , \ab[16][0] , \ab[15][31] , \ab[15][30] , \ab[15][29] ,
         \ab[15][28] , \ab[15][27] , \ab[15][26] , \ab[15][25] , \ab[15][24] ,
         \ab[15][23] , \ab[15][22] , \ab[15][21] , \ab[15][20] , \ab[15][19] ,
         \ab[15][18] , \ab[15][17] , \ab[15][16] , \ab[15][15] , \ab[15][14] ,
         \ab[15][13] , \ab[15][12] , \ab[15][11] , \ab[15][10] , \ab[15][9] ,
         \ab[15][8] , \ab[15][7] , \ab[15][6] , \ab[15][5] , \ab[15][4] ,
         \ab[15][3] , \ab[15][2] , \ab[15][1] , \ab[15][0] , \ab[14][31] ,
         \ab[14][30] , \ab[14][29] , \ab[14][28] , \ab[14][27] , \ab[14][26] ,
         \ab[14][25] , \ab[14][24] , \ab[14][23] , \ab[14][22] , \ab[14][21] ,
         \ab[14][20] , \ab[14][19] , \ab[14][18] , \ab[14][17] , \ab[14][16] ,
         \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] ,
         \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] ,
         \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] ,
         \ab[14][0] , \ab[13][31] , \ab[13][30] , \ab[13][29] , \ab[13][28] ,
         \ab[13][27] , \ab[13][26] , \ab[13][25] , \ab[13][24] , \ab[13][23] ,
         \ab[13][22] , \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] ,
         \ab[13][17] , \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][31] , \ab[12][30] ,
         \ab[12][29] , \ab[12][28] , \ab[12][27] , \ab[12][26] , \ab[12][25] ,
         \ab[12][24] , \ab[12][23] , \ab[12][22] , \ab[12][21] , \ab[12][20] ,
         \ab[12][19] , \ab[12][18] , \ab[12][17] , \ab[12][16] , \ab[12][15] ,
         \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] ,
         \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] ,
         \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][31] , \ab[11][30] , \ab[11][29] , \ab[11][28] , \ab[11][27] ,
         \ab[11][26] , \ab[11][25] , \ab[11][24] , \ab[11][23] , \ab[11][22] ,
         \ab[11][21] , \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] ,
         \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] ,
         \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] ,
         \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] ,
         \ab[11][1] , \ab[11][0] , \ab[10][31] , \ab[10][30] , \ab[10][29] ,
         \ab[10][28] , \ab[10][27] , \ab[10][26] , \ab[10][25] , \ab[10][24] ,
         \ab[10][23] , \ab[10][22] , \ab[10][21] , \ab[10][20] , \ab[10][19] ,
         \ab[10][18] , \ab[10][17] , \ab[10][16] , \ab[10][15] , \ab[10][14] ,
         \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] ,
         \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] ,
         \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][31] ,
         \ab[9][30] , \ab[9][29] , \ab[9][28] , \ab[9][27] , \ab[9][26] ,
         \ab[9][25] , \ab[9][24] , \ab[9][23] , \ab[9][22] , \ab[9][21] ,
         \ab[9][20] , \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] ,
         \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] ,
         \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] ,
         \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] ,
         \ab[9][0] , \ab[8][31] , \ab[8][30] , \ab[8][29] , \ab[8][28] ,
         \ab[8][27] , \ab[8][26] , \ab[8][25] , \ab[8][24] , \ab[8][23] ,
         \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] ,
         \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][31] , \ab[7][30] ,
         \ab[7][29] , \ab[7][28] , \ab[7][27] , \ab[7][26] , \ab[7][25] ,
         \ab[7][24] , \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] ,
         \ab[7][19] , \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][31] , \ab[6][30] , \ab[6][29] , \ab[6][28] , \ab[6][27] ,
         \ab[6][26] , \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] ,
         \ab[6][21] , \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] ,
         \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] ,
         \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] ,
         \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] ,
         \ab[6][1] , \ab[6][0] , \ab[5][31] , \ab[5][30] , \ab[5][29] ,
         \ab[5][28] , \ab[5][27] , \ab[5][26] , \ab[5][25] , \ab[5][24] ,
         \ab[5][23] , \ab[5][22] , \ab[5][21] , \ab[5][20] , \ab[5][19] ,
         \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][15] , \ab[5][14] ,
         \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] ,
         \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] ,
         \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][31] ,
         \ab[4][30] , \ab[4][29] , \ab[4][28] , \ab[4][27] , \ab[4][26] ,
         \ab[4][25] , \ab[4][24] , \ab[4][23] , \ab[4][22] , \ab[4][21] ,
         \ab[4][20] , \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] ,
         \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] ,
         \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] ,
         \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] ,
         \ab[4][0] , \ab[3][31] , \ab[3][30] , \ab[3][29] , \ab[3][28] ,
         \ab[3][27] , \ab[3][26] , \ab[3][25] , \ab[3][24] , \ab[3][23] ,
         \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] ,
         \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][31] , \ab[2][30] ,
         \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] , \ab[2][25] ,
         \ab[2][24] , \ab[2][23] , \ab[2][22] , \ab[2][21] , \ab[2][20] ,
         \ab[2][19] , \ab[2][18] , \ab[2][17] , \ab[2][16] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][31] , \ab[1][30] , \ab[1][29] , \ab[1][28] , \ab[1][27] ,
         \ab[1][26] , \ab[1][25] , \ab[1][24] , \ab[1][23] , \ab[1][22] ,
         \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] ,
         \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] ,
         \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] ,
         \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] ,
         \ab[1][1] , \ab[1][0] , \ab[0][31] , \ab[0][30] , \ab[0][29] ,
         \ab[0][28] , \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] ,
         \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] ,
         \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[15][30] ,
         \CARRYB[15][29] , \CARRYB[15][28] , \CARRYB[15][27] ,
         \CARRYB[15][26] , \CARRYB[15][25] , \CARRYB[15][24] ,
         \CARRYB[15][23] , \CARRYB[15][22] , \CARRYB[15][21] ,
         \CARRYB[15][20] , \CARRYB[15][19] , \CARRYB[15][18] ,
         \CARRYB[15][17] , \CARRYB[15][16] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][30] , \CARRYB[13][29] , \CARRYB[13][28] ,
         \CARRYB[13][27] , \CARRYB[13][26] , \CARRYB[13][25] ,
         \CARRYB[13][24] , \CARRYB[13][23] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][30] , \CARRYB[11][29] , \CARRYB[11][28] ,
         \CARRYB[11][27] , \CARRYB[11][26] , \CARRYB[11][25] ,
         \CARRYB[11][24] , \CARRYB[11][23] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][30] , \CARRYB[10][29] , \CARRYB[10][28] ,
         \CARRYB[10][27] , \CARRYB[10][26] , \CARRYB[10][25] ,
         \CARRYB[10][24] , \CARRYB[10][23] , \CARRYB[10][22] ,
         \CARRYB[10][21] , \CARRYB[10][20] , \CARRYB[10][19] ,
         \CARRYB[10][18] , \CARRYB[10][17] , \CARRYB[10][16] ,
         \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][30] , \CARRYB[9][29] , \CARRYB[9][28] ,
         \CARRYB[9][27] , \CARRYB[9][26] , \CARRYB[9][25] , \CARRYB[9][24] ,
         \CARRYB[9][23] , \CARRYB[9][22] , \CARRYB[9][21] , \CARRYB[9][20] ,
         \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] , \CARRYB[9][16] ,
         \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] ,
         \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] ,
         \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] ,
         \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] ,
         \CARRYB[8][30] , \CARRYB[8][29] , \CARRYB[8][28] , \CARRYB[8][27] ,
         \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] , \CARRYB[8][23] ,
         \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] , \CARRYB[8][19] ,
         \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] , \CARRYB[8][15] ,
         \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] ,
         \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] ,
         \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] ,
         \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][30] ,
         \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] , \CARRYB[7][26] ,
         \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] ,
         \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] ,
         \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][30] , \CARRYB[6][29] ,
         \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][30] , \CARRYB[5][29] , \CARRYB[5][28] ,
         \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] , \CARRYB[5][24] ,
         \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] , \CARRYB[5][20] ,
         \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] , \CARRYB[5][16] ,
         \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] ,
         \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] ,
         \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] ,
         \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] ,
         \CARRYB[4][30] , \CARRYB[4][29] , \CARRYB[4][28] , \CARRYB[4][27] ,
         \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] , \CARRYB[4][23] ,
         \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] , \CARRYB[4][19] ,
         \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][15] ,
         \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] ,
         \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] ,
         \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] ,
         \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][30] ,
         \CARRYB[3][29] , \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] ,
         \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][30] , \CARRYB[2][29] ,
         \CARRYB[2][28] , \CARRYB[2][27] , \CARRYB[2][26] , \CARRYB[2][25] ,
         \CARRYB[2][24] , \CARRYB[2][23] , \CARRYB[2][22] , \CARRYB[2][21] ,
         \CARRYB[2][20] , \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] ,
         \CARRYB[2][16] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \SUMB[15][30] , \SUMB[15][29] , \SUMB[15][28] ,
         \SUMB[15][27] , \SUMB[15][26] , \SUMB[15][25] , \SUMB[15][24] ,
         \SUMB[15][23] , \SUMB[15][22] , \SUMB[15][21] , \SUMB[15][20] ,
         \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] , \SUMB[15][16] ,
         \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] ,
         \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] ,
         \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] ,
         \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][30] ,
         \SUMB[14][29] , \SUMB[14][28] , \SUMB[14][27] , \SUMB[14][26] ,
         \SUMB[14][25] , \SUMB[14][24] , \SUMB[14][23] , \SUMB[14][22] ,
         \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] , \SUMB[14][18] ,
         \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][30] , \SUMB[13][29] , \SUMB[13][28] ,
         \SUMB[13][27] , \SUMB[13][26] , \SUMB[13][25] , \SUMB[13][24] ,
         \SUMB[13][23] , \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] ,
         \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] ,
         \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][30] ,
         \SUMB[12][29] , \SUMB[12][28] , \SUMB[12][27] , \SUMB[12][26] ,
         \SUMB[12][25] , \SUMB[12][24] , \SUMB[12][23] , \SUMB[12][22] ,
         \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] ,
         \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][30] , \SUMB[11][29] , \SUMB[11][28] ,
         \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] ,
         \SUMB[11][23] , \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] ,
         \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][30] ,
         \SUMB[10][29] , \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] ,
         \SUMB[10][25] , \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] ,
         \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] ,
         \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][30] , \SUMB[9][29] , \SUMB[9][28] ,
         \SUMB[9][27] , \SUMB[9][26] , \SUMB[9][25] , \SUMB[9][24] ,
         \SUMB[9][23] , \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] ,
         \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] ,
         \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][30] , \SUMB[8][29] ,
         \SUMB[8][28] , \SUMB[8][27] , \SUMB[8][26] , \SUMB[8][25] ,
         \SUMB[8][24] , \SUMB[8][23] , \SUMB[8][22] , \SUMB[8][21] ,
         \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] , \SUMB[8][17] ,
         \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][30] ,
         \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] , \SUMB[7][26] ,
         \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][30] ,
         \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] , \SUMB[6][26] ,
         \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][30] ,
         \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] , \SUMB[5][26] ,
         \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][30] ,
         \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] , \SUMB[4][26] ,
         \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][30] ,
         \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][30] ,
         \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] ,
         \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[31][31] , \CARRYB[31][30] , \CARRYB[31][29] ,
         \CARRYB[31][28] , \CARRYB[31][27] , \CARRYB[31][26] ,
         \CARRYB[31][25] , \CARRYB[31][24] , \CARRYB[31][23] ,
         \CARRYB[31][22] , \CARRYB[31][21] , \CARRYB[31][20] ,
         \CARRYB[31][19] , \CARRYB[31][18] , \CARRYB[31][17] ,
         \CARRYB[31][16] , \CARRYB[31][15] , \CARRYB[31][14] ,
         \CARRYB[31][13] , \CARRYB[31][12] , \CARRYB[31][11] ,
         \CARRYB[31][10] , \CARRYB[31][9] , \CARRYB[31][8] , \CARRYB[31][7] ,
         \CARRYB[31][6] , \CARRYB[31][5] , \CARRYB[31][4] , \CARRYB[31][3] ,
         \CARRYB[31][2] , \CARRYB[31][1] , \CARRYB[31][0] , \CARRYB[30][30] ,
         \CARRYB[30][29] , \CARRYB[30][28] , \CARRYB[30][27] ,
         \CARRYB[30][26] , \CARRYB[30][25] , \CARRYB[30][24] ,
         \CARRYB[30][23] , \CARRYB[30][22] , \CARRYB[30][21] ,
         \CARRYB[30][20] , \CARRYB[30][19] , \CARRYB[30][18] ,
         \CARRYB[30][17] , \CARRYB[30][16] , \CARRYB[30][15] ,
         \CARRYB[30][14] , \CARRYB[30][13] , \CARRYB[30][12] ,
         \CARRYB[30][11] , \CARRYB[30][10] , \CARRYB[30][9] , \CARRYB[30][8] ,
         \CARRYB[30][7] , \CARRYB[30][6] , \CARRYB[30][5] , \CARRYB[30][4] ,
         \CARRYB[30][3] , \CARRYB[30][2] , \CARRYB[30][1] , \CARRYB[30][0] ,
         \CARRYB[29][30] , \CARRYB[29][29] , \CARRYB[29][28] ,
         \CARRYB[29][27] , \CARRYB[29][26] , \CARRYB[29][25] ,
         \CARRYB[29][24] , \CARRYB[29][23] , \CARRYB[29][22] ,
         \CARRYB[29][21] , \CARRYB[29][20] , \CARRYB[29][19] ,
         \CARRYB[29][18] , \CARRYB[29][17] , \CARRYB[29][16] ,
         \CARRYB[29][15] , \CARRYB[29][14] , \CARRYB[29][13] ,
         \CARRYB[29][12] , \CARRYB[29][11] , \CARRYB[29][10] , \CARRYB[29][9] ,
         \CARRYB[29][8] , \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][5] ,
         \CARRYB[29][4] , \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][30] , \CARRYB[28][29] , \CARRYB[28][28] ,
         \CARRYB[28][27] , \CARRYB[28][26] , \CARRYB[28][25] ,
         \CARRYB[28][24] , \CARRYB[28][23] , \CARRYB[28][22] ,
         \CARRYB[28][21] , \CARRYB[28][20] , \CARRYB[28][19] ,
         \CARRYB[28][18] , \CARRYB[28][17] , \CARRYB[28][16] ,
         \CARRYB[28][15] , \CARRYB[28][14] , \CARRYB[28][13] ,
         \CARRYB[28][12] , \CARRYB[28][11] , \CARRYB[28][10] , \CARRYB[28][9] ,
         \CARRYB[28][8] , \CARRYB[28][7] , \CARRYB[28][6] , \CARRYB[28][5] ,
         \CARRYB[28][4] , \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][30] , \CARRYB[27][29] , \CARRYB[27][28] ,
         \CARRYB[27][27] , \CARRYB[27][26] , \CARRYB[27][25] ,
         \CARRYB[27][24] , \CARRYB[27][23] , \CARRYB[27][22] ,
         \CARRYB[27][21] , \CARRYB[27][20] , \CARRYB[27][19] ,
         \CARRYB[27][18] , \CARRYB[27][17] , \CARRYB[27][16] ,
         \CARRYB[27][15] , \CARRYB[27][14] , \CARRYB[27][13] ,
         \CARRYB[27][12] , \CARRYB[27][11] , \CARRYB[27][10] , \CARRYB[27][9] ,
         \CARRYB[27][8] , \CARRYB[27][7] , \CARRYB[27][6] , \CARRYB[27][5] ,
         \CARRYB[27][4] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][30] , \CARRYB[25][29] , \CARRYB[25][28] ,
         \CARRYB[25][27] , \CARRYB[25][26] , \CARRYB[25][25] ,
         \CARRYB[25][24] , \CARRYB[25][23] , \CARRYB[25][22] ,
         \CARRYB[25][21] , \CARRYB[25][20] , \CARRYB[25][19] ,
         \CARRYB[25][18] , \CARRYB[25][17] , \CARRYB[25][16] ,
         \CARRYB[25][15] , \CARRYB[25][14] , \CARRYB[25][13] ,
         \CARRYB[25][12] , \CARRYB[25][11] , \CARRYB[25][10] , \CARRYB[25][9] ,
         \CARRYB[25][8] , \CARRYB[25][7] , \CARRYB[25][6] , \CARRYB[25][5] ,
         \CARRYB[25][4] , \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] ,
         \CARRYB[25][0] , \CARRYB[24][30] , \CARRYB[24][29] , \CARRYB[24][28] ,
         \CARRYB[24][27] , \CARRYB[24][26] , \CARRYB[24][25] ,
         \CARRYB[24][24] , \CARRYB[24][23] , \CARRYB[24][22] ,
         \CARRYB[24][21] , \CARRYB[24][20] , \CARRYB[24][19] ,
         \CARRYB[24][18] , \CARRYB[24][17] , \CARRYB[24][16] ,
         \CARRYB[24][15] , \CARRYB[24][14] , \CARRYB[24][13] ,
         \CARRYB[24][12] , \CARRYB[24][11] , \CARRYB[24][10] , \CARRYB[24][9] ,
         \CARRYB[24][8] , \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] ,
         \CARRYB[24][4] , \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] ,
         \CARRYB[24][0] , \CARRYB[23][30] , \CARRYB[23][29] , \CARRYB[23][28] ,
         \CARRYB[23][27] , \CARRYB[23][26] , \CARRYB[23][25] ,
         \CARRYB[23][24] , \CARRYB[23][23] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][30] , \CARRYB[22][29] , \CARRYB[22][28] ,
         \CARRYB[22][27] , \CARRYB[22][26] , \CARRYB[22][25] ,
         \CARRYB[22][24] , \CARRYB[22][23] , \CARRYB[22][22] ,
         \CARRYB[22][21] , \CARRYB[22][20] , \CARRYB[22][19] ,
         \CARRYB[22][18] , \CARRYB[22][17] , \CARRYB[22][16] ,
         \CARRYB[22][15] , \CARRYB[22][14] , \CARRYB[22][13] ,
         \CARRYB[22][12] , \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] ,
         \CARRYB[22][8] , \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][30] , \CARRYB[21][29] , \CARRYB[21][28] ,
         \CARRYB[21][27] , \CARRYB[21][26] , \CARRYB[21][25] ,
         \CARRYB[21][24] , \CARRYB[21][23] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][30] , \CARRYB[19][29] , \CARRYB[19][28] ,
         \CARRYB[19][27] , \CARRYB[19][26] , \CARRYB[19][25] ,
         \CARRYB[19][24] , \CARRYB[19][23] , \CARRYB[19][22] ,
         \CARRYB[19][21] , \CARRYB[19][20] , \CARRYB[19][19] ,
         \CARRYB[19][18] , \CARRYB[19][17] , \CARRYB[19][16] ,
         \CARRYB[19][15] , \CARRYB[19][14] , \CARRYB[19][13] ,
         \CARRYB[19][12] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] ,
         \CARRYB[19][8] , \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] ,
         \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] ,
         \CARRYB[19][0] , \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][30] , \CARRYB[17][29] , \CARRYB[17][28] ,
         \CARRYB[17][27] , \CARRYB[17][26] , \CARRYB[17][25] ,
         \CARRYB[17][24] , \CARRYB[17][23] , \CARRYB[17][22] ,
         \CARRYB[17][21] , \CARRYB[17][20] , \CARRYB[17][19] ,
         \CARRYB[17][18] , \CARRYB[17][17] , \CARRYB[17][16] ,
         \CARRYB[17][15] , \CARRYB[17][14] , \CARRYB[17][13] ,
         \CARRYB[17][12] , \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] ,
         \CARRYB[17][8] , \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \SUMB[31][31] , \SUMB[31][30] , \SUMB[31][29] ,
         \SUMB[31][28] , \SUMB[31][27] , \SUMB[31][26] , \SUMB[31][25] ,
         \SUMB[31][24] , \SUMB[31][23] , \SUMB[31][22] , \SUMB[31][21] ,
         \SUMB[31][20] , \SUMB[31][19] , \SUMB[31][18] , \SUMB[31][17] ,
         \SUMB[31][16] , \SUMB[31][15] , \SUMB[31][14] , \SUMB[31][13] ,
         \SUMB[31][12] , \SUMB[31][11] , \SUMB[31][10] , \SUMB[31][9] ,
         \SUMB[31][8] , \SUMB[31][7] , \SUMB[31][6] , \SUMB[31][5] ,
         \SUMB[31][4] , \SUMB[31][3] , \SUMB[31][2] , \SUMB[31][1] ,
         \SUMB[31][0] , \SUMB[30][30] , \SUMB[30][29] , \SUMB[30][28] ,
         \SUMB[30][27] , \SUMB[30][26] , \SUMB[30][25] , \SUMB[30][24] ,
         \SUMB[30][23] , \SUMB[30][22] , \SUMB[30][21] , \SUMB[30][20] ,
         \SUMB[30][19] , \SUMB[30][18] , \SUMB[30][17] , \SUMB[30][16] ,
         \SUMB[30][15] , \SUMB[30][14] , \SUMB[30][13] , \SUMB[30][12] ,
         \SUMB[30][11] , \SUMB[30][10] , \SUMB[30][9] , \SUMB[30][8] ,
         \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][5] , \SUMB[30][4] ,
         \SUMB[30][3] , \SUMB[30][2] , \SUMB[30][1] , \SUMB[29][30] ,
         \SUMB[29][29] , \SUMB[29][28] , \SUMB[29][27] , \SUMB[29][26] ,
         \SUMB[29][25] , \SUMB[29][24] , \SUMB[29][23] , \SUMB[29][22] ,
         \SUMB[29][21] , \SUMB[29][20] , \SUMB[29][19] , \SUMB[29][18] ,
         \SUMB[29][17] , \SUMB[29][16] , \SUMB[29][15] , \SUMB[29][14] ,
         \SUMB[29][13] , \SUMB[29][12] , \SUMB[29][11] , \SUMB[29][10] ,
         \SUMB[29][9] , \SUMB[29][8] , \SUMB[29][7] , \SUMB[29][6] ,
         \SUMB[29][5] , \SUMB[29][4] , \SUMB[29][3] , \SUMB[29][2] ,
         \SUMB[29][1] , \SUMB[28][30] , \SUMB[28][29] , \SUMB[28][28] ,
         \SUMB[28][27] , \SUMB[28][26] , \SUMB[28][25] , \SUMB[28][24] ,
         \SUMB[28][23] , \SUMB[28][22] , \SUMB[28][21] , \SUMB[28][20] ,
         \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] , \SUMB[28][16] ,
         \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] , \SUMB[28][12] ,
         \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] , \SUMB[28][8] ,
         \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] , \SUMB[28][4] ,
         \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][30] ,
         \SUMB[27][29] , \SUMB[27][28] , \SUMB[27][27] , \SUMB[27][26] ,
         \SUMB[27][25] , \SUMB[27][24] , \SUMB[27][23] , \SUMB[27][22] ,
         \SUMB[27][21] , \SUMB[27][20] , \SUMB[27][19] , \SUMB[27][18] ,
         \SUMB[27][17] , \SUMB[27][16] , \SUMB[27][15] , \SUMB[27][14] ,
         \SUMB[27][13] , \SUMB[27][12] , \SUMB[27][11] , \SUMB[27][10] ,
         \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] , \SUMB[27][6] ,
         \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] , \SUMB[27][2] ,
         \SUMB[27][1] , \SUMB[26][30] , \SUMB[26][29] , \SUMB[26][28] ,
         \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] , \SUMB[26][24] ,
         \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] , \SUMB[26][20] ,
         \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] , \SUMB[26][16] ,
         \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] , \SUMB[26][12] ,
         \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] , \SUMB[26][8] ,
         \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][30] ,
         \SUMB[25][29] , \SUMB[25][28] , \SUMB[25][27] , \SUMB[25][26] ,
         \SUMB[25][25] , \SUMB[25][24] , \SUMB[25][23] , \SUMB[25][22] ,
         \SUMB[25][21] , \SUMB[25][20] , \SUMB[25][19] , \SUMB[25][18] ,
         \SUMB[25][17] , \SUMB[25][16] , \SUMB[25][15] , \SUMB[25][14] ,
         \SUMB[25][13] , \SUMB[25][12] , \SUMB[25][11] , \SUMB[25][10] ,
         \SUMB[25][9] , \SUMB[25][8] , \SUMB[25][7] , \SUMB[25][6] ,
         \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] ,
         \SUMB[25][1] , \SUMB[24][30] , \SUMB[24][29] , \SUMB[24][28] ,
         \SUMB[24][27] , \SUMB[24][26] , \SUMB[24][25] , \SUMB[24][24] ,
         \SUMB[24][23] , \SUMB[24][22] , \SUMB[24][21] , \SUMB[24][20] ,
         \SUMB[24][19] , \SUMB[24][18] , \SUMB[24][17] , \SUMB[24][16] ,
         \SUMB[24][15] , \SUMB[24][14] , \SUMB[24][13] , \SUMB[24][12] ,
         \SUMB[24][11] , \SUMB[24][10] , \SUMB[24][9] , \SUMB[24][8] ,
         \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][30] ,
         \SUMB[23][29] , \SUMB[23][28] , \SUMB[23][27] , \SUMB[23][26] ,
         \SUMB[23][25] , \SUMB[23][24] , \SUMB[23][23] , \SUMB[23][22] ,
         \SUMB[23][21] , \SUMB[23][20] , \SUMB[23][19] , \SUMB[23][18] ,
         \SUMB[23][17] , \SUMB[23][16] , \SUMB[23][15] , \SUMB[23][14] ,
         \SUMB[23][13] , \SUMB[23][12] , \SUMB[23][11] , \SUMB[23][10] ,
         \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] , \SUMB[23][6] ,
         \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] ,
         \SUMB[23][1] , \SUMB[22][30] , \SUMB[22][29] , \SUMB[22][28] ,
         \SUMB[22][27] , \SUMB[22][26] , \SUMB[22][25] , \SUMB[22][24] ,
         \SUMB[22][23] , \SUMB[22][22] , \SUMB[22][21] , \SUMB[22][20] ,
         \SUMB[22][19] , \SUMB[22][18] , \SUMB[22][17] , \SUMB[22][16] ,
         \SUMB[22][15] , \SUMB[22][14] , \SUMB[22][13] , \SUMB[22][12] ,
         \SUMB[22][11] , \SUMB[22][10] , \SUMB[22][9] , \SUMB[22][8] ,
         \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] ,
         \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][30] ,
         \SUMB[21][29] , \SUMB[21][28] , \SUMB[21][27] , \SUMB[21][26] ,
         \SUMB[21][25] , \SUMB[21][24] , \SUMB[21][23] , \SUMB[21][22] ,
         \SUMB[21][21] , \SUMB[21][20] , \SUMB[21][19] , \SUMB[21][18] ,
         \SUMB[21][17] , \SUMB[21][16] , \SUMB[21][15] , \SUMB[21][14] ,
         \SUMB[21][13] , \SUMB[21][12] , \SUMB[21][11] , \SUMB[21][10] ,
         \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] , \SUMB[21][6] ,
         \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] ,
         \SUMB[21][1] , \SUMB[20][30] , \SUMB[20][29] , \SUMB[20][28] ,
         \SUMB[20][27] , \SUMB[20][26] , \SUMB[20][25] , \SUMB[20][24] ,
         \SUMB[20][23] , \SUMB[20][22] , \SUMB[20][21] , \SUMB[20][20] ,
         \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] , \SUMB[20][16] ,
         \SUMB[20][15] , \SUMB[20][14] , \SUMB[20][13] , \SUMB[20][12] ,
         \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] ,
         \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][30] ,
         \SUMB[19][29] , \SUMB[19][28] , \SUMB[19][27] , \SUMB[19][26] ,
         \SUMB[19][25] , \SUMB[19][24] , \SUMB[19][23] , \SUMB[19][22] ,
         \SUMB[19][21] , \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] ,
         \SUMB[19][17] , \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] ,
         \SUMB[19][13] , \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] ,
         \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][30] , \SUMB[18][29] , \SUMB[18][28] ,
         \SUMB[18][27] , \SUMB[18][26] , \SUMB[18][25] , \SUMB[18][24] ,
         \SUMB[18][23] , \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] ,
         \SUMB[18][19] , \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] ,
         \SUMB[18][15] , \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] ,
         \SUMB[18][11] , \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] ,
         \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] ,
         \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][30] ,
         \SUMB[17][29] , \SUMB[17][28] , \SUMB[17][27] , \SUMB[17][26] ,
         \SUMB[17][25] , \SUMB[17][24] , \SUMB[17][23] , \SUMB[17][22] ,
         \SUMB[17][21] , \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] ,
         \SUMB[17][17] , \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] ,
         \SUMB[17][13] , \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] ,
         \SUMB[17][9] , \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] ,
         \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] ,
         \SUMB[17][1] , \SUMB[16][30] , \SUMB[16][29] , \SUMB[16][28] ,
         \SUMB[16][27] , \SUMB[16][26] , \SUMB[16][25] , \SUMB[16][24] ,
         \SUMB[16][23] , \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] ,
         \SUMB[16][19] , \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] ,
         \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] ,
         \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] ,
         \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , ZA, ZB, \A1[60] ,
         \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] ,
         \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] ,
         \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] ,
         \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] ,
         \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] ,
         \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] ,
         \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] ,
         \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] ,
         \A1[3] , \A1[2] , \A1[1] , \A1[0] , \A2[30] , n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239;
  assign ZA = A[31];
  assign ZB = B[31];

  FADDX1 S4_1 ( .A(\ab[31][1] ), .B(\CARRYB[30][1] ), .CI(\SUMB[30][2] ), .CO(
        \CARRYB[31][1] ), .S(\SUMB[31][1] ) );
  FADDX1 S4_5 ( .A(\ab[31][5] ), .B(\CARRYB[30][5] ), .CI(\SUMB[30][6] ), .CO(
        \CARRYB[31][5] ), .S(\SUMB[31][5] ) );
  FADDX1 S4_6 ( .A(\ab[31][6] ), .B(\CARRYB[30][6] ), .CI(\SUMB[30][7] ), .CO(
        \CARRYB[31][6] ), .S(\SUMB[31][6] ) );
  FADDX1 S4_12 ( .A(\ab[31][12] ), .B(\CARRYB[30][12] ), .CI(\SUMB[30][13] ), 
        .CO(\CARRYB[31][12] ), .S(\SUMB[31][12] ) );
  FADDX1 S4_13 ( .A(\ab[31][13] ), .B(\CARRYB[30][13] ), .CI(\SUMB[30][14] ), 
        .CO(\CARRYB[31][13] ), .S(\SUMB[31][13] ) );
  FADDX1 S4_14 ( .A(\ab[31][14] ), .B(\CARRYB[30][14] ), .CI(\SUMB[30][15] ), 
        .CO(\CARRYB[31][14] ), .S(\SUMB[31][14] ) );
  FADDX1 S4_15 ( .A(\ab[31][15] ), .B(\CARRYB[30][15] ), .CI(\SUMB[30][16] ), 
        .CO(\CARRYB[31][15] ), .S(\SUMB[31][15] ) );
  FADDX1 S4_16 ( .A(\ab[31][16] ), .B(\CARRYB[30][16] ), .CI(\SUMB[30][17] ), 
        .CO(\CARRYB[31][16] ), .S(\SUMB[31][16] ) );
  FADDX1 S4_17 ( .A(\ab[31][17] ), .B(\CARRYB[30][17] ), .CI(\SUMB[30][18] ), 
        .CO(\CARRYB[31][17] ), .S(\SUMB[31][17] ) );
  FADDX1 S4_18 ( .A(\ab[31][18] ), .B(\CARRYB[30][18] ), .CI(\SUMB[30][19] ), 
        .CO(\CARRYB[31][18] ), .S(\SUMB[31][18] ) );
  FADDX1 S4_19 ( .A(\ab[31][19] ), .B(\CARRYB[30][19] ), .CI(\SUMB[30][20] ), 
        .CO(\CARRYB[31][19] ), .S(\SUMB[31][19] ) );
  FADDX1 S4_20 ( .A(\ab[31][20] ), .B(\CARRYB[30][20] ), .CI(\SUMB[30][21] ), 
        .CO(\CARRYB[31][20] ), .S(\SUMB[31][20] ) );
  FADDX1 S4_23 ( .A(\ab[31][23] ), .B(\CARRYB[30][23] ), .CI(\SUMB[30][24] ), 
        .CO(\CARRYB[31][23] ), .S(\SUMB[31][23] ) );
  FADDX1 S4_26 ( .A(\ab[31][26] ), .B(\CARRYB[30][26] ), .CI(\SUMB[30][27] ), 
        .CO(\CARRYB[31][26] ), .S(\SUMB[31][26] ) );
  FADDX1 S4_27 ( .A(\ab[31][27] ), .B(\CARRYB[30][27] ), .CI(\SUMB[30][28] ), 
        .CO(\CARRYB[31][27] ), .S(\SUMB[31][27] ) );
  FADDX1 S4_28 ( .A(\ab[31][28] ), .B(\CARRYB[30][28] ), .CI(\SUMB[30][29] ), 
        .CO(\CARRYB[31][28] ), .S(\SUMB[31][28] ) );
  FADDX1 S4_29 ( .A(\ab[31][29] ), .B(\CARRYB[30][29] ), .CI(\SUMB[30][30] ), 
        .CO(\CARRYB[31][29] ), .S(\SUMB[31][29] ) );
  FADDX1 S5_30 ( .A(\ab[31][30] ), .B(\CARRYB[30][30] ), .CI(\ab[30][31] ), 
        .CO(\CARRYB[31][30] ), .S(\SUMB[31][30] ) );
  FADDX1 S14_31 ( .A(n2004), .B(n2094), .CI(\ab[31][31] ), .CO(
        \CARRYB[31][31] ), .S(\SUMB[31][31] ) );
  FADDX1 S2_30_5 ( .A(\ab[30][5] ), .B(\CARRYB[29][5] ), .CI(\SUMB[29][6] ), 
        .CO(\CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FADDX1 S2_30_9 ( .A(\ab[30][9] ), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), 
        .CO(\CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FADDX1 S2_30_13 ( .A(\ab[30][13] ), .B(\CARRYB[29][13] ), .CI(\SUMB[29][14] ), .CO(\CARRYB[30][13] ), .S(\SUMB[30][13] ) );
  FADDX1 S2_30_15 ( .A(\ab[30][15] ), .B(\CARRYB[29][15] ), .CI(\SUMB[29][16] ), .CO(\CARRYB[30][15] ), .S(\SUMB[30][15] ) );
  FADDX1 S2_30_19 ( .A(\ab[30][19] ), .B(\CARRYB[29][19] ), .CI(\SUMB[29][20] ), .CO(\CARRYB[30][19] ), .S(\SUMB[30][19] ) );
  FADDX1 S2_30_26 ( .A(\ab[30][26] ), .B(\CARRYB[29][26] ), .CI(\SUMB[29][27] ), .CO(\CARRYB[30][26] ), .S(\SUMB[30][26] ) );
  FADDX1 S2_30_27 ( .A(\ab[30][27] ), .B(\CARRYB[29][27] ), .CI(\SUMB[29][28] ), .CO(\CARRYB[30][27] ), .S(\SUMB[30][27] ) );
  FADDX1 S2_30_28 ( .A(\ab[30][28] ), .B(\CARRYB[29][28] ), .CI(\SUMB[29][29] ), .CO(\CARRYB[30][28] ), .S(\SUMB[30][28] ) );
  FADDX1 S2_30_29 ( .A(\ab[30][29] ), .B(\CARRYB[29][29] ), .CI(\SUMB[29][30] ), .CO(\CARRYB[30][29] ), .S(\SUMB[30][29] ) );
  FADDX1 S3_30_30 ( .A(\ab[30][30] ), .B(\CARRYB[29][30] ), .CI(\ab[29][31] ), 
        .CO(\CARRYB[30][30] ), .S(\SUMB[30][30] ) );
  FADDX1 S2_29_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), 
        .CO(\CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FADDX1 S2_29_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), 
        .CO(\CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FADDX1 S2_29_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FADDX1 S2_29_11 ( .A(\ab[29][11] ), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), .CO(\CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FADDX1 S2_29_13 ( .A(\ab[29][13] ), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), .CO(\CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FADDX1 S2_29_24 ( .A(\ab[29][24] ), .B(\CARRYB[28][24] ), .CI(\SUMB[28][25] ), .CO(\CARRYB[29][24] ), .S(\SUMB[29][24] ) );
  FADDX1 S2_29_25 ( .A(\ab[29][25] ), .B(\CARRYB[28][25] ), .CI(\SUMB[28][26] ), .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FADDX1 S2_29_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FADDX1 S2_29_29 ( .A(\ab[29][29] ), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), .CO(\CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FADDX1 S3_29_30 ( .A(\ab[29][30] ), .B(\CARRYB[28][30] ), .CI(\ab[28][31] ), 
        .CO(\CARRYB[29][30] ), .S(\SUMB[29][30] ) );
  FADDX1 S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(\A1[26] ) );
  FADDX1 S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FADDX1 S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FADDX1 S2_28_24 ( .A(\ab[28][24] ), .B(\CARRYB[27][24] ), .CI(\SUMB[27][25] ), .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FADDX1 S2_28_25 ( .A(\ab[28][25] ), .B(\CARRYB[27][25] ), .CI(\SUMB[27][26] ), .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FADDX1 S2_28_29 ( .A(\ab[28][29] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FADDX1 S3_28_30 ( .A(\ab[28][30] ), .B(\CARRYB[27][30] ), .CI(\ab[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FADDX1 S2_27_8 ( .A(\ab[27][8] ), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FADDX1 S2_27_12 ( .A(\ab[27][12] ), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), .CO(\CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FADDX1 S2_27_22 ( .A(\ab[27][22] ), .B(\CARRYB[26][22] ), .CI(\SUMB[26][23] ), .CO(\CARRYB[27][22] ), .S(\SUMB[27][22] ) );
  FADDX1 S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FADDX1 S2_27_28 ( .A(\ab[27][28] ), .B(\CARRYB[26][28] ), .CI(\SUMB[26][29] ), .CO(\CARRYB[27][28] ), .S(\SUMB[27][28] ) );
  FADDX1 S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(\A1[24] ) );
  FADDX1 S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FADDX1 S2_26_8 ( .A(\ab[26][8] ), .B(\CARRYB[25][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FADDX1 S2_26_9 ( .A(\ab[26][9] ), .B(\CARRYB[25][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FADDX1 S2_26_12 ( .A(\SUMB[25][13] ), .B(\ab[26][12] ), .CI(\CARRYB[25][12] ), .CO(\CARRYB[26][12] ), .S(\SUMB[26][12] ) );
  FADDX1 S2_26_13 ( .A(\ab[26][13] ), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), .CO(\CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FADDX1 S2_26_29 ( .A(\ab[26][29] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FADDX1 S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(\A1[23] ) );
  FADDX1 S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FADDX1 S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FADDX1 S2_25_8 ( .A(\ab[25][8] ), .B(\CARRYB[24][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FADDX1 S2_25_9 ( .A(\ab[25][9] ), .B(\CARRYB[24][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FADDX1 S2_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FADDX1 S2_25_12 ( .A(\ab[25][12] ), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), .CO(\CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FADDX1 S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FADDX1 S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FADDX1 S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FADDX1 S2_25_27 ( .A(\ab[25][27] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FADDX1 S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FADDX1 S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FADDX1 S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FADDX1 S2_24_9 ( .A(\ab[24][9] ), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FADDX1 S2_24_11 ( .A(\ab[24][11] ), .B(\CARRYB[23][11] ), .CI(\SUMB[23][12] ), .CO(\CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FADDX1 S2_24_13 ( .A(\ab[24][13] ), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), .CO(\CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FADDX1 S2_24_15 ( .A(\CARRYB[23][15] ), .B(\ab[24][15] ), .CI(\SUMB[23][16] ), .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FADDX1 S3_24_30 ( .A(\ab[24][30] ), .B(\CARRYB[23][30] ), .CI(\ab[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FADDX1 S2_23_6 ( .A(\CARRYB[22][6] ), .B(\ab[23][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FADDX1 S2_23_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FADDX1 S2_23_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FADDX1 S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FADDX1 S3_23_30 ( .A(\ab[23][30] ), .B(\CARRYB[22][30] ), .CI(\ab[22][31] ), 
        .CO(\CARRYB[23][30] ), .S(\SUMB[23][30] ) );
  FADDX1 S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FADDX1 S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FADDX1 S2_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FADDX1 S2_22_25 ( .A(\ab[22][25] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FADDX1 S2_22_26 ( .A(\ab[22][26] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FADDX1 S3_22_30 ( .A(\ab[22][30] ), .B(\CARRYB[21][30] ), .CI(\ab[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FADDX1 S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FADDX1 S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FADDX1 S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FADDX1 S2_21_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FADDX1 S2_21_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FADDX1 S2_21_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FADDX1 S3_21_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\ab[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FADDX1 S1_20_0 ( .A(\ab[20][0] ), .B(\SUMB[19][1] ), .CI(\CARRYB[19][0] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FADDX1 S2_20_8 ( .A(\CARRYB[19][8] ), .B(\ab[20][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FADDX1 S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FADDX1 S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FADDX1 S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FADDX1 S3_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\ab[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FADDX1 S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FADDX1 S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FADDX1 S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FADDX1 S3_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\ab[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FADDX1 S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FADDX1 S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FADDX1 S3_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\ab[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FADDX1 S2_17_14 ( .A(\ab[17][14] ), .B(\SUMB[16][15] ), .CI(\CARRYB[16][14] ), .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FADDX1 S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FADDX1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FADDX1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FADDX1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FADDX1 S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FADDX1 S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FADDX1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FADDX1 S2_15_12 ( .A(\CARRYB[14][12] ), .B(\ab[15][12] ), .CI(\SUMB[14][13] ), .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FADDX1 S3_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\ab[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FADDX1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FADDX1 S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FADDX1 S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FADDX1 S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FADDX1 S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FADDX1 S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FADDX1 S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FADDX1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FADDX1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FADDX1 S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FADDX1 S3_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\ab[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FADDX1 S2_11_19 ( .A(\CARRYB[10][19] ), .B(\ab[11][19] ), .CI(\SUMB[10][20] ), .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FADDX1 S2_11_24 ( .A(\CARRYB[10][24] ), .B(\ab[11][24] ), .CI(\SUMB[10][25] ), .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FADDX1 S2_11_25 ( .A(\CARRYB[10][25] ), .B(\ab[11][25] ), .CI(\SUMB[10][26] ), .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FADDX1 S3_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\ab[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FADDX1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), 
        .CO(\CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FADDX1 S3_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\ab[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FADDX1 S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FADDX1 S3_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\ab[8][31] ), 
        .CO(\CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FADDX1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FADDX1 S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FADDX1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FADDX1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FADDX1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FADDX1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FADDX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FADDX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FADDX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FADDX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FADDX1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FADDX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FADDX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FADDX1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FADDX1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FADDX1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FADDX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FADDX1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FADDX1 S2_2_1 ( .A(\ab[2][1] ), .B(n4), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FADDX1 S2_2_3 ( .A(\ab[2][3] ), .B(n1808), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FADDX1 S2_2_4 ( .A(\ab[2][4] ), .B(n3), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FADDX1 S2_2_5 ( .A(\SUMB[1][6] ), .B(n754), .CI(\ab[2][5] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FADDX1 S2_2_9 ( .A(\ab[2][9] ), .B(n1782), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FADDX1 S2_2_16 ( .A(\ab[2][16] ), .B(n294), .CI(\SUMB[1][17] ), .CO(
        \CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FADDX1 S2_2_19 ( .A(\ab[2][19] ), .B(n6), .CI(\SUMB[1][20] ), .CO(
        \CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FADDX1 S2_2_26 ( .A(\ab[2][26] ), .B(n165), .CI(\SUMB[1][27] ), .CO(
        \CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  VerilogMultiplier_DW01_add_0 FS_1 ( .A({n2175, \A1[60] , \A1[59] , \A1[58] , 
        \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , 
        \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , 
        \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , 
        \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , 
        \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , 
        \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , 
        \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , 
        \A1[0] }), .B({n16, n1987, n1994, n1999, n2001, n2000, n1998, n1997, 
        n1996, n1995, n1993, n1992, n1991, n1990, n1989, n1988, n1980, n1979, 
        n1983, n1972, n1985, n1976, n1981, n1975, n1973, n1978, n1982, n1974, 
        n1986, n1977, n1984, \A2[30] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[63:2]) );
  FADDX1 S4_2 ( .A(\ab[31][2] ), .B(\CARRYB[30][2] ), .CI(\SUMB[30][3] ), .CO(
        \CARRYB[31][2] ), .S(\SUMB[31][2] ) );
  FADDX1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FADDX1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FADDX1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FADDX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FADDX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FADDX1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FADDX1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FADDX1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FADDX1 S1_29_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), 
        .CO(\CARRYB[29][0] ), .S(\A1[27] ) );
  FADDX1 S2_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FADDX1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FADDX1 S1_2_0 ( .A(\ab[2][0] ), .B(n13), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FADDX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FADDX1 S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FADDX1 S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FADDX1 S2_25_11 ( .A(\ab[25][11] ), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), .CO(\CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FADDX1 S2_27_11 ( .A(\CARRYB[26][11] ), .B(\ab[27][11] ), .CI(\SUMB[26][12] ), .CO(\CARRYB[27][11] ), .S(\SUMB[27][11] ) );
  FADDX1 S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FADDX1 S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FADDX1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FADDX1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FADDX2 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FADDX1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FADDX1 S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FADDX1 S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FADDX1 S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FADDX1 S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FADDX1 S2_23_15 ( .A(\CARRYB[22][15] ), .B(\ab[23][15] ), .CI(\SUMB[22][16] ), .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FADDX1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), 
        .CO(\CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FADDX1 S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FADDX1 S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FADDX1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FADDX1 S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FADDX1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FADDX1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FADDX1 S2_26_7 ( .A(\ab[26][7] ), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FADDX1 S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FADDX1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FADDX1 S2_2_11 ( .A(\ab[2][11] ), .B(n1689), .CI(\SUMB[1][12] ), .CO(
        \CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FADDX1 S2_26_27 ( .A(\ab[26][27] ), .B(\CARRYB[25][27] ), .CI(\SUMB[25][28] ), .CO(\CARRYB[26][27] ), .S(\SUMB[26][27] ) );
  FADDX1 S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FADDX2 S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FADDX1 S2_8_15 ( .A(\SUMB[7][16] ), .B(\ab[8][15] ), .CI(\CARRYB[7][15] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FADDX1 S2_21_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FADDX1 S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FADDX2 S2_23_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FADDX1 S2_22_10 ( .A(\CARRYB[21][10] ), .B(\ab[22][10] ), .CI(\SUMB[21][11] ), .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FADDX1 S2_24_10 ( .A(\ab[24][10] ), .B(\CARRYB[23][10] ), .CI(\SUMB[23][11] ), .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FADDX1 S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FADDX1 S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FADDX1 S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FADDX1 S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FADDX1 S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FADDX1 S2_24_27 ( .A(\ab[24][27] ), .B(\CARRYB[23][27] ), .CI(\SUMB[23][28] ), .CO(\CARRYB[24][27] ), .S(\SUMB[24][27] ) );
  FADDX1 S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FADDX1 S2_12_15 ( .A(\CARRYB[11][15] ), .B(\ab[12][15] ), .CI(\SUMB[11][16] ), .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FADDX1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FADDX1 S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FADDX1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FADDX1 S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FADDX1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FADDX1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FADDX1 S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FADDX1 S2_28_21 ( .A(\ab[28][21] ), .B(\CARRYB[27][21] ), .CI(\SUMB[27][22] ), .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FADDX1 S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FADDX1 S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FADDX1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), 
        .CO(\CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FADDX1 S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FADDX1 S2_27_21 ( .A(\ab[27][21] ), .B(\CARRYB[26][21] ), .CI(\SUMB[26][22] ), .CO(\CARRYB[27][21] ), .S(\SUMB[27][21] ) );
  FADDX1 S2_21_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FADDX1 S2_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\SUMB[27][21] ), .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FADDX1 S2_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\SUMB[25][21] ), .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FADDX1 S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FADDX1 S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FADDX1 S2_7_8 ( .A(\ab[7][8] ), .B(\SUMB[6][9] ), .CI(\CARRYB[6][8] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FADDX1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FADDX1 S2_16_1 ( .A(\CARRYB[15][1] ), .B(\ab[16][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FADDX1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FADDX1 S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FADDX1 S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FADDX1 S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FADDX1 S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FADDX1 S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FADDX1 S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FADDX1 S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FADDX1 S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FADDX1 S2_9_20 ( .A(\CARRYB[8][20] ), .B(\ab[9][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FADDX1 S2_26_11 ( .A(\ab[26][11] ), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), .CO(\CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FADDX2 S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FADDX1 S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FADDX2 S3_3_30 ( .A(\ab[3][30] ), .B(\ab[2][31] ), .CI(\CARRYB[2][30] ), 
        .CO(\CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FADDX2 S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FADDX1 S2_20_5 ( .A(\SUMB[19][6] ), .B(\ab[20][5] ), .CI(\CARRYB[19][5] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FADDX1 S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FADDX2 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FADDX1 S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FADDX1 S2_22_28 ( .A(\CARRYB[21][28] ), .B(\ab[22][28] ), .CI(\SUMB[21][29] ), .CO(\CARRYB[22][28] ), .S(\SUMB[22][28] ) );
  FADDX1 S2_29_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FADDX1 S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FADDX1 S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FADDX2 S2_30_18 ( .A(\ab[30][18] ), .B(\CARRYB[29][18] ), .CI(\SUMB[29][19] ), .CO(\CARRYB[30][18] ), .S(\SUMB[30][18] ) );
  FADDX1 S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FADDX1 S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FADDX1 S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FADDX1 S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FADDX1 S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FADDX2 S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FADDX1 S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FADDX1 S2_2_20 ( .A(\ab[2][20] ), .B(n8), .CI(\SUMB[1][21] ), .CO(
        \CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FADDX1 S2_8_19 ( .A(\CARRYB[7][19] ), .B(\ab[8][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FADDX1 S2_6_21 ( .A(\CARRYB[5][21] ), .B(\ab[6][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FADDX1 S2_2_21 ( .A(\ab[2][21] ), .B(n1581), .CI(\SUMB[1][22] ), .CO(
        \CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FADDX1 S2_28_23 ( .A(\ab[28][23] ), .B(\CARRYB[27][23] ), .CI(\SUMB[27][24] ), .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FADDX2 S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FADDX1 S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FADDX1 S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FADDX1 S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FADDX1 S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FADDX1 S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FADDX1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FADDX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FADDX1 S2_9_4 ( .A(\ab[9][4] ), .B(\SUMB[8][5] ), .CI(\CARRYB[8][4] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FADDX1 S3_5_30 ( .A(\ab[5][30] ), .B(\ab[4][31] ), .CI(\CARRYB[4][30] ), 
        .CO(\CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FADDX1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FADDX1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FADDX1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FADDX1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FADDX1 S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FADDX1 S2_7_23 ( .A(\CARRYB[6][23] ), .B(\ab[7][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FADDX1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FADDX1 S2_13_21 ( .A(\ab[13][21] ), .B(\SUMB[12][22] ), .CI(\CARRYB[12][21] ), .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FADDX1 S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FADDX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FADDX1 S2_14_8 ( .A(\CARRYB[13][8] ), .B(\ab[14][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FADDX2 S2_7_20 ( .A(\CARRYB[6][20] ), .B(\ab[7][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FADDX1 S2_14_15 ( .A(\ab[14][15] ), .B(\SUMB[13][16] ), .CI(\CARRYB[13][15] ), .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FADDX1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FADDX2 S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FADDX1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FADDX1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FADDX1 S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(\A1[25] ) );
  FADDX1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FADDX1 S2_24_1 ( .A(\ab[24][1] ), .B(\SUMB[23][2] ), .CI(\CARRYB[23][1] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FADDX1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FADDX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FADDX1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FADDX1 S2_8_3 ( .A(\CARRYB[7][3] ), .B(\ab[8][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FADDX1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FADDX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FADDX1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FADDX1 S2_30_14 ( .A(\ab[30][14] ), .B(\CARRYB[29][14] ), .CI(\SUMB[29][15] ), .CO(\CARRYB[30][14] ), .S(\SUMB[30][14] ) );
  FADDX1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FADDX1 S2_27_29 ( .A(\ab[27][29] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FADDX1 S2_26_28 ( .A(\ab[26][28] ), .B(\CARRYB[25][28] ), .CI(\SUMB[25][29] ), .CO(\CARRYB[26][28] ), .S(\SUMB[26][28] ) );
  FADDX1 S2_26_26 ( .A(\ab[26][26] ), .B(\CARRYB[25][26] ), .CI(\SUMB[25][27] ), .CO(\CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FADDX1 S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FADDX1 S2_26_22 ( .A(\ab[26][22] ), .B(\CARRYB[25][22] ), .CI(\SUMB[25][23] ), .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FADDX1 S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FADDX1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FADDX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FADDX1 S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FADDX1 S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FADDX1 S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FADDX1 S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FADDX1 S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FADDX1 S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FADDX1 S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FADDX1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FADDX1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FADDX1 S2_2_28 ( .A(\ab[2][28] ), .B(n7), .CI(\SUMB[1][29] ), .CO(
        \CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  FADDX1 S3_2_30 ( .A(\ab[2][30] ), .B(\ab[1][31] ), .CI(n422), .CO(
        \CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  FADDX1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FADDX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FADDX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FADDX1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FADDX1 S2_6_2 ( .A(\SUMB[5][3] ), .B(\ab[6][2] ), .CI(\CARRYB[5][2] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FADDX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FADDX1 S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FADDX1 S2_25_28 ( .A(\ab[25][28] ), .B(\SUMB[24][29] ), .CI(\CARRYB[24][28] ), .CO(\CARRYB[25][28] ), .S(\SUMB[25][28] ) );
  FADDX1 S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FADDX1 S2_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FADDX1 S2_22_18 ( .A(\CARRYB[21][18] ), .B(\ab[22][18] ), .CI(\SUMB[21][19] ), .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FADDX1 S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FADDX1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FADDX1 S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FADDX1 S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FADDX1 S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FADDX1 S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FADDX1 S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FADDX1 S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FADDX1 S2_2_17 ( .A(\ab[2][17] ), .B(n5), .CI(\SUMB[1][18] ), .CO(
        \CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FADDX1 S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FADDX1 S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FADDX1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FADDX1 S2_2_29 ( .A(n687), .B(\ab[2][29] ), .CI(\SUMB[1][30] ), .CO(
        \CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FADDX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FADDX1 S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FADDX1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FADDX1 S2_29_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), 
        .CO(\CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FADDX1 S2_25_7 ( .A(\ab[25][7] ), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FADDX1 S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FADDX1 S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FADDX1 S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FADDX1 S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FADDX1 S2_7_27 ( .A(\ab[7][27] ), .B(\CARRYB[6][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FADDX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FADDX1 S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FADDX1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FADDX1 S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FADDX1 S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FADDX1 S2_14_21 ( .A(\SUMB[13][22] ), .B(\ab[14][21] ), .CI(\CARRYB[13][21] ), .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FADDX2 S2_28_11 ( .A(\ab[28][11] ), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), .CO(\CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FADDX2 S2_23_11 ( .A(\CARRYB[22][11] ), .B(\ab[23][11] ), .CI(\SUMB[22][12] ), .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FADDX2 S2_30_23 ( .A(\ab[30][23] ), .B(\CARRYB[29][23] ), .CI(\SUMB[29][24] ), .CO(\CARRYB[30][23] ), .S(\SUMB[30][23] ) );
  FADDX2 S2_30_1 ( .A(\ab[30][1] ), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), 
        .CO(\CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FADDX2 S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FADDX2 S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  AND2X4 U2 ( .IN1(\CARRYB[31][1] ), .IN2(\SUMB[31][2] ), .Q(n1977) );
  XOR2X2 U3 ( .IN1(n1456), .IN2(\CARRYB[2][25] ), .Q(\SUMB[3][25] ) );
  NAND3X4 U4 ( .IN1(n58), .IN2(n60), .IN3(n59), .QN(n22) );
  NAND3X1 U5 ( .IN1(n1304), .IN2(n1305), .IN3(n1306), .QN(\CARRYB[22][12] ) );
  NAND3X1 U6 ( .IN1(n1161), .IN2(n1163), .IN3(n1162), .QN(\CARRYB[15][22] ) );
  NAND3X1 U7 ( .IN1(n1896), .IN2(n1897), .IN3(n1898), .QN(\CARRYB[19][12] ) );
  NAND3X1 U8 ( .IN1(n774), .IN2(n775), .IN3(n776), .QN(\CARRYB[27][20] ) );
  NAND3X1 U9 ( .IN1(n934), .IN2(n935), .IN3(n936), .QN(\CARRYB[6][15] ) );
  NAND3X0 U10 ( .IN1(n233), .IN2(n234), .IN3(n235), .QN(\CARRYB[11][23] ) );
  NAND3X0 U11 ( .IN1(n562), .IN2(n561), .IN3(n563), .QN(\CARRYB[13][24] ) );
  NAND3X0 U12 ( .IN1(n253), .IN2(n254), .IN3(n255), .QN(\CARRYB[14][25] ) );
  XOR2X1 U13 ( .IN1(n1038), .IN2(\CARRYB[13][26] ), .Q(\SUMB[14][26] ) );
  NAND3X0 U14 ( .IN1(n1675), .IN2(n1676), .IN3(n1677), .QN(\CARRYB[13][11] )
         );
  NAND3X0 U15 ( .IN1(n1686), .IN2(n1687), .IN3(n1688), .QN(\CARRYB[19][14] )
         );
  NAND3X0 U16 ( .IN1(n1250), .IN2(n1249), .IN3(n1248), .QN(\CARRYB[22][15] )
         );
  XOR2X1 U17 ( .IN1(n1480), .IN2(\CARRYB[21][16] ), .Q(\SUMB[22][16] ) );
  XOR2X1 U18 ( .IN1(n269), .IN2(\CARRYB[14][10] ), .Q(\SUMB[15][10] ) );
  NAND3X0 U19 ( .IN1(n809), .IN2(n810), .IN3(n811), .QN(\CARRYB[27][9] ) );
  NAND3X0 U20 ( .IN1(n543), .IN2(n544), .IN3(n545), .QN(\CARRYB[4][5] ) );
  NAND3X0 U21 ( .IN1(n1813), .IN2(n1814), .IN3(n1815), .QN(\CARRYB[26][4] ) );
  XOR2X1 U22 ( .IN1(n542), .IN2(\CARRYB[3][5] ), .Q(\SUMB[4][5] ) );
  NAND3X0 U23 ( .IN1(n1201), .IN2(n1202), .IN3(n1203), .QN(\CARRYB[4][4] ) );
  NAND3X0 U24 ( .IN1(n1021), .IN2(n1022), .IN3(n1023), .QN(\CARRYB[5][26] ) );
  NAND3X0 U25 ( .IN1(n401), .IN2(n402), .IN3(n403), .QN(\CARRYB[2][27] ) );
  XOR2X1 U26 ( .IN1(n567), .IN2(\CARRYB[5][28] ), .Q(\SUMB[6][28] ) );
  NAND3X0 U27 ( .IN1(n915), .IN2(n916), .IN3(n917), .QN(\CARRYB[6][27] ) );
  NAND3X0 U28 ( .IN1(n209), .IN2(n210), .IN3(n211), .QN(\CARRYB[7][26] ) );
  NAND3X0 U29 ( .IN1(n1411), .IN2(n1412), .IN3(n1413), .QN(\CARRYB[10][27] )
         );
  NAND3X0 U30 ( .IN1(n1599), .IN2(n1600), .IN3(n1601), .QN(\CARRYB[4][19] ) );
  NAND3X0 U31 ( .IN1(n1496), .IN2(n1495), .IN3(n1497), .QN(\CARRYB[9][24] ) );
  XOR2X1 U32 ( .IN1(n1449), .IN2(\CARRYB[8][25] ), .Q(\SUMB[9][25] ) );
  XOR2X1 U33 ( .IN1(n1009), .IN2(\CARRYB[12][23] ), .Q(\SUMB[13][23] ) );
  NAND3X0 U34 ( .IN1(n989), .IN2(n990), .IN3(n991), .QN(\CARRYB[3][16] ) );
  XOR2X1 U35 ( .IN1(n232), .IN2(\SUMB[11][23] ), .Q(\SUMB[12][22] ) );
  XOR2X1 U36 ( .IN1(n252), .IN2(\CARRYB[13][25] ), .Q(\SUMB[14][25] ) );
  NAND3X0 U37 ( .IN1(n1738), .IN2(n1739), .IN3(n1740), .QN(\CARRYB[8][13] ) );
  NAND3X0 U38 ( .IN1(n652), .IN2(n653), .IN3(n654), .QN(\CARRYB[18][25] ) );
  XOR2X1 U39 ( .IN1(n901), .IN2(\CARRYB[16][24] ), .Q(\SUMB[17][24] ) );
  NAND3X0 U40 ( .IN1(n1185), .IN2(n1186), .IN3(n1187), .QN(\CARRYB[17][21] )
         );
  NAND3X0 U41 ( .IN1(n306), .IN2(n307), .IN3(n308), .QN(\CARRYB[20][16] ) );
  NAND3X0 U42 ( .IN1(n1651), .IN2(n1652), .IN3(n1653), .QN(\CARRYB[11][11] )
         );
  XOR2X1 U43 ( .IN1(n496), .IN2(\CARRYB[10][13] ), .Q(\SUMB[11][13] ) );
  NAND3X0 U44 ( .IN1(n1321), .IN2(n1322), .IN3(n1323), .QN(\CARRYB[11][12] )
         );
  NAND3X0 U45 ( .IN1(n1014), .IN2(n1015), .IN3(n1016), .QN(\CARRYB[21][19] )
         );
  NAND3X0 U46 ( .IN1(n1265), .IN2(n1266), .IN3(n1267), .QN(\CARRYB[21][29] )
         );
  NAND3X0 U47 ( .IN1(n1617), .IN2(n1618), .IN3(n1619), .QN(\CARRYB[14][12] )
         );
  NAND3X0 U48 ( .IN1(n1092), .IN2(n1093), .IN3(n1094), .QN(\CARRYB[22][14] )
         );
  XNOR2X1 U49 ( .IN1(n623), .IN2(\CARRYB[20][21] ), .Q(\SUMB[21][21] ) );
  NAND3X0 U50 ( .IN1(n571), .IN2(n572), .IN3(n573), .QN(\CARRYB[21][20] ) );
  NAND3X0 U51 ( .IN1(n892), .IN2(n893), .IN3(n894), .QN(\CARRYB[23][24] ) );
  NAND3X0 U52 ( .IN1(n1467), .IN2(n1468), .IN3(n1469), .QN(\CARRYB[24][25] )
         );
  NAND3X0 U53 ( .IN1(n588), .IN2(n589), .IN3(n590), .QN(\CARRYB[17][8] ) );
  NAND3X0 U54 ( .IN1(n606), .IN2(n607), .IN3(n608), .QN(\CARRYB[24][16] ) );
  NAND3X0 U55 ( .IN1(n1103), .IN2(n1104), .IN3(n1105), .QN(\CARRYB[25][14] )
         );
  XOR2X1 U56 ( .IN1(n1258), .IN2(\SUMB[23][29] ), .Q(\SUMB[24][28] ) );
  NAND3X0 U57 ( .IN1(n1295), .IN2(n1296), .IN3(n1297), .QN(\CARRYB[19][8] ) );
  NAND3X0 U58 ( .IN1(n1151), .IN2(n1152), .IN3(n1153), .QN(\CARRYB[27][19] )
         );
  NAND3X0 U59 ( .IN1(n692), .IN2(n693), .IN3(n694), .QN(\CARRYB[26][21] ) );
  NAND3X0 U60 ( .IN1(n1694), .IN2(n1695), .IN3(n1696), .QN(\CARRYB[28][6] ) );
  NAND3X0 U61 ( .IN1(n135), .IN2(n136), .IN3(n137), .QN(\CARRYB[27][23] ) );
  NAND3X0 U62 ( .IN1(n1197), .IN2(n1198), .IN3(n1199), .QN(\CARRYB[3][4] ) );
  NAND3X0 U63 ( .IN1(n103), .IN2(n104), .IN3(n105), .QN(\CARRYB[6][5] ) );
  NAND3X0 U64 ( .IN1(n733), .IN2(n734), .IN3(n735), .QN(\CARRYB[12][3] ) );
  NAND3X0 U65 ( .IN1(n1794), .IN2(n1795), .IN3(n1796), .QN(\CARRYB[15][3] ) );
  NAND3X0 U66 ( .IN1(n625), .IN2(n626), .IN3(n627), .QN(\CARRYB[20][3] ) );
  XOR2X1 U67 ( .IN1(n584), .IN2(\CARRYB[21][6] ), .Q(\SUMB[22][6] ) );
  XOR2X1 U68 ( .IN1(n290), .IN2(\CARRYB[26][5] ), .Q(\SUMB[27][5] ) );
  NAND3X0 U69 ( .IN1(n508), .IN2(n509), .IN3(n510), .QN(\CARRYB[29][7] ) );
  NAND3X0 U70 ( .IN1(n1728), .IN2(n1729), .IN3(n1730), .QN(\CARRYB[28][13] )
         );
  XOR2X1 U71 ( .IN1(n1116), .IN2(\SUMB[27][27] ), .Q(\SUMB[28][26] ) );
  NAND3X0 U72 ( .IN1(n862), .IN2(n863), .IN3(n864), .QN(\CARRYB[6][3] ) );
  NAND3X0 U73 ( .IN1(n331), .IN2(n332), .IN3(n333), .QN(\CARRYB[21][2] ) );
  NAND3X0 U74 ( .IN1(n1337), .IN2(n1338), .IN3(n1339), .QN(\CARRYB[24][3] ) );
  AND2X1 U75 ( .IN1(\ab[0][30] ), .IN2(\ab[1][29] ), .Q(n687) );
  XOR2X1 U76 ( .IN1(n141), .IN2(\SUMB[4][30] ), .Q(\SUMB[5][29] ) );
  NAND3X0 U77 ( .IN1(n564), .IN2(n565), .IN3(n566), .QN(\CARRYB[5][28] ) );
  XOR2X1 U78 ( .IN1(n411), .IN2(\CARRYB[4][27] ), .Q(\SUMB[5][27] ) );
  XOR2X1 U79 ( .IN1(n404), .IN2(\CARRYB[2][27] ), .Q(\SUMB[3][27] ) );
  NAND3X0 U80 ( .IN1(n1024), .IN2(n1025), .IN3(n1026), .QN(\CARRYB[3][26] ) );
  NAND3X0 U81 ( .IN1(n1457), .IN2(n1458), .IN3(n1459), .QN(\CARRYB[3][25] ) );
  NAND3X0 U82 ( .IN1(n178), .IN2(n179), .IN3(n180), .QN(\CARRYB[3][23] ) );
  NAND3X0 U83 ( .IN1(n780), .IN2(n782), .IN3(n781), .QN(\CARRYB[8][26] ) );
  NAND3X0 U84 ( .IN1(n115), .IN2(n116), .IN3(n117), .QN(\CARRYB[7][25] ) );
  XOR2X1 U85 ( .IN1(n208), .IN2(\CARRYB[6][26] ), .Q(\SUMB[7][26] ) );
  XOR2X1 U86 ( .IN1(\ab[9][29] ), .IN2(\SUMB[8][30] ), .Q(n338) );
  XOR2X1 U87 ( .IN1(\ab[1][21] ), .IN2(\ab[0][22] ), .Q(\SUMB[1][21] ) );
  NAND3X0 U88 ( .IN1(n159), .IN2(n160), .IN3(n161), .QN(\CARRYB[8][21] ) );
  NAND3X0 U89 ( .IN1(n912), .IN2(n913), .IN3(n914), .QN(\CARRYB[10][26] ) );
  NAND3X0 U90 ( .IN1(n771), .IN2(n772), .IN3(n773), .QN(\CARRYB[10][25] ) );
  XOR2X1 U91 ( .IN1(n970), .IN2(n349), .Q(\SUMB[11][29] ) );
  NAND3X0 U92 ( .IN1(n1603), .IN2(n1604), .IN3(n1605), .QN(\CARRYB[5][19] ) );
  NAND3X0 U93 ( .IN1(n614), .IN2(n615), .IN3(n616), .QN(\CARRYB[9][23] ) );
  NAND3X0 U94 ( .IN1(n1006), .IN2(n1007), .IN3(n1008), .QN(\CARRYB[12][23] )
         );
  XOR2X1 U95 ( .IN1(n908), .IN2(\CARRYB[11][26] ), .Q(\SUMB[12][26] ) );
  NAND3X0 U96 ( .IN1(n1415), .IN2(n1416), .IN3(n1417), .QN(\CARRYB[11][27] )
         );
  NAND3X0 U97 ( .IN1(n909), .IN2(n910), .IN3(n911), .QN(\CARRYB[12][26] ) );
  NAND3X0 U98 ( .IN1(n844), .IN2(n845), .IN3(n846), .QN(\CARRYB[13][30] ) );
  XOR2X1 U99 ( .IN1(n818), .IN2(\CARRYB[3][17] ), .Q(\SUMB[4][17] ) );
  NAND3X0 U100 ( .IN1(n993), .IN2(n994), .IN3(n995), .QN(\CARRYB[4][16] ) );
  NAND3X0 U101 ( .IN1(n819), .IN2(n820), .IN3(n821), .QN(\CARRYB[4][17] ) );
  XOR2X1 U102 ( .IN1(n1633), .IN2(\CARRYB[3][18] ), .Q(\SUMB[4][18] ) );
  XOR2X1 U103 ( .IN1(n613), .IN2(\SUMB[9][23] ), .Q(\SUMB[10][22] ) );
  NAND3X0 U104 ( .IN1(n314), .IN2(n313), .IN3(n315), .QN(\CARRYB[10][21] ) );
  NAND3X0 U105 ( .IN1(n515), .IN2(n516), .IN3(n517), .QN(\CARRYB[15][20] ) );
  XOR3X1 U106 ( .IN1(\ab[15][21] ), .IN2(\CARRYB[14][21] ), .IN3(
        \SUMB[14][22] ), .Q(\SUMB[15][21] ) );
  NAND3X0 U107 ( .IN1(n198), .IN2(n199), .IN3(n200), .QN(\CARRYB[14][23] ) );
  XOR2X1 U108 ( .IN1(n1240), .IN2(\CARRYB[7][17] ), .Q(\SUMB[8][17] ) );
  NAND3X0 U109 ( .IN1(n30), .IN2(n31), .IN3(n32), .QN(\CARRYB[8][16] ) );
  NAND3X0 U110 ( .IN1(n799), .IN2(n800), .IN3(n801), .QN(\CARRYB[11][18] ) );
  NAND3X0 U111 ( .IN1(n1039), .IN2(n1040), .IN3(n1041), .QN(\CARRYB[14][26] )
         );
  NAND3X0 U112 ( .IN1(n710), .IN2(n711), .IN3(n712), .QN(\CARRYB[15][21] ) );
  NAND3X0 U113 ( .IN1(n937), .IN2(n938), .IN3(n939), .QN(\CARRYB[7][14] ) );
  XOR2X1 U114 ( .IN1(n985), .IN2(\CARRYB[5][16] ), .Q(\SUMB[6][16] ) );
  XOR3X1 U115 ( .IN1(\ab[13][19] ), .IN2(\CARRYB[12][19] ), .IN3(
        \SUMB[12][20] ), .Q(\SUMB[13][19] ) );
  XOR3X1 U116 ( .IN1(\ab[17][20] ), .IN2(\SUMB[16][21] ), .IN3(
        \CARRYB[16][20] ), .Q(\SUMB[17][20] ) );
  NAND3X0 U117 ( .IN1(n519), .IN2(n520), .IN3(n521), .QN(\CARRYB[17][18] ) );
  XOR2X1 U118 ( .IN1(n1404), .IN2(\CARRYB[16][27] ), .Q(\SUMB[17][27] ) );
  NAND3X0 U119 ( .IN1(n1405), .IN2(n1406), .IN3(n1407), .QN(\CARRYB[17][27] )
         );
  NAND3X0 U120 ( .IN1(n1574), .IN2(n1575), .IN3(n1576), .QN(\CARRYB[16][30] )
         );
  NAND3X0 U121 ( .IN1(n1624), .IN2(n1625), .IN3(n1626), .QN(\CARRYB[5][13] )
         );
  XOR3X1 U122 ( .IN1(\ab[10][17] ), .IN2(\CARRYB[9][17] ), .IN3(\SUMB[9][18] ), 
        .Q(\SUMB[10][17] ) );
  NAND3X0 U123 ( .IN1(n826), .IN2(n827), .IN3(n828), .QN(\CARRYB[10][16] ) );
  NAND3X0 U124 ( .IN1(n964), .IN2(n965), .IN3(n966), .QN(\CARRYB[16][14] ) );
  XOR2X1 U125 ( .IN1(n832), .IN2(\CARRYB[15][15] ), .Q(\SUMB[16][15] ) );
  NAND3X0 U126 ( .IN1(n902), .IN2(n903), .IN3(n904), .QN(\CARRYB[17][24] ) );
  NAND3X0 U127 ( .IN1(n246), .IN2(n247), .IN3(n248), .QN(\CARRYB[18][24] ) );
  NAND3X0 U128 ( .IN1(n1032), .IN2(n1033), .IN3(n1034), .QN(\CARRYB[19][25] )
         );
  NAND3X0 U129 ( .IN1(n1327), .IN2(n1328), .IN3(n1329), .QN(\CARRYB[10][12] )
         );
  XOR3X1 U130 ( .IN1(\ab[9][13] ), .IN2(\CARRYB[8][13] ), .IN3(\SUMB[8][14] ), 
        .Q(\SUMB[9][13] ) );
  XOR3X1 U131 ( .IN1(\SUMB[15][15] ), .IN2(\ab[16][14] ), .IN3(
        \CARRYB[15][14] ), .Q(\SUMB[16][14] ) );
  NAND3X0 U132 ( .IN1(n451), .IN2(n452), .IN3(n453), .QN(\CARRYB[16][17] ) );
  NAND3X0 U133 ( .IN1(n1251), .IN2(n1252), .IN3(n1253), .QN(\CARRYB[20][15] )
         );
  XOR2X1 U134 ( .IN1(n353), .IN2(\CARRYB[2][14] ), .Q(\SUMB[3][14] ) );
  XOR2X1 U135 ( .IN1(n1623), .IN2(\CARRYB[4][13] ), .Q(\SUMB[5][13] ) );
  XOR3X1 U136 ( .IN1(\CARRYB[10][11] ), .IN2(\ab[11][11] ), .IN3(
        \SUMB[10][12] ), .Q(n591) );
  NAND3X0 U137 ( .IN1(n695), .IN2(n696), .IN3(n697), .QN(\CARRYB[11][10] ) );
  XOR2X1 U138 ( .IN1(n1616), .IN2(\CARRYB[13][12] ), .Q(\SUMB[14][12] ) );
  NAND3X0 U139 ( .IN1(n1679), .IN2(n1680), .IN3(n1681), .QN(\CARRYB[14][11] )
         );
  NAND3X0 U140 ( .IN1(n1721), .IN2(n1722), .IN3(n1723), .QN(\CARRYB[13][13] )
         );
  XOR2X1 U141 ( .IN1(n464), .IN2(\CARRYB[18][13] ), .Q(\SUMB[19][13] ) );
  NAND3X0 U142 ( .IN1(n1641), .IN2(n1642), .IN3(n1643), .QN(\CARRYB[21][18] )
         );
  XOR2X1 U143 ( .IN1(n1013), .IN2(\SUMB[20][20] ), .Q(\SUMB[21][19] ) );
  XOR2X1 U144 ( .IN1(n1664), .IN2(\CARRYB[20][17] ), .Q(\SUMB[21][17] ) );
  NAND3X0 U145 ( .IN1(n1477), .IN2(n1478), .IN3(n1479), .QN(\CARRYB[21][16] )
         );
  NAND3X0 U146 ( .IN1(n1086), .IN2(n1087), .IN3(n1088), .QN(\CARRYB[20][21] )
         );
  NAND3X0 U147 ( .IN1(n777), .IN2(n778), .IN3(n779), .QN(\CARRYB[22][23] ) );
  XOR2X1 U148 ( .IN1(\SUMB[1][13] ), .IN2(n9), .Q(n1899) );
  AND2X1 U149 ( .IN1(\ab[0][12] ), .IN2(\ab[1][11] ), .Q(n1689) );
  NAND3X0 U150 ( .IN1(n1648), .IN2(n1649), .IN3(n1650), .QN(\CARRYB[13][10] )
         );
  NAND3X0 U151 ( .IN1(n270), .IN2(n271), .IN3(n272), .QN(\CARRYB[15][10] ) );
  NAND3X0 U152 ( .IN1(n1269), .IN2(n1270), .IN3(n1271), .QN(\CARRYB[22][29] )
         );
  NAND3X0 U153 ( .IN1(n723), .IN2(n724), .IN3(n725), .QN(\CARRYB[5][10] ) );
  NAND3X0 U154 ( .IN1(n1560), .IN2(n1561), .IN3(n1562), .QN(\CARRYB[16][11] )
         );
  XOR2X1 U155 ( .IN1(n276), .IN2(\CARRYB[16][10] ), .Q(\SUMB[17][10] ) );
  NAND3X0 U156 ( .IN1(n1289), .IN2(n1290), .IN3(n1291), .QN(\CARRYB[17][9] )
         );
  NAND3X0 U157 ( .IN1(n1070), .IN2(n1071), .IN3(n1072), .QN(\CARRYB[22][9] )
         );
  NAND3X0 U158 ( .IN1(n1279), .IN2(n1280), .IN3(n1281), .QN(\CARRYB[23][13] )
         );
  XOR2X1 U159 ( .IN1(n1095), .IN2(\CARRYB[22][14] ), .Q(\SUMB[23][14] ) );
  XOR2X1 U160 ( .IN1(n605), .IN2(\CARRYB[23][16] ), .Q(\SUMB[24][16] ) );
  NAND3X0 U161 ( .IN1(n1099), .IN2(n1100), .IN3(n1101), .QN(\CARRYB[24][14] )
         );
  XOR2X1 U162 ( .IN1(n430), .IN2(\SUMB[22][21] ), .Q(\SUMB[23][20] ) );
  XNOR3X1 U163 ( .IN1(\CARRYB[23][24] ), .IN2(n659), .IN3(\SUMB[23][25] ), .Q(
        \SUMB[24][24] ) );
  NAND3X0 U164 ( .IN1(n1515), .IN2(n1516), .IN3(n1517), .QN(\CARRYB[24][23] )
         );
  XOR2X1 U165 ( .IN1(\ab[1][8] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][8] ) );
  NAND3X0 U166 ( .IN1(n639), .IN2(n640), .IN3(n641), .QN(\CARRYB[8][8] ) );
  NAND3X0 U167 ( .IN1(n1764), .IN2(n1765), .IN3(n1766), .QN(\CARRYB[19][9] )
         );
  NAND3X0 U168 ( .IN1(n1749), .IN2(n1750), .IN3(n1751), .QN(\CARRYB[20][7] )
         );
  NAND3X0 U169 ( .IN1(n1505), .IN2(n1506), .IN3(n1507), .QN(\CARRYB[25][24] )
         );
  NAND3X0 U170 ( .IN1(n1364), .IN2(n1365), .IN3(n1366), .QN(\CARRYB[24][29] )
         );
  NAND3X0 U171 ( .IN1(n1262), .IN2(n1263), .IN3(n1264), .QN(\CARRYB[24][28] )
         );
  NAND3X0 U172 ( .IN1(n1460), .IN2(n1461), .IN3(n1462), .QN(\CARRYB[25][25] )
         );
  NAND3X0 U173 ( .IN1(n1368), .IN2(n1369), .IN3(n1370), .QN(\CARRYB[25][29] )
         );
  NAND3X0 U174 ( .IN1(n1219), .IN2(n1220), .IN3(n1221), .QN(\CARRYB[2][8] ) );
  XOR2X1 U175 ( .IN1(n360), .IN2(\CARRYB[15][6] ), .Q(\SUMB[16][6] ) );
  XNOR2X1 U176 ( .IN1(n702), .IN2(\SUMB[17][9] ), .Q(\SUMB[18][8] ) );
  NAND3X0 U177 ( .IN1(n1213), .IN2(n1214), .IN3(n1215), .QN(\CARRYB[18][7] )
         );
  NAND3X0 U178 ( .IN1(n1286), .IN2(n1287), .IN3(n1288), .QN(\CARRYB[22][7] )
         );
  NAND3X0 U179 ( .IN1(n1905), .IN2(n1906), .IN3(n1907), .QN(\CARRYB[28][5] )
         );
  XOR3X1 U180 ( .IN1(\ab[26][10] ), .IN2(\CARRYB[25][10] ), .IN3(
        \SUMB[25][11] ), .Q(\SUMB[26][10] ) );
  NAND3X0 U181 ( .IN1(n511), .IN2(n512), .IN3(n513), .QN(\CARRYB[27][7] ) );
  NAND3X0 U182 ( .IN1(n1528), .IN2(n1529), .IN3(n1530), .QN(\CARRYB[26][15] )
         );
  NAND3X0 U183 ( .IN1(n1474), .IN2(n1475), .IN3(n1476), .QN(\CARRYB[26][14] )
         );
  NBUFFX2 U184 ( .INP(n2219), .Z(n2122) );
  NAND3X0 U185 ( .IN1(n1117), .IN2(n1118), .IN3(n1119), .QN(\CARRYB[27][27] )
         );
  NAND3X0 U186 ( .IN1(n1826), .IN2(n1827), .IN3(n1828), .QN(\CARRYB[11][4] )
         );
  NAND3X0 U187 ( .IN1(n1216), .IN2(n1217), .IN3(n1218), .QN(\CARRYB[19][6] )
         );
  XOR3X1 U188 ( .IN1(\ab[19][7] ), .IN2(\CARRYB[18][7] ), .IN3(\SUMB[18][8] ), 
        .Q(\SUMB[19][7] ) );
  NAND3X0 U189 ( .IN1(n872), .IN2(n873), .IN3(n874), .QN(\CARRYB[28][17] ) );
  NAND3X0 U190 ( .IN1(n256), .IN2(n257), .IN3(n258), .QN(\CARRYB[29][22] ) );
  NAND3X0 U191 ( .IN1(n750), .IN2(n751), .IN3(n752), .QN(\CARRYB[14][5] ) );
  NAND3X0 U192 ( .IN1(n1801), .IN2(n1802), .IN3(n1803), .QN(\CARRYB[17][3] )
         );
  NAND3X0 U193 ( .IN1(n1916), .IN2(n1917), .IN3(n1918), .QN(\CARRYB[19][5] )
         );
  XOR2X1 U194 ( .IN1(n1282), .IN2(\SUMB[21][8] ), .Q(\SUMB[22][7] ) );
  NAND3X0 U195 ( .IN1(n585), .IN2(n586), .IN3(n587), .QN(\CARRYB[22][6] ) );
  NAND3X0 U196 ( .IN1(n1809), .IN2(n1810), .IN3(n1811), .QN(\CARRYB[25][4] )
         );
  NAND3X0 U197 ( .IN1(n1787), .IN2(n1788), .IN3(n1789), .QN(\CARRYB[29][3] )
         );
  NAND3X0 U198 ( .IN1(n280), .IN2(n281), .IN3(n282), .QN(\CARRYB[30][4] ) );
  NAND3X0 U199 ( .IN1(n1909), .IN2(n1910), .IN3(n1911), .QN(\CARRYB[29][5] )
         );
  NAND3X0 U200 ( .IN1(n1746), .IN2(n1747), .IN3(n1748), .QN(\CARRYB[30][7] )
         );
  NAND3X0 U201 ( .IN1(n1836), .IN2(n1837), .IN3(n1838), .QN(\CARRYB[30][8] )
         );
  XOR2X1 U202 ( .IN1(n298), .IN2(\CARRYB[28][14] ), .Q(\SUMB[29][14] ) );
  NAND3X0 U203 ( .IN1(n865), .IN2(n866), .IN3(n867), .QN(\CARRYB[29][16] ) );
  NAND3X0 U204 ( .IN1(n787), .IN2(n788), .IN3(n789), .QN(\CARRYB[29][15] ) );
  XOR2X1 U205 ( .IN1(n999), .IN2(\CARRYB[28][18] ), .Q(\SUMB[29][18] ) );
  NAND3X0 U206 ( .IN1(n1000), .IN2(n1001), .IN3(n1002), .QN(\CARRYB[29][18] )
         );
  NAND3X0 U207 ( .IN1(n895), .IN2(n896), .IN3(n897), .QN(\CARRYB[29][21] ) );
  NAND3X0 U208 ( .IN1(n1484), .IN2(n1485), .IN3(n1486), .QN(\CARRYB[30][24] )
         );
  NAND3X0 U209 ( .IN1(n1439), .IN2(n1440), .IN3(n1441), .QN(\CARRYB[30][25] )
         );
  XOR2X1 U210 ( .IN1(n1421), .IN2(\CARRYB[28][27] ), .Q(\SUMB[29][27] ) );
  NAND3X0 U211 ( .IN1(n858), .IN2(n859), .IN3(n860), .QN(\CARRYB[5][3] ) );
  XOR2X1 U212 ( .IN1(n1797), .IN2(\CARRYB[15][3] ), .Q(\SUMB[16][3] ) );
  NAND3X0 U213 ( .IN1(n1204), .IN2(n1205), .IN3(n1206), .QN(\CARRYB[19][2] )
         );
  XOR2X1 U214 ( .IN1(n1786), .IN2(\CARRYB[28][3] ), .Q(\SUMB[29][3] ) );
  AND2X1 U215 ( .IN1(\ab[1][3] ), .IN2(\ab[0][4] ), .Q(n1808) );
  NAND3X0 U216 ( .IN1(n660), .IN2(n661), .IN3(n662), .QN(\CARRYB[2][2] ) );
  NAND3X0 U217 ( .IN1(n737), .IN2(n738), .IN3(n739), .QN(\CARRYB[13][3] ) );
  XNOR2X1 U218 ( .IN1(n381), .IN2(\CARRYB[20][4] ), .Q(\SUMB[21][4] ) );
  NAND3X0 U219 ( .IN1(n629), .IN2(n630), .IN3(n631), .QN(\CARRYB[21][3] ) );
  NAND3X0 U220 ( .IN1(n1132), .IN2(n1133), .IN3(n1134), .QN(\CARRYB[22][2] )
         );
  NAND3X0 U221 ( .IN1(n128), .IN2(n129), .IN3(n130), .QN(\CARRYB[9][1] ) );
  XOR2X1 U222 ( .IN1(n1435), .IN2(n19), .Q(\SUMB[18][1] ) );
  NAND3X0 U223 ( .IN1(n918), .IN2(n919), .IN3(n920), .QN(\CARRYB[18][0] ) );
  XOR2X1 U224 ( .IN1(n1932), .IN2(\CARRYB[24][2] ), .Q(\SUMB[25][2] ) );
  NAND3X0 U225 ( .IN1(n1933), .IN2(n1934), .IN3(n1935), .QN(\CARRYB[25][2] )
         );
  XOR2X1 U226 ( .IN1(n925), .IN2(\SUMB[12][2] ), .Q(\SUMB[13][1] ) );
  AND2X1 U227 ( .IN1(n2206), .IN2(n148), .Q(\ab[1][31] ) );
  NAND3X0 U228 ( .IN1(n216), .IN2(n217), .IN3(n218), .QN(\CARRYB[4][28] ) );
  XOR2X1 U229 ( .IN1(\ab[4][28] ), .IN2(\SUMB[3][29] ), .Q(n215) );
  XOR2X1 U230 ( .IN1(n1020), .IN2(\CARRYB[4][26] ), .Q(\SUMB[5][26] ) );
  XOR2X1 U231 ( .IN1(\ab[1][29] ), .IN2(\ab[0][30] ), .Q(\SUMB[1][29] ) );
  AND2X1 U232 ( .IN1(\ab[1][26] ), .IN2(\ab[0][27] ), .Q(n165) );
  AND2X1 U233 ( .IN1(\ab[0][24] ), .IN2(\ab[1][23] ), .Q(n1123) );
  NAND3X0 U234 ( .IN1(n568), .IN2(n569), .IN3(n570), .QN(\CARRYB[6][28] ) );
  NAND3X0 U235 ( .IN1(n205), .IN2(n206), .IN3(n207), .QN(\CARRYB[6][26] ) );
  XOR2X1 U236 ( .IN1(\ab[8][30] ), .IN2(\ab[7][31] ), .Q(n854) );
  NAND3X0 U237 ( .IN1(n1502), .IN2(n1503), .IN3(n1504), .QN(\CARRYB[3][24] )
         );
  NAND3X0 U238 ( .IN1(n182), .IN2(n183), .IN3(n184), .QN(\CARRYB[4][23] ) );
  XOR2X1 U239 ( .IN1(n99), .IN2(\CARRYB[6][24] ), .Q(\SUMB[7][24] ) );
  XOR2X1 U240 ( .IN1(\ab[7][25] ), .IN2(\SUMB[6][26] ), .Q(n114) );
  NAND3X0 U241 ( .IN1(n100), .IN2(n101), .IN3(n102), .QN(\CARRYB[7][24] ) );
  NAND3X0 U242 ( .IN1(n1408), .IN2(n1409), .IN3(n1410), .QN(\CARRYB[9][27] )
         );
  NAND3X0 U243 ( .IN1(n768), .IN2(n769), .IN3(n770), .QN(\CARRYB[9][26] ) );
  NAND3X0 U244 ( .IN1(n1542), .IN2(n1543), .IN3(n1544), .QN(\CARRYB[5][22] )
         );
  XOR2X1 U245 ( .IN1(n1602), .IN2(\CARRYB[4][19] ), .Q(\SUMB[5][19] ) );
  NAND3X0 U246 ( .IN1(n1446), .IN2(n1447), .IN3(n1448), .QN(\CARRYB[8][25] )
         );
  NAND3X0 U247 ( .IN1(n656), .IN2(n657), .IN3(n658), .QN(\CARRYB[10][28] ) );
  NAND3X0 U248 ( .IN1(n905), .IN2(n906), .IN3(n907), .QN(\CARRYB[11][26] ) );
  XOR2X1 U249 ( .IN1(n1414), .IN2(\CARRYB[10][27] ), .Q(\SUMB[11][27] ) );
  XOR2X1 U250 ( .IN1(\ab[1][19] ), .IN2(\ab[0][20] ), .Q(\SUMB[1][19] ) );
  NAND3X0 U251 ( .IN1(n1003), .IN2(n1004), .IN3(n1005), .QN(\CARRYB[10][23] )
         );
  XOR3X1 U252 ( .IN1(\ab[8][22] ), .IN2(\CARRYB[7][22] ), .IN3(\SUMB[7][23] ), 
        .Q(n27) );
  NAND3X0 U253 ( .IN1(n1385), .IN2(n1386), .IN3(n1387), .QN(\CARRYB[12][28] )
         );
  XOR2X1 U254 ( .IN1(n1384), .IN2(\CARRYB[11][28] ), .Q(\SUMB[12][28] ) );
  XOR2X1 U255 ( .IN1(n560), .IN2(\CARRYB[12][24] ), .Q(\SUMB[13][24] ) );
  NAND3X0 U256 ( .IN1(n1010), .IN2(n1011), .IN3(n1012), .QN(\CARRYB[13][23] )
         );
  NAND3X0 U257 ( .IN1(n1634), .IN2(n1635), .IN3(n1636), .QN(\CARRYB[4][18] )
         );
  XOR3X1 U258 ( .IN1(\ab[7][21] ), .IN2(\CARRYB[6][21] ), .IN3(\SUMB[6][22] ), 
        .Q(\SUMB[7][21] ) );
  XOR2X1 U259 ( .IN1(n959), .IN2(\CARRYB[6][18] ), .Q(\SUMB[7][18] ) );
  NAND3X0 U260 ( .IN1(n50), .IN2(n51), .IN3(n52), .QN(\CARRYB[7][16] ) );
  NOR2X0 U261 ( .IN1(n2134), .IN2(n2071), .QN(\ab[8][16] ) );
  NAND3X0 U262 ( .IN1(n236), .IN2(n237), .IN3(n238), .QN(\CARRYB[12][22] ) );
  NAND3X0 U263 ( .IN1(n617), .IN2(n618), .IN3(n619), .QN(\CARRYB[10][22] ) );
  XOR3X1 U264 ( .IN1(\ab[11][23] ), .IN2(\CARRYB[10][23] ), .IN3(
        \SUMB[10][24] ), .Q(\SUMB[11][23] ) );
  NAND3X0 U265 ( .IN1(n249), .IN2(n250), .IN3(n251), .QN(\CARRYB[13][25] ) );
  NAND3X0 U266 ( .IN1(n1035), .IN2(n1036), .IN3(n1037), .QN(\CARRYB[13][26] )
         );
  NAND3X0 U267 ( .IN1(n982), .IN2(n983), .IN3(n984), .QN(\CARRYB[5][16] ) );
  NAND3X0 U268 ( .IN1(n960), .IN2(n961), .IN3(n962), .QN(\CARRYB[7][18] ) );
  XOR2X1 U269 ( .IN1(n172), .IN2(\CARRYB[6][19] ), .Q(\SUMB[7][19] ) );
  NAND3X0 U270 ( .IN1(n444), .IN2(n445), .IN3(n446), .QN(\CARRYB[14][18] ) );
  XOR3X1 U271 ( .IN1(\CARRYB[15][21] ), .IN2(\ab[16][21] ), .IN3(
        \SUMB[15][22] ), .Q(\SUMB[16][21] ) );
  NAND3X0 U272 ( .IN1(n713), .IN2(n714), .IN3(n715), .QN(\CARRYB[16][20] ) );
  XNOR2X1 U273 ( .IN1(n624), .IN2(\SUMB[15][21] ), .Q(\SUMB[16][20] ) );
  NAND3X0 U274 ( .IN1(n1610), .IN2(n1611), .IN3(n1612), .QN(\CARRYB[16][19] )
         );
  XOR2X1 U275 ( .IN1(n201), .IN2(\CARRYB[14][23] ), .Q(\SUMB[15][23] ) );
  NAND3X0 U276 ( .IN1(n202), .IN2(n203), .IN3(n204), .QN(\CARRYB[15][23] ) );
  NAND3X0 U277 ( .IN1(n703), .IN2(n704), .IN3(n705), .QN(\CARRYB[17][20] ) );
  NAND3X0 U278 ( .IN1(n848), .IN2(n849), .IN3(n850), .QN(\CARRYB[14][30] ) );
  XOR2X1 U279 ( .IN1(n992), .IN2(\CARRYB[3][16] ), .Q(\SUMB[4][16] ) );
  XOR2X1 U280 ( .IN1(\ab[1][17] ), .IN2(\ab[0][18] ), .Q(\SUMB[1][17] ) );
  AND2X1 U281 ( .IN1(\ab[0][17] ), .IN2(\ab[1][16] ), .Q(n294) );
  NAND3X0 U282 ( .IN1(n1168), .IN2(n1169), .IN3(n1170), .QN(\CARRYB[8][14] )
         );
  XOR3X1 U283 ( .IN1(\ab[10][15] ), .IN2(\CARRYB[9][15] ), .IN3(\SUMB[9][16] ), 
        .Q(\SUMB[10][15] ) );
  NAND3X0 U284 ( .IN1(n822), .IN2(n823), .IN3(n824), .QN(\CARRYB[9][16] ) );
  NAND3X0 U285 ( .IN1(n1525), .IN2(n1526), .IN3(n1527), .QN(\CARRYB[13][16] )
         );
  NAND3X0 U286 ( .IN1(n441), .IN2(n442), .IN3(n443), .QN(\CARRYB[13][19] ) );
  XNOR2X1 U287 ( .IN1(n316), .IN2(\CARRYB[12][20] ), .Q(\SUMB[13][20] ) );
  NAND3X0 U288 ( .IN1(n418), .IN2(n419), .IN3(n420), .QN(\CARRYB[13][20] ) );
  XOR3X1 U289 ( .IN1(\ab[15][18] ), .IN2(\CARRYB[14][18] ), .IN3(
        \SUMB[14][19] ), .Q(\SUMB[15][18] ) );
  XOR2X1 U290 ( .IN1(\SUMB[17][21] ), .IN2(\ab[18][20] ), .Q(n706) );
  NAND3X0 U291 ( .IN1(n243), .IN2(n244), .IN3(n245), .QN(\CARRYB[17][25] ) );
  NAND3X0 U292 ( .IN1(n898), .IN2(n899), .IN3(n900), .QN(\CARRYB[16][24] ) );
  NAND3X0 U293 ( .IN1(n1181), .IN2(n1182), .IN3(n1183), .QN(\CARRYB[16][21] )
         );
  NAND3X0 U294 ( .IN1(n1361), .IN2(n1362), .IN3(n1363), .QN(\CARRYB[6][13] )
         );
  NAND3X0 U295 ( .IN1(n1324), .IN2(n1325), .IN3(n1326), .QN(\CARRYB[9][13] )
         );
  XOR3X1 U296 ( .IN1(\CARRYB[12][16] ), .IN2(\ab[13][16] ), .IN3(
        \SUMB[12][17] ), .Q(\SUMB[13][16] ) );
  XOR3X1 U297 ( .IN1(\ab[10][15] ), .IN2(\CARRYB[9][15] ), .IN3(\SUMB[9][16] ), 
        .Q(n49) );
  XOR2X1 U298 ( .IN1(n440), .IN2(\SUMB[13][19] ), .Q(\SUMB[14][18] ) );
  NAND3X0 U299 ( .IN1(n522), .IN2(n523), .IN3(n524), .QN(\CARRYB[18][17] ) );
  NAND3X0 U300 ( .IN1(n1158), .IN2(n1159), .IN3(n1160), .QN(\CARRYB[20][19] )
         );
  NAND3X0 U301 ( .IN1(n1029), .IN2(n1030), .IN3(n1031), .QN(\CARRYB[18][26] )
         );
  NAND3X0 U302 ( .IN1(n1578), .IN2(n1579), .IN3(n1580), .QN(\CARRYB[17][30] )
         );
  AND2X1 U303 ( .IN1(\ab[0][14] ), .IN2(\ab[1][13] ), .Q(n1425) );
  XOR2X1 U304 ( .IN1(\ab[1][14] ), .IN2(\ab[0][15] ), .Q(\SUMB[1][14] ) );
  AND2X1 U305 ( .IN1(\ab[0][15] ), .IN2(\ab[1][14] ), .Q(n948) );
  NAND3X0 U306 ( .IN1(n354), .IN2(n355), .IN3(n356), .QN(\CARRYB[3][14] ) );
  XOR2X1 U307 ( .IN1(n943), .IN2(\CARRYB[2][15] ), .Q(\SUMB[3][15] ) );
  NAND3X0 U308 ( .IN1(n1620), .IN2(n1621), .IN3(n1622), .QN(\CARRYB[4][13] )
         );
  NAND3X0 U309 ( .IN1(n190), .IN2(n191), .IN3(n192), .QN(\CARRYB[12][14] ) );
  NAND3X0 U310 ( .IN1(n1110), .IN2(n1111), .IN3(n1112), .QN(\CARRYB[11][15] )
         );
  NAND3X0 U311 ( .IN1(n1682), .IN2(n1683), .IN3(n1684), .QN(\CARRYB[18][14] )
         );
  XOR2X1 U312 ( .IN1(n1157), .IN2(\CARRYB[19][19] ), .Q(\SUMB[20][19] ) );
  NAND3X0 U313 ( .IN1(n1637), .IN2(n1638), .IN3(n1639), .QN(\CARRYB[20][18] )
         );
  NAND3X0 U314 ( .IN1(n1244), .IN2(n1245), .IN3(n1246), .QN(\CARRYB[21][15] )
         );
  XOR2X1 U315 ( .IN1(n1028), .IN2(\SUMB[18][26] ), .Q(\SUMB[19][25] ) );
  XOR2X1 U316 ( .IN1(n242), .IN2(\SUMB[17][25] ), .Q(\SUMB[18][24] ) );
  NAND3X0 U317 ( .IN1(n575), .IN2(n576), .IN3(n577), .QN(\CARRYB[20][20] ) );
  NAND3X0 U318 ( .IN1(n1645), .IN2(n1646), .IN3(n1647), .QN(\CARRYB[12][11] )
         );
  XNOR2X1 U319 ( .IN1(n1310), .IN2(\CARRYB[18][12] ), .Q(\SUMB[19][12] ) );
  NAND3X0 U320 ( .IN1(n465), .IN2(n466), .IN3(n467), .QN(\CARRYB[19][13] ) );
  XOR2X1 U321 ( .IN1(n518), .IN2(\SUMB[17][18] ), .Q(\SUMB[18][17] ) );
  NOR2X0 U322 ( .IN1(n2132), .IN2(n2029), .QN(\ab[22][17] ) );
  NAND3X0 U323 ( .IN1(n888), .IN2(n889), .IN3(n890), .QN(\CARRYB[22][24] ) );
  NAND3X0 U324 ( .IN1(n1375), .IN2(n1376), .IN3(n1377), .QN(\CARRYB[4][12] )
         );
  NAND3X0 U325 ( .IN1(n698), .IN2(n699), .IN3(n700), .QN(\CARRYB[12][10] ) );
  XOR3X1 U326 ( .IN1(\CARRYB[10][11] ), .IN2(\ab[11][11] ), .IN3(
        \SUMB[10][12] ), .Q(\SUMB[11][11] ) );
  XOR2X1 U327 ( .IN1(n1678), .IN2(\CARRYB[13][11] ), .Q(\SUMB[14][11] ) );
  NAND3X0 U328 ( .IN1(n1556), .IN2(n1557), .IN3(n1558), .QN(\CARRYB[15][11] )
         );
  NAND3X0 U329 ( .IN1(n273), .IN2(n274), .IN3(n275), .QN(\CARRYB[16][10] ) );
  NAND3X0 U330 ( .IN1(n979), .IN2(n980), .IN3(n981), .QN(\CARRYB[18][11] ) );
  NAND3X0 U331 ( .IN1(n1067), .IN2(n1068), .IN3(n1069), .QN(\CARRYB[21][10] )
         );
  NAND3X0 U332 ( .IN1(n472), .IN2(n473), .IN3(n474), .QN(\CARRYB[22][11] ) );
  NAND3X0 U333 ( .IN1(n620), .IN2(n621), .IN3(n622), .QN(\CARRYB[22][17] ) );
  NAND3X0 U334 ( .IN1(n1481), .IN2(n1482), .IN3(n1483), .QN(\CARRYB[22][16] )
         );
  NAND3X0 U335 ( .IN1(n1096), .IN2(n1097), .IN3(n1098), .QN(\CARRYB[23][14] )
         );
  NAND3X0 U336 ( .IN1(n1089), .IN2(n1090), .IN3(n1091), .QN(\CARRYB[21][21] )
         );
  NAND3X0 U337 ( .IN1(n1080), .IN2(n1081), .IN3(n1082), .QN(\CARRYB[23][22] )
         );
  XOR2X1 U338 ( .IN1(n763), .IN2(\CARRYB[22][23] ), .Q(\SUMB[23][23] ) );
  NAND3X0 U339 ( .IN1(n764), .IN2(n765), .IN3(n766), .QN(\CARRYB[23][23] ) );
  NAND3X0 U340 ( .IN1(n649), .IN2(n650), .IN3(n651), .QN(\CARRYB[23][25] ) );
  NBUFFX2 U341 ( .INP(n2231), .Z(n2156) );
  NBUFFX2 U342 ( .INP(n2230), .Z(n2154) );
  XOR3X1 U343 ( .IN1(\CARRYB[2][11] ), .IN2(\ab[3][11] ), .IN3(\SUMB[2][12] ), 
        .Q(\SUMB[3][11] ) );
  XOR2X1 U344 ( .IN1(\ab[4][11] ), .IN2(\SUMB[3][12] ), .Q(n1076) );
  NAND3X0 U345 ( .IN1(n718), .IN2(n719), .IN3(n720), .QN(\CARRYB[6][10] ) );
  NAND3X0 U346 ( .IN1(n266), .IN2(n267), .IN3(n268), .QN(\CARRYB[14][10] ) );
  NOR2X0 U347 ( .IN1(n2150), .IN2(n2038), .QN(\ab[19][10] ) );
  NAND3X0 U348 ( .IN1(n602), .IN2(n603), .IN3(n604), .QN(\CARRYB[23][16] ) );
  NAND3X0 U349 ( .IN1(n434), .IN2(n435), .IN3(n436), .QN(\CARRYB[23][20] ) );
  NAND3X0 U350 ( .IN1(n1083), .IN2(n1084), .IN3(n1085), .QN(\CARRYB[24][21] )
         );
  NAND3X0 U351 ( .IN1(n1512), .IN2(n1513), .IN3(n1514), .QN(\CARRYB[24][24] )
         );
  NAND3X0 U352 ( .IN1(n335), .IN2(n336), .IN3(n337), .QN(\CARRYB[23][28] ) );
  NAND3X0 U353 ( .IN1(n1259), .IN2(n1260), .IN3(n1261), .QN(\CARRYB[23][29] )
         );
  AND2X1 U354 ( .IN1(\ab[0][9] ), .IN2(\ab[1][8] ), .Q(n1354) );
  XOR2X1 U355 ( .IN1(\ab[1][9] ), .IN2(\ab[0][10] ), .Q(\SUMB[1][9] ) );
  AND2X1 U356 ( .IN1(B[10]), .IN2(A[1]), .Q(\ab[1][10] ) );
  NAND3X0 U357 ( .IN1(n1223), .IN2(n1224), .IN3(n1225), .QN(\CARRYB[3][8] ) );
  NOR2X0 U358 ( .IN1(n2157), .IN2(n2067), .QN(\ab[10][8] ) );
  XOR2X1 U359 ( .IN1(\ab[15][7] ), .IN2(\SUMB[14][8] ), .Q(n1045) );
  NAND3X0 U360 ( .IN1(n121), .IN2(n122), .IN3(n123), .QN(\CARRYB[15][8] ) );
  XOR2X1 U361 ( .IN1(n1771), .IN2(\CARRYB[17][9] ), .Q(\SUMB[18][9] ) );
  NAND3X0 U362 ( .IN1(n1292), .IN2(n1293), .IN3(n1294), .QN(\CARRYB[18][8] )
         );
  NAND3X0 U363 ( .IN1(n277), .IN2(n278), .IN3(n279), .QN(\CARRYB[17][10] ) );
  NAND3X0 U364 ( .IN1(n1772), .IN2(n1773), .IN3(n1774), .QN(\CARRYB[18][9] )
         );
  NAND3X0 U365 ( .IN1(n1843), .IN2(n1844), .IN3(n1845), .QN(\CARRYB[23][8] )
         );
  NAND3X0 U366 ( .IN1(n1471), .IN2(n1472), .IN3(n1473), .QN(\CARRYB[25][15] )
         );
  NAND3X0 U367 ( .IN1(n1731), .IN2(n1732), .IN3(n1733), .QN(\CARRYB[25][13] )
         );
  XOR2X1 U368 ( .IN1(n1102), .IN2(\CARRYB[24][14] ), .Q(\SUMB[25][14] ) );
  XOR2X1 U369 ( .IN1(n1470), .IN2(\SUMB[25][15] ), .Q(\SUMB[26][14] ) );
  NAND3X0 U370 ( .IN1(n1147), .IN2(n1148), .IN3(n1149), .QN(\CARRYB[26][19] )
         );
  XOR2X1 U371 ( .IN1(n1538), .IN2(\CARRYB[24][22] ), .Q(\SUMB[25][22] ) );
  XOR2X1 U372 ( .IN1(n1518), .IN2(\CARRYB[24][23] ), .Q(\SUMB[25][23] ) );
  NAND3X0 U373 ( .IN1(n1539), .IN2(n1540), .IN3(n1541), .QN(\CARRYB[25][22] )
         );
  XNOR2X1 U374 ( .IN1(n974), .IN2(\CARRYB[24][26] ), .Q(n836) );
  NAND3X0 U375 ( .IN1(n1571), .IN2(n1572), .IN3(n1573), .QN(\CARRYB[25][30] )
         );
  XOR2X1 U376 ( .IN1(n1778), .IN2(\CARRYB[6][9] ), .Q(\SUMB[7][9] ) );
  NOR2X0 U377 ( .IN1(n2159), .IN2(n2067), .QN(\ab[10][7] ) );
  NAND3X0 U378 ( .IN1(n593), .IN2(n594), .IN3(n595), .QN(\CARRYB[19][7] ) );
  XOR2X1 U379 ( .IN1(n1752), .IN2(\CARRYB[20][7] ), .Q(\SUMB[21][7] ) );
  NAND3X0 U380 ( .IN1(n1753), .IN2(n1754), .IN3(n1755), .QN(\CARRYB[21][7] )
         );
  XOR2X1 U381 ( .IN1(n1842), .IN2(\CARRYB[22][8] ), .Q(\SUMB[23][8] ) );
  NAND3X0 U382 ( .IN1(n1690), .IN2(n1691), .IN3(n1692), .QN(\CARRYB[27][6] )
         );
  NAND3X0 U383 ( .IN1(n806), .IN2(n807), .IN3(n808), .QN(\CARRYB[26][10] ) );
  XOR2X1 U384 ( .IN1(n1727), .IN2(\CARRYB[27][13] ), .Q(\SUMB[28][13] ) );
  XOR2X1 U385 ( .IN1(n1671), .IN2(\CARRYB[26][16] ), .Q(\SUMB[27][16] ) );
  NAND3X0 U386 ( .IN1(n1532), .IN2(n1533), .IN3(n1534), .QN(\CARRYB[27][15] )
         );
  NAND3X0 U387 ( .IN1(n229), .IN2(n230), .IN3(n231), .QN(\CARRYB[27][17] ) );
  NAND3X0 U388 ( .IN1(n226), .IN2(n227), .IN3(n228), .QN(\CARRYB[26][18] ) );
  XOR2X1 U389 ( .IN1(n1508), .IN2(\CARRYB[25][24] ), .Q(\SUMB[26][24] ) );
  NAND3X0 U390 ( .IN1(n131), .IN2(n132), .IN3(n133), .QN(\CARRYB[26][23] ) );
  NAND3X0 U391 ( .IN1(n1509), .IN2(n1510), .IN3(n1511), .QN(\CARRYB[26][24] )
         );
  NAND3X0 U392 ( .IN1(n1429), .IN2(n1430), .IN3(n1431), .QN(\CARRYB[25][26] )
         );
  NAND3X0 U393 ( .IN1(n1563), .IN2(n1564), .IN3(n1565), .QN(\CARRYB[26][30] )
         );
  XOR2X1 U394 ( .IN1(n1713), .IN2(\CARRYB[2][6] ), .Q(\SUMB[3][6] ) );
  NAND3X0 U395 ( .IN1(n1714), .IN2(n1715), .IN3(n1716), .QN(\CARRYB[3][6] ) );
  XOR2X1 U396 ( .IN1(n1222), .IN2(\CARRYB[2][8] ), .Q(\SUMB[3][8] ) );
  NAND3X0 U397 ( .IN1(n1145), .IN2(n1144), .IN3(n1146), .QN(\CARRYB[7][7] ) );
  XOR2X1 U398 ( .IN1(n1759), .IN2(\CARRYB[11][7] ), .Q(\SUMB[12][7] ) );
  NAND3X0 U399 ( .IN1(n747), .IN2(n748), .IN3(n749), .QN(\CARRYB[13][5] ) );
  XOR2X1 U400 ( .IN1(n952), .IN2(\CARRYB[16][5] ), .Q(\SUMB[17][5] ) );
  NAND3X0 U401 ( .IN1(n596), .IN2(n597), .IN3(n598), .QN(\CARRYB[20][6] ) );
  NAND3X0 U402 ( .IN1(n581), .IN2(n582), .IN3(n583), .QN(\CARRYB[21][6] ) );
  NAND3X0 U403 ( .IN1(n670), .IN2(n671), .IN3(n672), .QN(\CARRYB[24][5] ) );
  NAND3X0 U404 ( .IN1(n674), .IN2(n675), .IN3(n676), .QN(\CARRYB[25][5] ) );
  NAND3X0 U405 ( .IN1(n287), .IN2(n288), .IN3(n289), .QN(\CARRYB[26][5] ) );
  NAND3X0 U406 ( .IN1(n291), .IN2(n292), .IN3(n293), .QN(\CARRYB[27][5] ) );
  XOR2X1 U407 ( .IN1(n1908), .IN2(\CARRYB[28][5] ), .Q(\SUMB[29][5] ) );
  XOR2X1 U408 ( .IN1(n805), .IN2(\SUMB[26][10] ), .Q(\SUMB[27][9] ) );
  NAND3X0 U409 ( .IN1(n504), .IN2(n505), .IN3(n506), .QN(\CARRYB[28][7] ) );
  NAND3X0 U410 ( .IN1(n302), .IN2(n303), .IN3(n304), .QN(\CARRYB[27][14] ) );
  NAND3X0 U411 ( .IN1(n1883), .IN2(n1884), .IN3(n1885), .QN(\CARRYB[29][12] )
         );
  NAND3X0 U412 ( .IN1(n221), .IN2(n222), .IN3(n223), .QN(\CARRYB[28][16] ) );
  NAND3X0 U413 ( .IN1(n395), .IN2(n396), .IN3(n397), .QN(\CARRYB[28][19] ) );
  NAND3X0 U414 ( .IN1(n1418), .IN2(n1419), .IN3(n1420), .QN(\CARRYB[28][27] )
         );
  NAND3X0 U415 ( .IN1(n539), .IN2(n540), .IN3(n541), .QN(\CARRYB[3][5] ) );
  XOR2X1 U416 ( .IN1(n1829), .IN2(\CARRYB[11][4] ), .Q(\SUMB[12][4] ) );
  XOR2X1 U417 ( .IN1(n592), .IN2(\SUMB[19][7] ), .Q(\SUMB[20][6] ) );
  XOR2X1 U418 ( .IN1(n673), .IN2(\CARRYB[24][5] ), .Q(\SUMB[25][5] ) );
  NAND3X0 U419 ( .IN1(n1791), .IN2(n1792), .IN3(n1793), .QN(\CARRYB[27][3] )
         );
  NAND3X0 U420 ( .IN1(n1783), .IN2(n1784), .IN3(n1785), .QN(\CARRYB[28][3] )
         );
  NAND3X0 U421 ( .IN1(n1697), .IN2(n1698), .IN3(n1699), .QN(\CARRYB[29][6] )
         );
  NOR2X0 U422 ( .IN1(B[7]), .IN2(n2004), .QN(\ab[31][7] ) );
  NOR2X0 U423 ( .IN1(B[10]), .IN2(n2004), .QN(\ab[31][10] ) );
  NAND3X0 U424 ( .IN1(n299), .IN2(n300), .IN3(n301), .QN(\CARRYB[29][14] ) );
  XOR2X1 U425 ( .IN1(n786), .IN2(\CARRYB[28][15] ), .Q(\SUMB[29][15] ) );
  NAND3X0 U426 ( .IN1(n239), .IN2(n240), .IN3(n241), .QN(\CARRYB[30][22] ) );
  NAND3X0 U427 ( .IN1(n881), .IN2(n882), .IN3(n883), .QN(\CARRYB[30][21] ) );
  NAND3X0 U428 ( .IN1(n1422), .IN2(n1423), .IN3(n1424), .QN(\CARRYB[29][27] )
         );
  NAND3X0 U429 ( .IN1(n1567), .IN2(n1568), .IN3(n1569), .QN(\CARRYB[27][30] )
         );
  NBUFFX2 U430 ( .INP(n2236), .Z(n2167) );
  XOR2X1 U431 ( .IN1(n1200), .IN2(\CARRYB[3][4] ), .Q(\SUMB[4][4] ) );
  XOR2X1 U432 ( .IN1(n106), .IN2(\CARRYB[6][5] ), .Q(\SUMB[7][5] ) );
  XOR2X1 U433 ( .IN1(n736), .IN2(\CARRYB[12][3] ), .Q(\SUMB[13][3] ) );
  NAND3X0 U434 ( .IN1(n1798), .IN2(n1799), .IN3(n1800), .QN(\CARRYB[16][3] )
         );
  NAND3X0 U435 ( .IN1(n1128), .IN2(n1129), .IN3(n1130), .QN(\CARRYB[19][3] )
         );
  XOR2X1 U436 ( .IN1(n628), .IN2(\CARRYB[20][3] ), .Q(\SUMB[21][3] ) );
  NAND3X0 U437 ( .IN1(n1344), .IN2(n1345), .IN3(n1346), .QN(\CARRYB[23][3] )
         );
  NAND3X0 U438 ( .IN1(n1334), .IN2(n1335), .IN3(n1336), .QN(\CARRYB[30][2] )
         );
  XOR2X1 U439 ( .IN1(n45), .IN2(\CARRYB[30][3] ), .Q(\SUMB[31][3] ) );
  XOR2X1 U440 ( .IN1(n283), .IN2(\CARRYB[30][4] ), .Q(\SUMB[31][4] ) );
  NAND3X0 U441 ( .IN1(n284), .IN2(n285), .IN3(n286), .QN(\CARRYB[31][4] ) );
  XNOR2X1 U442 ( .IN1(n1311), .IN2(\CARRYB[29][6] ), .Q(\SUMB[30][6] ) );
  NAND3X0 U443 ( .IN1(n1700), .IN2(n1701), .IN3(n1702), .QN(\CARRYB[30][6] )
         );
  XOR2X1 U444 ( .IN1(n1745), .IN2(\CARRYB[29][7] ), .Q(\SUMB[30][7] ) );
  NAND3X0 U445 ( .IN1(n1742), .IN2(n1743), .IN3(n1744), .QN(\CARRYB[31][7] )
         );
  NAND3X0 U446 ( .IN1(n1833), .IN2(n1834), .IN3(n1835), .QN(\CARRYB[31][8] )
         );
  INVX0 U447 ( .INP(\ab[31][10] ), .ZN(n176) );
  NAND3X0 U448 ( .IN1(n1227), .IN2(n1228), .IN3(n1229), .QN(\CARRYB[31][11] )
         );
  NAND3X0 U449 ( .IN1(n1887), .IN2(n1888), .IN3(n1889), .QN(\CARRYB[30][12] )
         );
  XOR2X1 U450 ( .IN1(n868), .IN2(\CARRYB[29][16] ), .Q(\SUMB[30][16] ) );
  NAND3X0 U451 ( .IN1(n869), .IN2(n870), .IN3(n871), .QN(\CARRYB[30][16] ) );
  XOR2X1 U452 ( .IN1(n1657), .IN2(\CARRYB[29][17] ), .Q(\SUMB[30][17] ) );
  NAND3X0 U453 ( .IN1(n1658), .IN2(n1659), .IN3(n1660), .QN(\CARRYB[30][17] )
         );
  XOR2X1 U454 ( .IN1(n759), .IN2(\CARRYB[29][20] ), .Q(\SUMB[30][20] ) );
  XOR2X1 U455 ( .IN1(n884), .IN2(\CARRYB[30][21] ), .Q(\SUMB[31][21] ) );
  NAND3X0 U456 ( .IN1(n760), .IN2(n761), .IN3(n762), .QN(\CARRYB[30][20] ) );
  NAND3X0 U457 ( .IN1(n885), .IN2(n886), .IN3(n887), .QN(\CARRYB[31][21] ) );
  XOR2X1 U458 ( .IN1(n1487), .IN2(\CARRYB[30][24] ), .Q(\SUMB[31][24] ) );
  XOR2X1 U459 ( .IN1(n1442), .IN2(\CARRYB[30][25] ), .Q(\SUMB[31][25] ) );
  NAND3X0 U460 ( .IN1(n1488), .IN2(n1489), .IN3(n1490), .QN(\CARRYB[31][24] )
         );
  NAND3X0 U461 ( .IN1(n1443), .IN2(n1444), .IN3(n1445), .QN(\CARRYB[31][25] )
         );
  NAND3X0 U462 ( .IN1(n664), .IN2(n665), .IN3(n666), .QN(\CARRYB[3][2] ) );
  XOR2X1 U463 ( .IN1(n861), .IN2(\CARRYB[5][3] ), .Q(\SUMB[6][3] ) );
  XNOR2X1 U464 ( .IN1(n755), .IN2(\CARRYB[15][2] ), .Q(\SUMB[16][2] ) );
  NAND3X0 U465 ( .IN1(n1210), .IN2(n1211), .IN3(n1212), .QN(\CARRYB[17][2] )
         );
  NAND3X0 U466 ( .IN1(n1954), .IN2(n1955), .IN3(n1956), .QN(\CARRYB[21][0] )
         );
  NAND3X0 U467 ( .IN1(n1208), .IN2(n1207), .IN3(n1209), .QN(\CARRYB[20][2] )
         );
  XOR3X1 U468 ( .IN1(\ab[20][3] ), .IN2(\CARRYB[19][3] ), .IN3(\SUMB[19][4] ), 
        .Q(\SUMB[20][3] ) );
  NAND3X0 U469 ( .IN1(n1929), .IN2(n1930), .IN3(n1931), .QN(\CARRYB[24][2] )
         );
  NAND3X0 U470 ( .IN1(n1340), .IN2(n1341), .IN3(n1342), .QN(\CARRYB[25][3] )
         );
  XOR2X1 U471 ( .IN1(n1333), .IN2(\CARRYB[29][2] ), .Q(\SUMB[30][2] ) );
  XOR2X1 U472 ( .IN1(\CARRYB[31][2] ), .IN2(\SUMB[31][3] ), .Q(\A1[32] ) );
  XOR2X1 U473 ( .IN1(\CARRYB[31][3] ), .IN2(\SUMB[31][4] ), .Q(\A1[33] ) );
  XOR2X1 U474 ( .IN1(\CARRYB[31][6] ), .IN2(\SUMB[31][7] ), .Q(\A1[36] ) );
  XOR2X1 U475 ( .IN1(\CARRYB[31][7] ), .IN2(\SUMB[31][8] ), .Q(\A1[37] ) );
  XOR2X1 U476 ( .IN1(\CARRYB[31][8] ), .IN2(\SUMB[31][9] ), .Q(\A1[38] ) );
  AND2X1 U477 ( .IN1(\CARRYB[31][8] ), .IN2(\SUMB[31][9] ), .Q(n1981) );
  AND2X1 U478 ( .IN1(\CARRYB[31][9] ), .IN2(\SUMB[31][10] ), .Q(n1976) );
  XOR2X1 U479 ( .IN1(\CARRYB[31][10] ), .IN2(\SUMB[31][11] ), .Q(\A1[40] ) );
  AND2X1 U480 ( .IN1(\SUMB[31][21] ), .IN2(\CARRYB[31][20] ), .Q(n1993) );
  NBUFFX4 U481 ( .INP(B[30]), .Z(n546) );
  AND2X1 U482 ( .IN1(B[0]), .IN2(A[1]), .Q(\ab[1][0] ) );
  XOR2X1 U483 ( .IN1(n663), .IN2(\CARRYB[2][2] ), .Q(\SUMB[3][2] ) );
  NAND3X0 U484 ( .IN1(n1867), .IN2(n1868), .IN3(n1869), .QN(\CARRYB[11][1] )
         );
  XOR3X1 U485 ( .IN1(\ab[14][1] ), .IN2(\CARRYB[13][1] ), .IN3(\SUMB[13][2] ), 
        .Q(\SUMB[14][1] ) );
  NOR2X0 U486 ( .IN1(n2173), .IN2(n2050), .QN(\ab[15][0] ) );
  NOR2X0 U487 ( .IN1(n2173), .IN2(n2044), .QN(\ab[17][0] ) );
  XOR2X1 U488 ( .IN1(n535), .IN2(n18), .Q(\SUMB[21][1] ) );
  NAND3X0 U489 ( .IN1(n1135), .IN2(n1136), .IN3(n1137), .QN(\CARRYB[23][1] )
         );
  NAND3X0 U490 ( .IN1(n324), .IN2(n325), .IN3(n326), .QN(\CARRYB[27][1] ) );
  XOR2X1 U491 ( .IN1(n320), .IN2(\CARRYB[28][1] ), .Q(\SUMB[29][1] ) );
  NAND3X0 U492 ( .IN1(n1965), .IN2(n1966), .IN3(n1967), .QN(\CARRYB[10][0] )
         );
  NAND3X0 U493 ( .IN1(n63), .IN2(n64), .IN3(n65), .QN(\CARRYB[15][0] ) );
  XOR2X1 U494 ( .IN1(\ab[19][0] ), .IN2(\SUMB[18][1] ), .Q(n921) );
  NAND3X0 U495 ( .IN1(n922), .IN2(n923), .IN3(n924), .QN(\CARRYB[19][0] ) );
  INVX0 U496 ( .INP(\CARRYB[31][31] ), .ZN(n2175) );
  NBUFFX2 U497 ( .INP(n2232), .Z(n2159) );
  AND2X1 U498 ( .IN1(\ab[0][5] ), .IN2(\ab[1][4] ), .Q(n3) );
  AND2X1 U499 ( .IN1(\ab[0][2] ), .IN2(\ab[1][1] ), .Q(n4) );
  AND2X1 U500 ( .IN1(\ab[0][18] ), .IN2(\ab[1][17] ), .Q(n5) );
  AND2X1 U501 ( .IN1(\ab[0][20] ), .IN2(\ab[1][19] ), .Q(n6) );
  AND2X1 U502 ( .IN1(\ab[0][29] ), .IN2(\ab[1][28] ), .Q(n7) );
  AND2X1 U503 ( .IN1(\ab[0][21] ), .IN2(\ab[1][20] ), .Q(n8) );
  AND2X1 U504 ( .IN1(\ab[0][13] ), .IN2(\ab[1][12] ), .Q(n9) );
  AND2X1 U505 ( .IN1(\ab[0][26] ), .IN2(\ab[1][25] ), .Q(n10) );
  AND2X1 U506 ( .IN1(\ab[0][25] ), .IN2(\ab[1][24] ), .Q(n11) );
  AND2X1 U507 ( .IN1(\ab[1][6] ), .IN2(\ab[0][7] ), .Q(n12) );
  AND2X1 U508 ( .IN1(\ab[0][1] ), .IN2(\ab[1][0] ), .Q(n13) );
  AND2X1 U509 ( .IN1(\ab[0][19] ), .IN2(\ab[1][18] ), .Q(n14) );
  AND2X1 U510 ( .IN1(\ab[0][16] ), .IN2(\ab[1][15] ), .Q(n15) );
  AND2X1 U511 ( .IN1(\CARRYB[31][30] ), .IN2(\SUMB[31][31] ), .Q(n16) );
  INVX0 U512 ( .INP(\ab[24][24] ), .ZN(n659) );
  INVX0 U513 ( .INP(\ab[25][3] ), .ZN(n23) );
  INVX0 U514 ( .INP(\ab[24][22] ), .ZN(n1027) );
  XNOR2X1 U515 ( .IN1(n17), .IN2(\SUMB[7][22] ), .Q(\SUMB[8][21] ) );
  XNOR2X1 U516 ( .IN1(\ab[8][21] ), .IN2(\CARRYB[7][21] ), .Q(n17) );
  NAND3X1 U517 ( .IN1(n532), .IN2(n533), .IN3(n534), .QN(n18) );
  XOR2X1 U518 ( .IN1(n327), .IN2(\CARRYB[9][7] ), .Q(\SUMB[10][7] ) );
  NAND2X0 U519 ( .IN1(\ab[6][9] ), .IN2(\CARRYB[5][9] ), .QN(n1775) );
  NAND3X1 U520 ( .IN1(n1433), .IN2(n1432), .IN3(n1434), .QN(n19) );
  NBUFFX2 U521 ( .INP(\SUMB[8][22] ), .Z(n57) );
  INVX0 U522 ( .INP(n2134), .ZN(n20) );
  DELLN1X2 U523 ( .INP(n2223), .Z(n2134) );
  XNOR2X1 U524 ( .IN1(n21), .IN2(\CARRYB[13][5] ), .Q(\SUMB[14][5] ) );
  XNOR2X1 U525 ( .IN1(\ab[14][5] ), .IN2(\SUMB[13][6] ), .Q(n21) );
  XOR2X1 U526 ( .IN1(n23), .IN2(\SUMB[24][4] ), .Q(n394) );
  XOR2X1 U527 ( .IN1(\ab[1][23] ), .IN2(\ab[0][24] ), .Q(\SUMB[1][23] ) );
  NAND2X0 U528 ( .IN1(\ab[2][22] ), .IN2(\SUMB[1][23] ), .QN(n387) );
  NAND3X0 U529 ( .IN1(n386), .IN2(n387), .IN3(n388), .QN(\CARRYB[2][22] ) );
  XOR2X2 U530 ( .IN1(\ab[1][12] ), .IN2(\ab[0][13] ), .Q(\SUMB[1][12] ) );
  XOR3X1 U531 ( .IN1(\CARRYB[14][9] ), .IN2(\ab[15][9] ), .IN3(\SUMB[14][10] ), 
        .Q(\SUMB[15][9] ) );
  NAND2X1 U532 ( .IN1(\CARRYB[14][9] ), .IN2(\SUMB[14][10] ), .QN(n24) );
  NAND2X1 U533 ( .IN1(\CARRYB[14][9] ), .IN2(\ab[15][9] ), .QN(n25) );
  NAND2X1 U534 ( .IN1(\SUMB[14][10] ), .IN2(\ab[15][9] ), .QN(n26) );
  NAND3X0 U535 ( .IN1(n24), .IN2(n25), .IN3(n26), .QN(\CARRYB[15][9] ) );
  NAND3X0 U536 ( .IN1(n118), .IN2(n119), .IN3(n120), .QN(\CARRYB[14][9] ) );
  NAND2X0 U537 ( .IN1(\ab[9][21] ), .IN2(n57), .QN(n310) );
  INVX0 U538 ( .INP(n2145), .ZN(n28) );
  XNOR2X2 U539 ( .IN1(n177), .IN2(\SUMB[10][19] ), .Q(\SUMB[11][18] ) );
  XNOR2X2 U540 ( .IN1(n29), .IN2(\CARRYB[11][9] ), .Q(\SUMB[12][9] ) );
  XNOR2X1 U541 ( .IN1(\ab[12][9] ), .IN2(\SUMB[11][10] ), .Q(n29) );
  XOR3X1 U542 ( .IN1(\SUMB[7][17] ), .IN2(\ab[8][16] ), .IN3(\CARRYB[7][16] ), 
        .Q(\SUMB[8][16] ) );
  NAND2X0 U543 ( .IN1(\SUMB[7][17] ), .IN2(\CARRYB[7][16] ), .QN(n30) );
  NAND2X0 U544 ( .IN1(\SUMB[7][17] ), .IN2(\ab[8][16] ), .QN(n31) );
  NAND2X0 U545 ( .IN1(\CARRYB[7][16] ), .IN2(\ab[8][16] ), .QN(n32) );
  XOR3X1 U546 ( .IN1(\CARRYB[12][15] ), .IN2(\ab[13][15] ), .IN3(
        \SUMB[12][16] ), .Q(\SUMB[13][15] ) );
  NAND2X1 U547 ( .IN1(\CARRYB[12][15] ), .IN2(\SUMB[12][16] ), .QN(n33) );
  NAND2X0 U548 ( .IN1(\CARRYB[12][15] ), .IN2(\ab[13][15] ), .QN(n34) );
  NAND2X1 U549 ( .IN1(\SUMB[12][16] ), .IN2(\ab[13][15] ), .QN(n35) );
  NAND3X0 U550 ( .IN1(n33), .IN2(n34), .IN3(n35), .QN(\CARRYB[13][15] ) );
  NAND3X1 U551 ( .IN1(n1063), .IN2(n1064), .IN3(n1065), .QN(\CARRYB[9][11] )
         );
  XOR3X1 U552 ( .IN1(\SUMB[11][17] ), .IN2(\ab[12][16] ), .IN3(
        \CARRYB[11][16] ), .Q(\SUMB[12][16] ) );
  NAND2X0 U553 ( .IN1(\SUMB[11][17] ), .IN2(\CARRYB[11][16] ), .QN(n36) );
  NAND2X0 U554 ( .IN1(\SUMB[11][17] ), .IN2(\ab[12][16] ), .QN(n37) );
  NAND2X1 U555 ( .IN1(\CARRYB[11][16] ), .IN2(\ab[12][16] ), .QN(n38) );
  NAND3X0 U556 ( .IN1(n36), .IN2(n37), .IN3(n38), .QN(\CARRYB[12][16] ) );
  NAND3X0 U557 ( .IN1(n1312), .IN2(n1313), .IN3(n1314), .QN(\CARRYB[11][16] )
         );
  XOR2X1 U558 ( .IN1(n1233), .IN2(\CARRYB[10][17] ), .Q(\SUMB[11][17] ) );
  XNOR2X2 U559 ( .IN1(n39), .IN2(\CARRYB[7][12] ), .Q(\SUMB[8][12] ) );
  XNOR2X1 U560 ( .IN1(\ab[8][12] ), .IN2(\SUMB[7][13] ), .Q(n39) );
  XNOR2X2 U561 ( .IN1(n40), .IN2(\CARRYB[8][11] ), .Q(\SUMB[9][11] ) );
  XNOR2X1 U562 ( .IN1(\SUMB[8][12] ), .IN2(\ab[9][11] ), .Q(n40) );
  DELLN2X2 U563 ( .INP(n2223), .Z(n2136) );
  NAND2X0 U564 ( .IN1(\ab[11][10] ), .IN2(\CARRYB[10][10] ), .QN(n695) );
  NAND2X0 U565 ( .IN1(\CARRYB[16][13] ), .IN2(\ab[17][13] ), .QN(n1316) );
  NAND2X0 U566 ( .IN1(\ab[18][13] ), .IN2(\CARRYB[17][13] ), .QN(n461) );
  XOR2X2 U567 ( .IN1(\ab[1][26] ), .IN2(\ab[0][27] ), .Q(\SUMB[1][26] ) );
  XNOR2X2 U568 ( .IN1(n41), .IN2(\SUMB[14][9] ), .Q(\SUMB[15][8] ) );
  XNOR2X1 U569 ( .IN1(\ab[15][8] ), .IN2(\CARRYB[14][8] ), .Q(n41) );
  AND2X1 U570 ( .IN1(B[28]), .IN2(n599), .Q(\ab[0][28] ) );
  NAND3X1 U571 ( .IN1(n1890), .IN2(n1891), .IN3(n1892), .QN(\CARRYB[17][12] )
         );
  NAND2X0 U572 ( .IN1(\SUMB[16][13] ), .IN2(\ab[17][12] ), .QN(n1892) );
  NAND2X0 U573 ( .IN1(\CARRYB[16][12] ), .IN2(\SUMB[16][13] ), .QN(n1890) );
  NAND2X0 U574 ( .IN1(\CARRYB[10][16] ), .IN2(\ab[11][16] ), .QN(n1313) );
  NAND2X0 U575 ( .IN1(\ab[12][8] ), .IN2(\SUMB[11][9] ), .QN(n1847) );
  XOR3X1 U576 ( .IN1(\ab[30][3] ), .IN2(\CARRYB[29][3] ), .IN3(\SUMB[29][4] ), 
        .Q(\SUMB[30][3] ) );
  NAND2X1 U577 ( .IN1(\ab[30][3] ), .IN2(\CARRYB[29][3] ), .QN(n42) );
  NAND2X1 U578 ( .IN1(\ab[30][3] ), .IN2(\SUMB[29][4] ), .QN(n43) );
  NAND2X0 U579 ( .IN1(\CARRYB[29][3] ), .IN2(\SUMB[29][4] ), .QN(n44) );
  NAND3X0 U580 ( .IN1(n42), .IN2(n43), .IN3(n44), .QN(\CARRYB[30][3] ) );
  XOR2X1 U581 ( .IN1(\ab[31][3] ), .IN2(\SUMB[30][4] ), .Q(n45) );
  NAND2X0 U582 ( .IN1(\ab[31][3] ), .IN2(\SUMB[30][4] ), .QN(n46) );
  NAND2X0 U583 ( .IN1(\ab[31][3] ), .IN2(\CARRYB[30][3] ), .QN(n47) );
  NAND2X0 U584 ( .IN1(\SUMB[30][4] ), .IN2(\CARRYB[30][3] ), .QN(n48) );
  NAND3X0 U585 ( .IN1(n46), .IN2(n47), .IN3(n48), .QN(\CARRYB[31][3] ) );
  XOR3X1 U586 ( .IN1(\SUMB[6][17] ), .IN2(\ab[7][16] ), .IN3(\CARRYB[6][16] ), 
        .Q(\SUMB[7][16] ) );
  NAND2X1 U587 ( .IN1(\SUMB[6][17] ), .IN2(\CARRYB[6][16] ), .QN(n50) );
  NAND2X0 U588 ( .IN1(\SUMB[6][17] ), .IN2(\ab[7][16] ), .QN(n51) );
  NAND2X1 U589 ( .IN1(\CARRYB[6][16] ), .IN2(\ab[7][16] ), .QN(n52) );
  NAND3X0 U590 ( .IN1(n986), .IN2(n987), .IN3(n988), .QN(\CARRYB[6][16] ) );
  XOR2X1 U591 ( .IN1(\ab[1][3] ), .IN2(\ab[0][4] ), .Q(\SUMB[1][3] ) );
  XOR2X1 U592 ( .IN1(\ab[12][21] ), .IN2(\SUMB[11][22] ), .Q(n53) );
  XOR2X1 U593 ( .IN1(n53), .IN2(\CARRYB[11][21] ), .Q(\SUMB[12][21] ) );
  NAND2X0 U594 ( .IN1(\CARRYB[11][21] ), .IN2(\SUMB[11][22] ), .QN(n54) );
  NAND2X0 U595 ( .IN1(\CARRYB[11][21] ), .IN2(\ab[12][21] ), .QN(n55) );
  NAND2X1 U596 ( .IN1(\SUMB[11][22] ), .IN2(\ab[12][21] ), .QN(n56) );
  NAND3X0 U597 ( .IN1(n54), .IN2(n55), .IN3(n56), .QN(\CARRYB[12][21] ) );
  XOR3X1 U598 ( .IN1(n61), .IN2(\ab[10][8] ), .IN3(\CARRYB[9][8] ), .Q(
        \SUMB[10][8] ) );
  NAND2X0 U599 ( .IN1(\CARRYB[9][8] ), .IN2(n61), .QN(n58) );
  NAND2X0 U600 ( .IN1(\SUMB[9][9] ), .IN2(\ab[10][8] ), .QN(n59) );
  NAND2X0 U601 ( .IN1(\CARRYB[9][8] ), .IN2(\ab[10][8] ), .QN(n60) );
  NAND3X1 U602 ( .IN1(n58), .IN2(n60), .IN3(n59), .QN(\CARRYB[10][8] ) );
  XOR2X1 U603 ( .IN1(n371), .IN2(\SUMB[8][10] ), .Q(n61) );
  NAND3X0 U604 ( .IN1(n643), .IN2(n644), .IN3(n645), .QN(\CARRYB[9][8] ) );
  DELLN1X2 U605 ( .INP(n2220), .Z(n2126) );
  NAND3X1 U606 ( .IN1(n162), .IN2(n163), .IN3(n164), .QN(\CARRYB[6][23] ) );
  NAND2X0 U607 ( .IN1(\ab[20][1] ), .IN2(\CARRYB[19][1] ), .QN(n532) );
  XOR2X2 U608 ( .IN1(\ab[1][4] ), .IN2(\ab[0][5] ), .Q(\SUMB[1][4] ) );
  NAND3X1 U609 ( .IN1(n918), .IN2(n919), .IN3(n920), .QN(n62) );
  XOR3X1 U610 ( .IN1(\CARRYB[14][0] ), .IN2(\ab[15][0] ), .IN3(\SUMB[14][1] ), 
        .Q(\A1[13] ) );
  NAND2X0 U611 ( .IN1(\CARRYB[14][0] ), .IN2(\SUMB[14][1] ), .QN(n63) );
  NAND2X0 U612 ( .IN1(\CARRYB[14][0] ), .IN2(\ab[15][0] ), .QN(n64) );
  NAND2X0 U613 ( .IN1(\SUMB[14][1] ), .IN2(\ab[15][0] ), .QN(n65) );
  XOR3X1 U614 ( .IN1(\CARRYB[5][0] ), .IN2(\ab[6][0] ), .IN3(\SUMB[5][1] ), 
        .Q(\A1[4] ) );
  NAND2X0 U615 ( .IN1(\CARRYB[5][0] ), .IN2(\SUMB[5][1] ), .QN(n66) );
  NAND2X0 U616 ( .IN1(\CARRYB[5][0] ), .IN2(\ab[6][0] ), .QN(n67) );
  NAND2X1 U617 ( .IN1(\SUMB[5][1] ), .IN2(\ab[6][0] ), .QN(n68) );
  NAND3X0 U618 ( .IN1(n66), .IN2(n67), .IN3(n68), .QN(\CARRYB[6][0] ) );
  DELLN1X2 U619 ( .INP(n2238), .Z(n2171) );
  DELLN1X2 U620 ( .INP(n2219), .Z(n2124) );
  XNOR2X2 U621 ( .IN1(n69), .IN2(\SUMB[18][7] ), .Q(\SUMB[19][6] ) );
  XNOR2X1 U622 ( .IN1(\ab[19][6] ), .IN2(\CARRYB[18][6] ), .Q(n69) );
  NAND2X0 U623 ( .IN1(n1425), .IN2(\ab[2][13] ), .QN(n1379) );
  NAND3X1 U624 ( .IN1(n1378), .IN2(n1379), .IN3(n1380), .QN(\CARRYB[2][13] )
         );
  NAND2X0 U625 ( .IN1(\CARRYB[8][0] ), .IN2(\SUMB[8][1] ), .QN(n1963) );
  NAND2X0 U626 ( .IN1(\ab[9][0] ), .IN2(\CARRYB[8][0] ), .QN(n1961) );
  XOR3X1 U627 ( .IN1(\CARRYB[5][30] ), .IN2(\ab[5][31] ), .IN3(\ab[6][30] ), 
        .Q(\SUMB[6][30] ) );
  NAND2X0 U628 ( .IN1(\CARRYB[5][30] ), .IN2(\ab[6][30] ), .QN(n70) );
  NAND2X0 U629 ( .IN1(\CARRYB[5][30] ), .IN2(\ab[5][31] ), .QN(n71) );
  NAND2X0 U630 ( .IN1(\ab[6][30] ), .IN2(\ab[5][31] ), .QN(n72) );
  NAND3X1 U631 ( .IN1(n70), .IN2(n71), .IN3(n72), .QN(\CARRYB[6][30] ) );
  XOR3X1 U632 ( .IN1(\SUMB[26][26] ), .IN2(\ab[27][25] ), .IN3(
        \CARRYB[26][25] ), .Q(\SUMB[27][25] ) );
  NAND2X1 U633 ( .IN1(\SUMB[26][26] ), .IN2(\CARRYB[26][25] ), .QN(n73) );
  NAND2X0 U634 ( .IN1(\SUMB[26][26] ), .IN2(\ab[27][25] ), .QN(n74) );
  NAND2X1 U635 ( .IN1(\CARRYB[26][25] ), .IN2(\ab[27][25] ), .QN(n75) );
  NAND3X0 U636 ( .IN1(n73), .IN2(n74), .IN3(n75), .QN(\CARRYB[27][25] ) );
  NAND3X0 U637 ( .IN1(n1464), .IN2(n1465), .IN3(n1466), .QN(\CARRYB[26][25] )
         );
  XOR3X1 U638 ( .IN1(\ab[7][4] ), .IN2(\CARRYB[6][4] ), .IN3(\SUMB[6][5] ), 
        .Q(\SUMB[7][4] ) );
  NAND2X1 U639 ( .IN1(\ab[7][4] ), .IN2(\CARRYB[6][4] ), .QN(n76) );
  NAND2X1 U640 ( .IN1(\ab[7][4] ), .IN2(\SUMB[6][5] ), .QN(n77) );
  NAND2X1 U641 ( .IN1(\CARRYB[6][4] ), .IN2(\SUMB[6][5] ), .QN(n78) );
  NAND3X0 U642 ( .IN1(n76), .IN2(n77), .IN3(n78), .QN(\CARRYB[7][4] ) );
  XOR2X1 U643 ( .IN1(\ab[8][4] ), .IN2(\SUMB[7][5] ), .Q(n79) );
  XOR2X1 U644 ( .IN1(n79), .IN2(\CARRYB[7][4] ), .Q(\SUMB[8][4] ) );
  NAND2X1 U645 ( .IN1(\ab[8][4] ), .IN2(\SUMB[7][5] ), .QN(n80) );
  NAND2X0 U646 ( .IN1(\ab[8][4] ), .IN2(\CARRYB[7][4] ), .QN(n81) );
  NAND2X0 U647 ( .IN1(\SUMB[7][5] ), .IN2(\CARRYB[7][4] ), .QN(n82) );
  NAND3X0 U648 ( .IN1(n80), .IN2(n81), .IN3(n82), .QN(\CARRYB[8][4] ) );
  XOR3X1 U649 ( .IN1(\SUMB[1][8] ), .IN2(\ab[2][7] ), .IN3(n1763), .Q(
        \SUMB[2][7] ) );
  NAND2X0 U650 ( .IN1(\SUMB[1][8] ), .IN2(n1763), .QN(n83) );
  NAND2X0 U651 ( .IN1(\SUMB[1][8] ), .IN2(\ab[2][7] ), .QN(n84) );
  NAND2X0 U652 ( .IN1(n1763), .IN2(\ab[2][7] ), .QN(n85) );
  NAND3X1 U653 ( .IN1(n83), .IN2(n84), .IN3(n85), .QN(\CARRYB[2][7] ) );
  XOR3X1 U654 ( .IN1(\CARRYB[9][4] ), .IN2(\ab[10][4] ), .IN3(\SUMB[9][5] ), 
        .Q(\SUMB[10][4] ) );
  NAND2X1 U655 ( .IN1(\CARRYB[9][4] ), .IN2(\SUMB[9][5] ), .QN(n86) );
  NAND2X1 U656 ( .IN1(\CARRYB[9][4] ), .IN2(\ab[10][4] ), .QN(n87) );
  NAND2X1 U657 ( .IN1(\SUMB[9][5] ), .IN2(\ab[10][4] ), .QN(n88) );
  NAND3X0 U658 ( .IN1(n86), .IN2(n87), .IN3(n88), .QN(\CARRYB[10][4] ) );
  AND2X1 U659 ( .IN1(\ab[1][7] ), .IN2(\ab[0][8] ), .Q(n1763) );
  XOR2X1 U660 ( .IN1(n1922), .IN2(\CARRYB[8][5] ), .Q(\SUMB[9][5] ) );
  XOR2X1 U661 ( .IN1(\ab[8][20] ), .IN2(\CARRYB[7][20] ), .Q(n89) );
  XOR2X1 U662 ( .IN1(n89), .IN2(\SUMB[7][21] ), .Q(\SUMB[8][20] ) );
  NAND2X0 U663 ( .IN1(\ab[7][21] ), .IN2(\CARRYB[6][21] ), .QN(n90) );
  NAND2X0 U664 ( .IN1(\ab[7][21] ), .IN2(\SUMB[6][22] ), .QN(n91) );
  NAND2X0 U665 ( .IN1(\CARRYB[6][21] ), .IN2(\SUMB[6][22] ), .QN(n92) );
  NAND3X1 U666 ( .IN1(n90), .IN2(n91), .IN3(n92), .QN(\CARRYB[7][21] ) );
  NAND2X0 U667 ( .IN1(\ab[8][20] ), .IN2(\CARRYB[7][20] ), .QN(n93) );
  NAND2X0 U668 ( .IN1(\ab[8][20] ), .IN2(\SUMB[7][21] ), .QN(n94) );
  NAND2X0 U669 ( .IN1(\CARRYB[7][20] ), .IN2(\SUMB[7][21] ), .QN(n95) );
  NAND3X1 U670 ( .IN1(n93), .IN2(n94), .IN3(n95), .QN(\CARRYB[8][20] ) );
  XOR3X1 U671 ( .IN1(\ab[6][24] ), .IN2(\CARRYB[5][24] ), .IN3(\SUMB[5][25] ), 
        .Q(\SUMB[6][24] ) );
  NAND2X0 U672 ( .IN1(\ab[6][24] ), .IN2(\CARRYB[5][24] ), .QN(n96) );
  NAND2X0 U673 ( .IN1(\ab[6][24] ), .IN2(\SUMB[5][25] ), .QN(n97) );
  NAND2X0 U674 ( .IN1(\CARRYB[5][24] ), .IN2(\SUMB[5][25] ), .QN(n98) );
  NAND3X1 U675 ( .IN1(n96), .IN2(n97), .IN3(n98), .QN(\CARRYB[6][24] ) );
  XOR2X1 U676 ( .IN1(\ab[7][24] ), .IN2(\SUMB[6][25] ), .Q(n99) );
  NAND2X0 U677 ( .IN1(\ab[7][24] ), .IN2(\SUMB[6][25] ), .QN(n100) );
  NAND2X0 U678 ( .IN1(\ab[7][24] ), .IN2(\CARRYB[6][24] ), .QN(n101) );
  NAND2X0 U679 ( .IN1(\SUMB[6][25] ), .IN2(\CARRYB[6][24] ), .QN(n102) );
  DELLN1X2 U680 ( .INP(n2216), .Z(n2115) );
  XOR3X1 U681 ( .IN1(\ab[6][5] ), .IN2(\CARRYB[5][5] ), .IN3(\SUMB[5][6] ), 
        .Q(\SUMB[6][5] ) );
  NAND2X1 U682 ( .IN1(\ab[6][5] ), .IN2(\CARRYB[5][5] ), .QN(n103) );
  NAND2X0 U683 ( .IN1(\ab[6][5] ), .IN2(\SUMB[5][6] ), .QN(n104) );
  NAND2X0 U684 ( .IN1(\CARRYB[5][5] ), .IN2(\SUMB[5][6] ), .QN(n105) );
  XOR2X1 U685 ( .IN1(\ab[7][5] ), .IN2(\SUMB[6][6] ), .Q(n106) );
  NAND2X0 U686 ( .IN1(\ab[7][5] ), .IN2(\SUMB[6][6] ), .QN(n107) );
  NAND2X0 U687 ( .IN1(\ab[7][5] ), .IN2(\CARRYB[6][5] ), .QN(n108) );
  NAND2X0 U688 ( .IN1(\SUMB[6][6] ), .IN2(\CARRYB[6][5] ), .QN(n109) );
  NAND3X1 U689 ( .IN1(n107), .IN2(n108), .IN3(n109), .QN(\CARRYB[7][5] ) );
  XOR2X1 U690 ( .IN1(n740), .IN2(\SUMB[12][5] ), .Q(\SUMB[13][4] ) );
  XNOR2X2 U691 ( .IN1(n110), .IN2(\SUMB[23][22] ), .Q(\SUMB[24][21] ) );
  XNOR2X1 U692 ( .IN1(\ab[24][21] ), .IN2(\CARRYB[23][21] ), .Q(n110) );
  NAND2X0 U693 ( .IN1(\ab[18][4] ), .IN2(\CARRYB[17][4] ), .QN(n1125) );
  XOR3X1 U694 ( .IN1(\ab[6][25] ), .IN2(\CARRYB[5][25] ), .IN3(\SUMB[5][26] ), 
        .Q(\SUMB[6][25] ) );
  NAND2X0 U695 ( .IN1(\ab[6][25] ), .IN2(\CARRYB[5][25] ), .QN(n111) );
  NAND2X0 U696 ( .IN1(\ab[6][25] ), .IN2(\SUMB[5][26] ), .QN(n112) );
  NAND2X0 U697 ( .IN1(\CARRYB[5][25] ), .IN2(\SUMB[5][26] ), .QN(n113) );
  NAND3X1 U698 ( .IN1(n111), .IN2(n112), .IN3(n113), .QN(\CARRYB[6][25] ) );
  XOR2X1 U699 ( .IN1(n114), .IN2(\CARRYB[6][25] ), .Q(\SUMB[7][25] ) );
  NAND2X0 U700 ( .IN1(\ab[7][25] ), .IN2(\SUMB[6][26] ), .QN(n115) );
  NAND2X0 U701 ( .IN1(\ab[7][25] ), .IN2(\CARRYB[6][25] ), .QN(n116) );
  NAND2X0 U702 ( .IN1(\SUMB[6][26] ), .IN2(\CARRYB[6][25] ), .QN(n117) );
  XOR3X1 U703 ( .IN1(\ab[14][9] ), .IN2(\CARRYB[13][9] ), .IN3(\SUMB[13][10] ), 
        .Q(\SUMB[14][9] ) );
  NAND2X0 U704 ( .IN1(\ab[14][9] ), .IN2(\CARRYB[13][9] ), .QN(n118) );
  NAND2X0 U705 ( .IN1(\ab[14][9] ), .IN2(\SUMB[13][10] ), .QN(n119) );
  NAND2X0 U706 ( .IN1(\CARRYB[13][9] ), .IN2(\SUMB[13][10] ), .QN(n120) );
  NAND2X0 U707 ( .IN1(\ab[15][8] ), .IN2(\CARRYB[14][8] ), .QN(n121) );
  NAND2X0 U708 ( .IN1(\ab[15][8] ), .IN2(\SUMB[14][9] ), .QN(n122) );
  NAND2X0 U709 ( .IN1(\CARRYB[14][8] ), .IN2(\SUMB[14][9] ), .QN(n123) );
  XOR3X1 U710 ( .IN1(\CARRYB[12][9] ), .IN2(\ab[13][9] ), .IN3(\SUMB[12][10] ), 
        .Q(\SUMB[13][9] ) );
  NAND2X0 U711 ( .IN1(\CARRYB[12][9] ), .IN2(\SUMB[12][10] ), .QN(n124) );
  NAND2X0 U712 ( .IN1(\CARRYB[12][9] ), .IN2(\ab[13][9] ), .QN(n125) );
  NAND2X0 U713 ( .IN1(\SUMB[12][10] ), .IN2(\ab[13][9] ), .QN(n126) );
  NAND3X0 U714 ( .IN1(n124), .IN2(n125), .IN3(n126), .QN(\CARRYB[13][9] ) );
  NAND3X0 U715 ( .IN1(n1301), .IN2(n1302), .IN3(n1303), .QN(\CARRYB[12][9] )
         );
  NAND2X0 U716 ( .IN1(\ab[7][13] ), .IN2(\SUMB[6][14] ), .QN(n1735) );
  XOR2X1 U717 ( .IN1(\ab[9][1] ), .IN2(\SUMB[8][2] ), .Q(n127) );
  XOR2X1 U718 ( .IN1(n127), .IN2(\CARRYB[8][1] ), .Q(\SUMB[9][1] ) );
  NAND2X0 U719 ( .IN1(\CARRYB[8][1] ), .IN2(\SUMB[8][2] ), .QN(n128) );
  NAND2X0 U720 ( .IN1(\CARRYB[8][1] ), .IN2(\ab[9][1] ), .QN(n129) );
  NAND2X1 U721 ( .IN1(\SUMB[8][2] ), .IN2(\ab[9][1] ), .QN(n130) );
  XOR3X1 U722 ( .IN1(\ab[26][23] ), .IN2(\CARRYB[25][23] ), .IN3(
        \SUMB[25][24] ), .Q(\SUMB[26][23] ) );
  NAND2X1 U723 ( .IN1(\ab[26][23] ), .IN2(\CARRYB[25][23] ), .QN(n131) );
  NAND2X1 U724 ( .IN1(\ab[26][23] ), .IN2(\SUMB[25][24] ), .QN(n132) );
  NAND2X1 U725 ( .IN1(\CARRYB[25][23] ), .IN2(\SUMB[25][24] ), .QN(n133) );
  XOR2X1 U726 ( .IN1(\ab[27][23] ), .IN2(\SUMB[26][24] ), .Q(n134) );
  XOR2X1 U727 ( .IN1(n134), .IN2(\CARRYB[26][23] ), .Q(\SUMB[27][23] ) );
  NAND2X0 U728 ( .IN1(\ab[27][23] ), .IN2(\SUMB[26][24] ), .QN(n135) );
  NAND2X0 U729 ( .IN1(\ab[27][23] ), .IN2(\CARRYB[26][23] ), .QN(n136) );
  NAND2X0 U730 ( .IN1(\SUMB[26][24] ), .IN2(\CARRYB[26][23] ), .QN(n137) );
  XOR3X1 U731 ( .IN1(\CARRYB[22][26] ), .IN2(\ab[23][26] ), .IN3(
        \SUMB[22][27] ), .Q(\SUMB[23][26] ) );
  NAND2X0 U732 ( .IN1(\CARRYB[22][26] ), .IN2(\SUMB[22][27] ), .QN(n138) );
  NAND2X0 U733 ( .IN1(\CARRYB[22][26] ), .IN2(\ab[23][26] ), .QN(n139) );
  NAND2X0 U734 ( .IN1(\SUMB[22][27] ), .IN2(\ab[23][26] ), .QN(n140) );
  NAND3X0 U735 ( .IN1(n138), .IN2(n139), .IN3(n140), .QN(\CARRYB[23][26] ) );
  XOR3X2 U736 ( .IN1(\ab[4][30] ), .IN2(\ab[3][31] ), .IN3(\CARRYB[3][30] ), 
        .Q(\SUMB[4][30] ) );
  XOR2X1 U737 ( .IN1(\ab[5][29] ), .IN2(\CARRYB[4][29] ), .Q(n141) );
  NAND2X0 U738 ( .IN1(\ab[4][30] ), .IN2(\ab[3][31] ), .QN(n142) );
  NAND2X0 U739 ( .IN1(\ab[4][30] ), .IN2(\CARRYB[3][30] ), .QN(n143) );
  NAND2X0 U740 ( .IN1(\ab[3][31] ), .IN2(\CARRYB[3][30] ), .QN(n144) );
  NAND3X1 U741 ( .IN1(n142), .IN2(n143), .IN3(n144), .QN(\CARRYB[4][30] ) );
  NAND2X0 U742 ( .IN1(\ab[5][29] ), .IN2(\CARRYB[4][29] ), .QN(n145) );
  NAND2X0 U743 ( .IN1(\ab[5][29] ), .IN2(\SUMB[4][30] ), .QN(n146) );
  NAND2X0 U744 ( .IN1(\CARRYB[4][29] ), .IN2(\SUMB[4][30] ), .QN(n147) );
  NAND3X1 U745 ( .IN1(n145), .IN2(n146), .IN3(n147), .QN(\CARRYB[5][29] ) );
  DELLN1X2 U746 ( .INP(ZB), .Z(n148) );
  NAND2X0 U747 ( .IN1(\ab[11][9] ), .IN2(\SUMB[10][10] ), .QN(n1299) );
  XOR3X1 U748 ( .IN1(n1123), .IN2(\ab[2][23] ), .IN3(\SUMB[1][24] ), .Q(
        \SUMB[2][23] ) );
  NAND2X0 U749 ( .IN1(n1123), .IN2(\SUMB[1][24] ), .QN(n149) );
  NAND2X0 U750 ( .IN1(n1123), .IN2(\ab[2][23] ), .QN(n150) );
  NAND2X0 U751 ( .IN1(\SUMB[1][24] ), .IN2(\ab[2][23] ), .QN(n151) );
  NAND3X1 U752 ( .IN1(n149), .IN2(n150), .IN3(n151), .QN(\CARRYB[2][23] ) );
  NAND3X1 U753 ( .IN1(n1395), .IN2(n1396), .IN3(n1397), .QN(\CARRYB[9][28] )
         );
  NAND2X0 U754 ( .IN1(\ab[25][24] ), .IN2(\SUMB[24][25] ), .QN(n1506) );
  XOR2X1 U755 ( .IN1(\ab[1][30] ), .IN2(\ab[0][31] ), .Q(\SUMB[1][30] ) );
  XOR2X1 U756 ( .IN1(\ab[3][21] ), .IN2(\SUMB[2][22] ), .Q(n152) );
  XOR2X1 U757 ( .IN1(n152), .IN2(\CARRYB[2][21] ), .Q(\SUMB[3][21] ) );
  NAND2X0 U758 ( .IN1(\CARRYB[2][21] ), .IN2(\SUMB[2][22] ), .QN(n153) );
  NAND2X0 U759 ( .IN1(\CARRYB[2][21] ), .IN2(\ab[3][21] ), .QN(n154) );
  NAND2X1 U760 ( .IN1(\SUMB[2][22] ), .IN2(\ab[3][21] ), .QN(n155) );
  NAND3X1 U761 ( .IN1(n153), .IN2(n154), .IN3(n155), .QN(\CARRYB[3][21] ) );
  DELLN1X2 U762 ( .INP(n2216), .Z(n2113) );
  XOR3X1 U763 ( .IN1(\ab[7][22] ), .IN2(\CARRYB[6][22] ), .IN3(\SUMB[6][23] ), 
        .Q(\SUMB[7][22] ) );
  NAND2X1 U764 ( .IN1(\ab[7][22] ), .IN2(\CARRYB[6][22] ), .QN(n156) );
  NAND2X0 U765 ( .IN1(\ab[7][22] ), .IN2(\SUMB[6][23] ), .QN(n157) );
  NAND2X0 U766 ( .IN1(\CARRYB[6][22] ), .IN2(\SUMB[6][23] ), .QN(n158) );
  NAND3X1 U767 ( .IN1(n156), .IN2(n157), .IN3(n158), .QN(\CARRYB[7][22] ) );
  NAND2X0 U768 ( .IN1(\ab[8][21] ), .IN2(\CARRYB[7][21] ), .QN(n159) );
  NAND2X0 U769 ( .IN1(\ab[8][21] ), .IN2(\SUMB[7][22] ), .QN(n160) );
  NAND2X0 U770 ( .IN1(\CARRYB[7][21] ), .IN2(\SUMB[7][22] ), .QN(n161) );
  XOR3X1 U771 ( .IN1(\SUMB[5][24] ), .IN2(\ab[6][23] ), .IN3(\CARRYB[5][23] ), 
        .Q(\SUMB[6][23] ) );
  NAND2X0 U772 ( .IN1(\CARRYB[5][23] ), .IN2(\SUMB[5][24] ), .QN(n162) );
  NAND2X0 U773 ( .IN1(\ab[6][23] ), .IN2(\SUMB[5][24] ), .QN(n163) );
  NAND2X1 U774 ( .IN1(\CARRYB[5][23] ), .IN2(\ab[6][23] ), .QN(n164) );
  NAND3X0 U775 ( .IN1(n1522), .IN2(n1523), .IN3(n1524), .QN(\CARRYB[5][23] )
         );
  DELLN1X2 U776 ( .INP(n2218), .Z(n2120) );
  AND2X1 U777 ( .IN1(\ab[0][22] ), .IN2(\ab[1][21] ), .Q(n1581) );
  XOR3X1 U778 ( .IN1(\CARRYB[2][20] ), .IN2(\ab[3][20] ), .IN3(\SUMB[2][21] ), 
        .Q(\SUMB[3][20] ) );
  NAND2X0 U779 ( .IN1(\CARRYB[2][20] ), .IN2(\SUMB[2][21] ), .QN(n166) );
  NAND2X0 U780 ( .IN1(\CARRYB[2][20] ), .IN2(\ab[3][20] ), .QN(n167) );
  NAND2X1 U781 ( .IN1(\SUMB[2][21] ), .IN2(\ab[3][20] ), .QN(n168) );
  NAND3X1 U782 ( .IN1(n166), .IN2(n167), .IN3(n168), .QN(\CARRYB[3][20] ) );
  XOR3X1 U783 ( .IN1(\ab[6][19] ), .IN2(\CARRYB[5][19] ), .IN3(\SUMB[5][20] ), 
        .Q(\SUMB[6][19] ) );
  NAND2X0 U784 ( .IN1(\ab[6][19] ), .IN2(\CARRYB[5][19] ), .QN(n169) );
  NAND2X1 U785 ( .IN1(\ab[6][19] ), .IN2(\SUMB[5][20] ), .QN(n170) );
  NAND2X0 U786 ( .IN1(\CARRYB[5][19] ), .IN2(\SUMB[5][20] ), .QN(n171) );
  NAND3X1 U787 ( .IN1(n169), .IN2(n170), .IN3(n171), .QN(\CARRYB[6][19] ) );
  XOR2X1 U788 ( .IN1(\ab[7][19] ), .IN2(\SUMB[6][20] ), .Q(n172) );
  NAND2X0 U789 ( .IN1(\ab[7][19] ), .IN2(\SUMB[6][20] ), .QN(n173) );
  NAND2X0 U790 ( .IN1(\ab[7][19] ), .IN2(\CARRYB[6][19] ), .QN(n174) );
  NAND2X0 U791 ( .IN1(\SUMB[6][20] ), .IN2(\CARRYB[6][19] ), .QN(n175) );
  NAND3X1 U792 ( .IN1(n173), .IN2(n174), .IN3(n175), .QN(\CARRYB[7][19] ) );
  XOR2X1 U793 ( .IN1(n176), .IN2(\SUMB[30][11] ), .Q(n485) );
  XNOR2X1 U794 ( .IN1(\ab[11][18] ), .IN2(\CARRYB[10][18] ), .Q(n177) );
  NAND2X0 U795 ( .IN1(\CARRYB[12][16] ), .IN2(\ab[13][16] ), .QN(n1526) );
  NAND3X1 U796 ( .IN1(n1188), .IN2(n1189), .IN3(n1190), .QN(\CARRYB[4][21] )
         );
  NAND2X0 U797 ( .IN1(\ab[4][21] ), .IN2(\CARRYB[3][21] ), .QN(n1188) );
  XOR2X2 U798 ( .IN1(n382), .IN2(\SUMB[12][18] ), .Q(\SUMB[13][17] ) );
  NAND3X1 U799 ( .IN1(n875), .IN2(n876), .IN3(n877), .QN(\CARRYB[10][18] ) );
  XOR3X1 U800 ( .IN1(\ab[3][23] ), .IN2(\CARRYB[2][23] ), .IN3(\SUMB[2][24] ), 
        .Q(\SUMB[3][23] ) );
  NAND2X0 U801 ( .IN1(\ab[3][23] ), .IN2(\CARRYB[2][23] ), .QN(n178) );
  NAND2X1 U802 ( .IN1(\ab[3][23] ), .IN2(\SUMB[2][24] ), .QN(n179) );
  NAND2X0 U803 ( .IN1(\CARRYB[2][23] ), .IN2(\SUMB[2][24] ), .QN(n180) );
  XOR2X1 U804 ( .IN1(\ab[4][23] ), .IN2(\SUMB[3][24] ), .Q(n181) );
  XOR2X2 U805 ( .IN1(n181), .IN2(\CARRYB[3][23] ), .Q(\SUMB[4][23] ) );
  NAND2X0 U806 ( .IN1(\ab[4][23] ), .IN2(\SUMB[3][24] ), .QN(n182) );
  NAND2X0 U807 ( .IN1(\ab[4][23] ), .IN2(\CARRYB[3][23] ), .QN(n183) );
  NAND2X0 U808 ( .IN1(\SUMB[3][24] ), .IN2(\CARRYB[3][23] ), .QN(n184) );
  XNOR2X2 U809 ( .IN1(n185), .IN2(\CARRYB[4][21] ), .Q(\SUMB[5][21] ) );
  XNOR2X1 U810 ( .IN1(\ab[5][21] ), .IN2(\SUMB[4][22] ), .Q(n185) );
  XOR2X1 U811 ( .IN1(n478), .IN2(\SUMB[13][18] ), .Q(\SUMB[14][17] ) );
  XOR3X1 U812 ( .IN1(\CARRYB[19][11] ), .IN2(\ab[20][11] ), .IN3(
        \SUMB[19][12] ), .Q(\SUMB[20][11] ) );
  NAND2X0 U813 ( .IN1(\CARRYB[19][11] ), .IN2(\SUMB[19][12] ), .QN(n186) );
  NAND2X0 U814 ( .IN1(\CARRYB[19][11] ), .IN2(\ab[20][11] ), .QN(n187) );
  NAND2X0 U815 ( .IN1(\SUMB[19][12] ), .IN2(\ab[20][11] ), .QN(n188) );
  NAND3X1 U816 ( .IN1(n186), .IN2(n187), .IN3(n188), .QN(\CARRYB[20][11] ) );
  XOR2X1 U817 ( .IN1(\ab[12][14] ), .IN2(\CARRYB[11][14] ), .Q(n189) );
  XOR2X1 U818 ( .IN1(n189), .IN2(\SUMB[11][15] ), .Q(\SUMB[12][14] ) );
  NAND2X0 U819 ( .IN1(\SUMB[11][15] ), .IN2(\CARRYB[11][14] ), .QN(n190) );
  NAND2X0 U820 ( .IN1(\SUMB[11][15] ), .IN2(\ab[12][14] ), .QN(n191) );
  NAND2X0 U821 ( .IN1(\CARRYB[11][14] ), .IN2(\ab[12][14] ), .QN(n192) );
  XOR2X1 U822 ( .IN1(\ab[9][17] ), .IN2(\CARRYB[8][17] ), .Q(n193) );
  XOR2X1 U823 ( .IN1(n193), .IN2(\SUMB[8][18] ), .Q(\SUMB[9][17] ) );
  NAND2X0 U824 ( .IN1(\SUMB[8][18] ), .IN2(\CARRYB[8][17] ), .QN(n194) );
  NAND2X0 U825 ( .IN1(\SUMB[8][18] ), .IN2(\ab[9][17] ), .QN(n195) );
  NAND2X1 U826 ( .IN1(\CARRYB[8][17] ), .IN2(\ab[9][17] ), .QN(n196) );
  NAND3X1 U827 ( .IN1(n194), .IN2(n195), .IN3(n196), .QN(\CARRYB[9][17] ) );
  NAND3X0 U828 ( .IN1(n1553), .IN2(n1554), .IN3(n1555), .QN(\CARRYB[11][14] )
         );
  NAND2X0 U829 ( .IN1(\CARRYB[12][14] ), .IN2(\SUMB[12][15] ), .QN(n1318) );
  NAND2X0 U830 ( .IN1(\CARRYB[12][14] ), .IN2(\ab[13][14] ), .QN(n1319) );
  NAND3X0 U831 ( .IN1(n1241), .IN2(n1242), .IN3(n1243), .QN(\CARRYB[8][17] )
         );
  NAND3X1 U832 ( .IN1(n1954), .IN2(n1955), .IN3(n1956), .QN(n197) );
  XOR3X1 U833 ( .IN1(\ab[14][23] ), .IN2(\CARRYB[13][23] ), .IN3(
        \SUMB[13][24] ), .Q(\SUMB[14][23] ) );
  NAND2X1 U834 ( .IN1(\ab[14][23] ), .IN2(\CARRYB[13][23] ), .QN(n198) );
  NAND2X0 U835 ( .IN1(\ab[14][23] ), .IN2(\SUMB[13][24] ), .QN(n199) );
  NAND2X0 U836 ( .IN1(\CARRYB[13][23] ), .IN2(\SUMB[13][24] ), .QN(n200) );
  XOR2X1 U837 ( .IN1(\ab[15][23] ), .IN2(\SUMB[14][24] ), .Q(n201) );
  NAND2X0 U838 ( .IN1(\ab[15][23] ), .IN2(\SUMB[14][24] ), .QN(n202) );
  NAND2X0 U839 ( .IN1(\ab[15][23] ), .IN2(\CARRYB[14][23] ), .QN(n203) );
  NAND2X0 U840 ( .IN1(\SUMB[14][24] ), .IN2(\CARRYB[14][23] ), .QN(n204) );
  XOR3X1 U841 ( .IN1(\ab[6][26] ), .IN2(\CARRYB[5][26] ), .IN3(\SUMB[5][27] ), 
        .Q(\SUMB[6][26] ) );
  NAND2X0 U842 ( .IN1(\ab[6][26] ), .IN2(\CARRYB[5][26] ), .QN(n205) );
  NAND2X0 U843 ( .IN1(\ab[6][26] ), .IN2(\SUMB[5][27] ), .QN(n206) );
  NAND2X0 U844 ( .IN1(\CARRYB[5][26] ), .IN2(\SUMB[5][27] ), .QN(n207) );
  XOR2X1 U845 ( .IN1(\ab[7][26] ), .IN2(\SUMB[6][27] ), .Q(n208) );
  NAND2X0 U846 ( .IN1(\ab[7][26] ), .IN2(\SUMB[6][27] ), .QN(n209) );
  NAND2X0 U847 ( .IN1(\ab[7][26] ), .IN2(\CARRYB[6][26] ), .QN(n210) );
  NAND2X0 U848 ( .IN1(\SUMB[6][27] ), .IN2(\CARRYB[6][26] ), .QN(n211) );
  XOR3X1 U849 ( .IN1(\ab[3][28] ), .IN2(\CARRYB[2][28] ), .IN3(\SUMB[2][29] ), 
        .Q(\SUMB[3][28] ) );
  NAND2X0 U850 ( .IN1(\ab[3][28] ), .IN2(\CARRYB[2][28] ), .QN(n212) );
  NAND2X0 U851 ( .IN1(\ab[3][28] ), .IN2(\SUMB[2][29] ), .QN(n213) );
  NAND2X0 U852 ( .IN1(\CARRYB[2][28] ), .IN2(\SUMB[2][29] ), .QN(n214) );
  NAND3X1 U853 ( .IN1(n212), .IN2(n213), .IN3(n214), .QN(\CARRYB[3][28] ) );
  XOR2X1 U854 ( .IN1(n215), .IN2(\CARRYB[3][28] ), .Q(\SUMB[4][28] ) );
  NAND2X0 U855 ( .IN1(\ab[4][28] ), .IN2(\SUMB[3][29] ), .QN(n216) );
  NAND2X0 U856 ( .IN1(\ab[4][28] ), .IN2(\CARRYB[3][28] ), .QN(n217) );
  NAND2X0 U857 ( .IN1(\SUMB[3][29] ), .IN2(\CARRYB[3][28] ), .QN(n218) );
  XOR2X1 U858 ( .IN1(\ab[1][20] ), .IN2(\ab[0][21] ), .Q(\SUMB[1][20] ) );
  XOR3X1 U859 ( .IN1(\ab[13][18] ), .IN2(\CARRYB[12][18] ), .IN3(
        \SUMB[12][19] ), .Q(\SUMB[13][18] ) );
  NAND2X0 U860 ( .IN1(\ab[13][18] ), .IN2(\CARRYB[12][18] ), .QN(n479) );
  XNOR2X2 U861 ( .IN1(n219), .IN2(\CARRYB[28][19] ), .Q(\SUMB[29][19] ) );
  XNOR2X1 U862 ( .IN1(\ab[29][19] ), .IN2(\SUMB[28][20] ), .Q(n219) );
  NAND2X0 U863 ( .IN1(\CARRYB[8][27] ), .IN2(\ab[9][27] ), .QN(n1409) );
  INVX0 U864 ( .INP(\ab[15][19] ), .ZN(n421) );
  NAND2X0 U865 ( .IN1(\CARRYB[26][20] ), .IN2(\ab[27][20] ), .QN(n775) );
  XOR2X1 U866 ( .IN1(\ab[28][16] ), .IN2(\CARRYB[27][16] ), .Q(n220) );
  XOR2X1 U867 ( .IN1(n220), .IN2(\SUMB[27][17] ), .Q(\SUMB[28][16] ) );
  NAND2X0 U868 ( .IN1(\SUMB[27][17] ), .IN2(\CARRYB[27][16] ), .QN(n221) );
  NAND2X0 U869 ( .IN1(\SUMB[27][17] ), .IN2(\ab[28][16] ), .QN(n222) );
  NAND2X1 U870 ( .IN1(\CARRYB[27][16] ), .IN2(\ab[28][16] ), .QN(n223) );
  XOR2X1 U871 ( .IN1(\ab[8][26] ), .IN2(\SUMB[7][27] ), .Q(n224) );
  XOR2X1 U872 ( .IN1(n224), .IN2(\CARRYB[7][26] ), .Q(\SUMB[8][26] ) );
  XOR3X1 U873 ( .IN1(\ab[26][18] ), .IN2(\CARRYB[25][18] ), .IN3(
        \SUMB[25][19] ), .Q(\SUMB[26][18] ) );
  XOR2X1 U874 ( .IN1(\ab[27][17] ), .IN2(\CARRYB[26][17] ), .Q(n225) );
  XOR2X2 U875 ( .IN1(n225), .IN2(\SUMB[26][18] ), .Q(\SUMB[27][17] ) );
  NAND2X1 U876 ( .IN1(\ab[26][18] ), .IN2(\CARRYB[25][18] ), .QN(n226) );
  NAND2X0 U877 ( .IN1(\ab[26][18] ), .IN2(\SUMB[25][19] ), .QN(n227) );
  NAND2X0 U878 ( .IN1(\CARRYB[25][18] ), .IN2(\SUMB[25][19] ), .QN(n228) );
  NAND2X0 U879 ( .IN1(\ab[27][17] ), .IN2(\CARRYB[26][17] ), .QN(n229) );
  NAND2X0 U880 ( .IN1(\ab[27][17] ), .IN2(\SUMB[26][18] ), .QN(n230) );
  NAND2X0 U881 ( .IN1(\CARRYB[26][17] ), .IN2(\SUMB[26][18] ), .QN(n231) );
  XOR2X1 U882 ( .IN1(\ab[12][22] ), .IN2(\CARRYB[11][22] ), .Q(n232) );
  NAND2X1 U883 ( .IN1(\ab[11][23] ), .IN2(\CARRYB[10][23] ), .QN(n233) );
  NAND2X0 U884 ( .IN1(\ab[11][23] ), .IN2(\SUMB[10][24] ), .QN(n234) );
  NAND2X0 U885 ( .IN1(\CARRYB[10][23] ), .IN2(\SUMB[10][24] ), .QN(n235) );
  NAND2X0 U886 ( .IN1(\ab[12][22] ), .IN2(\CARRYB[11][22] ), .QN(n236) );
  NAND2X0 U887 ( .IN1(\ab[12][22] ), .IN2(\SUMB[11][23] ), .QN(n237) );
  NAND2X0 U888 ( .IN1(\CARRYB[11][22] ), .IN2(\SUMB[11][23] ), .QN(n238) );
  NAND3X0 U889 ( .IN1(n1672), .IN2(n1673), .IN3(n1674), .QN(\CARRYB[27][16] )
         );
  XOR3X1 U890 ( .IN1(\CARRYB[29][22] ), .IN2(\ab[30][22] ), .IN3(
        \SUMB[29][23] ), .Q(\SUMB[30][22] ) );
  NAND2X0 U891 ( .IN1(\CARRYB[29][22] ), .IN2(\SUMB[29][23] ), .QN(n239) );
  NAND2X0 U892 ( .IN1(\CARRYB[29][22] ), .IN2(\ab[30][22] ), .QN(n240) );
  NAND2X1 U893 ( .IN1(\SUMB[29][23] ), .IN2(\ab[30][22] ), .QN(n241) );
  XOR3X1 U894 ( .IN1(\ab[17][25] ), .IN2(\CARRYB[16][25] ), .IN3(
        \SUMB[16][26] ), .Q(\SUMB[17][25] ) );
  XOR2X1 U895 ( .IN1(\ab[18][24] ), .IN2(\CARRYB[17][24] ), .Q(n242) );
  NAND2X0 U896 ( .IN1(\ab[17][25] ), .IN2(\CARRYB[16][25] ), .QN(n243) );
  NAND2X0 U897 ( .IN1(\ab[17][25] ), .IN2(\SUMB[16][26] ), .QN(n244) );
  NAND2X0 U898 ( .IN1(\CARRYB[16][25] ), .IN2(\SUMB[16][26] ), .QN(n245) );
  NAND2X0 U899 ( .IN1(\ab[18][24] ), .IN2(\CARRYB[17][24] ), .QN(n246) );
  NAND2X0 U900 ( .IN1(\ab[18][24] ), .IN2(\SUMB[17][25] ), .QN(n247) );
  NAND2X0 U901 ( .IN1(\CARRYB[17][24] ), .IN2(\SUMB[17][25] ), .QN(n248) );
  XOR3X1 U902 ( .IN1(\CARRYB[12][25] ), .IN2(\ab[13][25] ), .IN3(
        \SUMB[12][26] ), .Q(\SUMB[13][25] ) );
  NAND2X0 U903 ( .IN1(\CARRYB[12][25] ), .IN2(\ab[13][25] ), .QN(n249) );
  NAND2X0 U904 ( .IN1(\CARRYB[12][25] ), .IN2(\SUMB[12][26] ), .QN(n250) );
  NAND2X0 U905 ( .IN1(\ab[13][25] ), .IN2(\SUMB[12][26] ), .QN(n251) );
  XOR2X1 U906 ( .IN1(\ab[14][25] ), .IN2(\SUMB[13][26] ), .Q(n252) );
  NAND2X0 U907 ( .IN1(\ab[14][25] ), .IN2(\SUMB[13][26] ), .QN(n253) );
  NAND2X0 U908 ( .IN1(\ab[14][25] ), .IN2(\CARRYB[13][25] ), .QN(n254) );
  NAND2X0 U909 ( .IN1(\SUMB[13][26] ), .IN2(\CARRYB[13][25] ), .QN(n255) );
  XOR3X1 U910 ( .IN1(\CARRYB[28][22] ), .IN2(\ab[29][22] ), .IN3(
        \SUMB[28][23] ), .Q(\SUMB[29][22] ) );
  NAND2X0 U911 ( .IN1(\CARRYB[28][22] ), .IN2(\SUMB[28][23] ), .QN(n256) );
  NAND2X0 U912 ( .IN1(\CARRYB[28][22] ), .IN2(\ab[29][22] ), .QN(n257) );
  NAND2X1 U913 ( .IN1(\SUMB[28][23] ), .IN2(\ab[29][22] ), .QN(n258) );
  XOR3X1 U914 ( .IN1(\CARRYB[4][14] ), .IN2(\ab[5][14] ), .IN3(\SUMB[4][15] ), 
        .Q(\SUMB[5][14] ) );
  NAND2X0 U915 ( .IN1(\CARRYB[4][14] ), .IN2(\ab[5][14] ), .QN(n259) );
  NAND2X0 U916 ( .IN1(\CARRYB[4][14] ), .IN2(\SUMB[4][15] ), .QN(n260) );
  NAND2X1 U917 ( .IN1(\ab[5][14] ), .IN2(\SUMB[4][15] ), .QN(n261) );
  NAND3X1 U918 ( .IN1(n259), .IN2(n260), .IN3(n261), .QN(\CARRYB[5][14] ) );
  XOR2X1 U919 ( .IN1(\ab[6][14] ), .IN2(\SUMB[5][15] ), .Q(n262) );
  XOR2X2 U920 ( .IN1(n262), .IN2(\CARRYB[5][14] ), .Q(\SUMB[6][14] ) );
  NAND2X0 U921 ( .IN1(\ab[6][14] ), .IN2(\SUMB[5][15] ), .QN(n263) );
  NAND2X0 U922 ( .IN1(\ab[6][14] ), .IN2(\CARRYB[5][14] ), .QN(n264) );
  NAND2X0 U923 ( .IN1(\SUMB[5][15] ), .IN2(\CARRYB[5][14] ), .QN(n265) );
  NAND3X1 U924 ( .IN1(n263), .IN2(n264), .IN3(n265), .QN(\CARRYB[6][14] ) );
  XOR3X1 U925 ( .IN1(\ab[14][10] ), .IN2(\CARRYB[13][10] ), .IN3(
        \SUMB[13][11] ), .Q(\SUMB[14][10] ) );
  NAND2X1 U926 ( .IN1(\ab[14][10] ), .IN2(\CARRYB[13][10] ), .QN(n266) );
  NAND2X0 U927 ( .IN1(\ab[14][10] ), .IN2(\SUMB[13][11] ), .QN(n267) );
  NAND2X0 U928 ( .IN1(\CARRYB[13][10] ), .IN2(\SUMB[13][11] ), .QN(n268) );
  XOR2X1 U929 ( .IN1(\ab[15][10] ), .IN2(\SUMB[14][11] ), .Q(n269) );
  NAND2X0 U930 ( .IN1(\ab[15][10] ), .IN2(\SUMB[14][11] ), .QN(n270) );
  NAND2X0 U931 ( .IN1(\ab[15][10] ), .IN2(\CARRYB[14][10] ), .QN(n271) );
  NAND2X0 U932 ( .IN1(\SUMB[14][11] ), .IN2(\CARRYB[14][10] ), .QN(n272) );
  XOR3X1 U933 ( .IN1(\ab[16][10] ), .IN2(\CARRYB[15][10] ), .IN3(
        \SUMB[15][11] ), .Q(\SUMB[16][10] ) );
  NAND2X1 U934 ( .IN1(\ab[16][10] ), .IN2(\CARRYB[15][10] ), .QN(n273) );
  NAND2X0 U935 ( .IN1(\ab[16][10] ), .IN2(\SUMB[15][11] ), .QN(n274) );
  NAND2X0 U936 ( .IN1(\CARRYB[15][10] ), .IN2(\SUMB[15][11] ), .QN(n275) );
  XOR2X1 U937 ( .IN1(\ab[17][10] ), .IN2(\SUMB[16][11] ), .Q(n276) );
  NAND2X0 U938 ( .IN1(\ab[17][10] ), .IN2(\SUMB[16][11] ), .QN(n277) );
  NAND2X0 U939 ( .IN1(\ab[17][10] ), .IN2(\CARRYB[16][10] ), .QN(n278) );
  NAND2X0 U940 ( .IN1(\SUMB[16][11] ), .IN2(\CARRYB[16][10] ), .QN(n279) );
  XOR3X1 U941 ( .IN1(\ab[30][4] ), .IN2(\CARRYB[29][4] ), .IN3(\SUMB[29][5] ), 
        .Q(\SUMB[30][4] ) );
  NAND2X0 U942 ( .IN1(\ab[30][4] ), .IN2(\CARRYB[29][4] ), .QN(n280) );
  NAND2X1 U943 ( .IN1(\ab[30][4] ), .IN2(\SUMB[29][5] ), .QN(n281) );
  NAND2X0 U944 ( .IN1(\CARRYB[29][4] ), .IN2(\SUMB[29][5] ), .QN(n282) );
  XOR2X1 U945 ( .IN1(\ab[31][4] ), .IN2(\SUMB[30][5] ), .Q(n283) );
  NAND2X0 U946 ( .IN1(\ab[31][4] ), .IN2(\SUMB[30][5] ), .QN(n284) );
  NAND2X0 U947 ( .IN1(\ab[31][4] ), .IN2(\CARRYB[30][4] ), .QN(n285) );
  NAND2X0 U948 ( .IN1(\SUMB[30][5] ), .IN2(\CARRYB[30][4] ), .QN(n286) );
  XOR3X1 U949 ( .IN1(\ab[26][5] ), .IN2(\CARRYB[25][5] ), .IN3(\SUMB[25][6] ), 
        .Q(\SUMB[26][5] ) );
  NAND2X1 U950 ( .IN1(\ab[26][5] ), .IN2(\CARRYB[25][5] ), .QN(n287) );
  NAND2X0 U951 ( .IN1(\ab[26][5] ), .IN2(\SUMB[25][6] ), .QN(n288) );
  NAND2X0 U952 ( .IN1(\CARRYB[25][5] ), .IN2(\SUMB[25][6] ), .QN(n289) );
  XOR2X1 U953 ( .IN1(\ab[27][5] ), .IN2(\SUMB[26][6] ), .Q(n290) );
  NAND2X0 U954 ( .IN1(\ab[27][5] ), .IN2(\SUMB[26][6] ), .QN(n291) );
  NAND2X0 U955 ( .IN1(\ab[27][5] ), .IN2(\CARRYB[26][5] ), .QN(n292) );
  NAND2X0 U956 ( .IN1(\SUMB[26][6] ), .IN2(\CARRYB[26][5] ), .QN(n293) );
  XOR3X1 U957 ( .IN1(\ab[28][14] ), .IN2(\CARRYB[27][14] ), .IN3(
        \SUMB[27][15] ), .Q(\SUMB[28][14] ) );
  NAND2X0 U958 ( .IN1(\ab[28][14] ), .IN2(\CARRYB[27][14] ), .QN(n295) );
  NAND2X1 U959 ( .IN1(\ab[28][14] ), .IN2(\SUMB[27][15] ), .QN(n296) );
  NAND2X0 U960 ( .IN1(\CARRYB[27][14] ), .IN2(\SUMB[27][15] ), .QN(n297) );
  NAND3X1 U961 ( .IN1(n295), .IN2(n296), .IN3(n297), .QN(\CARRYB[28][14] ) );
  XOR2X1 U962 ( .IN1(\ab[29][14] ), .IN2(\SUMB[28][15] ), .Q(n298) );
  NAND2X0 U963 ( .IN1(\ab[29][14] ), .IN2(\SUMB[28][15] ), .QN(n299) );
  NAND2X0 U964 ( .IN1(\ab[29][14] ), .IN2(\CARRYB[28][14] ), .QN(n300) );
  NAND2X0 U965 ( .IN1(\SUMB[28][15] ), .IN2(\CARRYB[28][14] ), .QN(n301) );
  XOR3X1 U966 ( .IN1(\SUMB[26][15] ), .IN2(\ab[27][14] ), .IN3(
        \CARRYB[26][14] ), .Q(\SUMB[27][14] ) );
  NAND2X0 U967 ( .IN1(\SUMB[26][15] ), .IN2(\CARRYB[26][14] ), .QN(n302) );
  NAND2X0 U968 ( .IN1(\SUMB[26][15] ), .IN2(\ab[27][14] ), .QN(n303) );
  NAND2X0 U969 ( .IN1(\CARRYB[26][14] ), .IN2(\ab[27][14] ), .QN(n304) );
  XOR2X1 U970 ( .IN1(\ab[21][16] ), .IN2(\SUMB[20][17] ), .Q(n305) );
  XOR2X2 U971 ( .IN1(n305), .IN2(\CARRYB[20][16] ), .Q(\SUMB[21][16] ) );
  XOR3X1 U972 ( .IN1(\CARRYB[19][16] ), .IN2(\ab[20][16] ), .IN3(
        \SUMB[19][17] ), .Q(\SUMB[20][16] ) );
  NAND2X0 U973 ( .IN1(\CARRYB[19][16] ), .IN2(\SUMB[19][17] ), .QN(n306) );
  NAND2X0 U974 ( .IN1(\CARRYB[19][16] ), .IN2(\ab[20][16] ), .QN(n307) );
  NAND2X0 U975 ( .IN1(\SUMB[19][17] ), .IN2(\ab[20][16] ), .QN(n308) );
  XOR3X1 U976 ( .IN1(\ab[9][21] ), .IN2(\CARRYB[8][21] ), .IN3(n27), .Q(
        \SUMB[9][21] ) );
  NAND2X0 U977 ( .IN1(\ab[9][21] ), .IN2(\CARRYB[8][21] ), .QN(n309) );
  NAND2X0 U978 ( .IN1(\CARRYB[8][21] ), .IN2(n57), .QN(n311) );
  NAND3X1 U979 ( .IN1(n309), .IN2(n310), .IN3(n311), .QN(\CARRYB[9][21] ) );
  XOR2X1 U980 ( .IN1(\ab[10][21] ), .IN2(\SUMB[9][22] ), .Q(n312) );
  XOR2X2 U981 ( .IN1(n312), .IN2(\CARRYB[9][21] ), .Q(\SUMB[10][21] ) );
  NAND2X0 U982 ( .IN1(\ab[10][21] ), .IN2(\SUMB[9][22] ), .QN(n313) );
  NAND2X0 U983 ( .IN1(\ab[10][21] ), .IN2(\CARRYB[9][21] ), .QN(n314) );
  NAND2X0 U984 ( .IN1(\SUMB[9][22] ), .IN2(\CARRYB[9][21] ), .QN(n315) );
  DELLN1X2 U985 ( .INP(n1971), .Z(n2092) );
  NAND2X0 U986 ( .IN1(\ab[8][25] ), .IN2(\SUMB[7][26] ), .QN(n1447) );
  XNOR2X1 U987 ( .IN1(\ab[13][20] ), .IN2(\SUMB[12][21] ), .Q(n316) );
  XOR3X1 U988 ( .IN1(\ab[26][15] ), .IN2(\CARRYB[25][15] ), .IN3(
        \SUMB[25][16] ), .Q(\SUMB[26][15] ) );
  XOR3X1 U989 ( .IN1(\ab[28][1] ), .IN2(\CARRYB[27][1] ), .IN3(\SUMB[27][2] ), 
        .Q(\SUMB[28][1] ) );
  NAND2X0 U990 ( .IN1(\ab[28][1] ), .IN2(\CARRYB[27][1] ), .QN(n317) );
  NAND2X0 U991 ( .IN1(\ab[28][1] ), .IN2(\SUMB[27][2] ), .QN(n318) );
  NAND2X0 U992 ( .IN1(\CARRYB[27][1] ), .IN2(\SUMB[27][2] ), .QN(n319) );
  NAND3X1 U993 ( .IN1(n317), .IN2(n318), .IN3(n319), .QN(\CARRYB[28][1] ) );
  XOR2X1 U994 ( .IN1(\ab[29][1] ), .IN2(\SUMB[28][2] ), .Q(n320) );
  NAND2X0 U995 ( .IN1(\ab[29][1] ), .IN2(\SUMB[28][2] ), .QN(n321) );
  NAND2X0 U996 ( .IN1(\ab[29][1] ), .IN2(\CARRYB[28][1] ), .QN(n322) );
  NAND2X0 U997 ( .IN1(\SUMB[28][2] ), .IN2(\CARRYB[28][1] ), .QN(n323) );
  NAND3X1 U998 ( .IN1(n321), .IN2(n322), .IN3(n323), .QN(\CARRYB[29][1] ) );
  XOR3X1 U999 ( .IN1(\CARRYB[26][1] ), .IN2(\ab[27][1] ), .IN3(\SUMB[26][2] ), 
        .Q(\SUMB[27][1] ) );
  NAND2X0 U1000 ( .IN1(\CARRYB[26][1] ), .IN2(\SUMB[26][2] ), .QN(n324) );
  NAND2X1 U1001 ( .IN1(\CARRYB[26][1] ), .IN2(\ab[27][1] ), .QN(n325) );
  NAND2X0 U1002 ( .IN1(\SUMB[26][2] ), .IN2(\ab[27][1] ), .QN(n326) );
  XOR2X1 U1003 ( .IN1(\ab[10][7] ), .IN2(\SUMB[9][8] ), .Q(n327) );
  NAND2X0 U1004 ( .IN1(\CARRYB[9][7] ), .IN2(\SUMB[9][8] ), .QN(n328) );
  NAND2X0 U1005 ( .IN1(\CARRYB[9][7] ), .IN2(\ab[10][7] ), .QN(n329) );
  NAND2X0 U1006 ( .IN1(\SUMB[9][8] ), .IN2(\ab[10][7] ), .QN(n330) );
  NAND3X1 U1007 ( .IN1(n328), .IN2(n329), .IN3(n330), .QN(\CARRYB[10][7] ) );
  XOR3X1 U1008 ( .IN1(\CARRYB[20][2] ), .IN2(\ab[21][2] ), .IN3(\SUMB[20][3] ), 
        .Q(\SUMB[21][2] ) );
  NAND2X0 U1009 ( .IN1(\CARRYB[20][2] ), .IN2(\SUMB[20][3] ), .QN(n331) );
  NAND2X0 U1010 ( .IN1(\CARRYB[20][2] ), .IN2(\ab[21][2] ), .QN(n332) );
  NAND2X1 U1011 ( .IN1(\SUMB[20][3] ), .IN2(\ab[21][2] ), .QN(n333) );
  XOR3X1 U1012 ( .IN1(\CARRYB[22][2] ), .IN2(\ab[23][2] ), .IN3(\SUMB[22][3] ), 
        .Q(\SUMB[23][2] ) );
  XOR2X1 U1013 ( .IN1(\ab[23][28] ), .IN2(\SUMB[22][29] ), .Q(n334) );
  XOR2X1 U1014 ( .IN1(n334), .IN2(\CARRYB[22][28] ), .Q(\SUMB[23][28] ) );
  NAND2X0 U1015 ( .IN1(\CARRYB[22][28] ), .IN2(\SUMB[22][29] ), .QN(n335) );
  NAND2X0 U1016 ( .IN1(\CARRYB[22][28] ), .IN2(\ab[23][28] ), .QN(n336) );
  NAND2X0 U1017 ( .IN1(\SUMB[22][29] ), .IN2(\ab[23][28] ), .QN(n337) );
  XOR2X1 U1018 ( .IN1(n338), .IN2(\CARRYB[8][29] ), .Q(\SUMB[9][29] ) );
  NAND2X0 U1019 ( .IN1(\CARRYB[8][29] ), .IN2(\SUMB[8][30] ), .QN(n339) );
  NAND2X0 U1020 ( .IN1(\CARRYB[8][29] ), .IN2(\ab[9][29] ), .QN(n340) );
  NAND2X0 U1021 ( .IN1(\SUMB[8][30] ), .IN2(\ab[9][29] ), .QN(n341) );
  NAND3X1 U1022 ( .IN1(n339), .IN2(n340), .IN3(n341), .QN(\CARRYB[9][29] ) );
  XOR3X1 U1023 ( .IN1(\ab[28][28] ), .IN2(\CARRYB[27][28] ), .IN3(
        \SUMB[27][29] ), .Q(\SUMB[28][28] ) );
  NAND2X0 U1024 ( .IN1(\ab[28][28] ), .IN2(\CARRYB[27][28] ), .QN(n342) );
  NAND2X1 U1025 ( .IN1(\ab[28][28] ), .IN2(\SUMB[27][29] ), .QN(n343) );
  NAND2X0 U1026 ( .IN1(\CARRYB[27][28] ), .IN2(\SUMB[27][29] ), .QN(n344) );
  NAND3X0 U1027 ( .IN1(n342), .IN2(n343), .IN3(n344), .QN(\CARRYB[28][28] ) );
  XOR2X1 U1028 ( .IN1(\ab[29][28] ), .IN2(\SUMB[28][29] ), .Q(n345) );
  XOR2X1 U1029 ( .IN1(n345), .IN2(\CARRYB[28][28] ), .Q(\SUMB[29][28] ) );
  NAND2X1 U1030 ( .IN1(\ab[29][28] ), .IN2(\SUMB[28][29] ), .QN(n346) );
  NAND2X0 U1031 ( .IN1(\ab[29][28] ), .IN2(\CARRYB[28][28] ), .QN(n347) );
  NAND2X0 U1032 ( .IN1(\SUMB[28][29] ), .IN2(\CARRYB[28][28] ), .QN(n348) );
  NAND3X0 U1033 ( .IN1(n346), .IN2(n347), .IN3(n348), .QN(\CARRYB[29][28] ) );
  NAND2X0 U1034 ( .IN1(\SUMB[22][24] ), .IN2(\ab[23][23] ), .QN(n766) );
  XOR2X1 U1035 ( .IN1(n767), .IN2(\SUMB[9][26] ), .Q(\SUMB[10][25] ) );
  NAND2X0 U1036 ( .IN1(\CARRYB[7][26] ), .IN2(\ab[8][26] ), .QN(n781) );
  NAND3X1 U1037 ( .IN1(n967), .IN2(n968), .IN3(n969), .QN(n349) );
  AND2X1 U1038 ( .IN1(\ab[0][31] ), .IN2(\ab[1][30] ), .Q(n422) );
  XOR2X1 U1039 ( .IN1(\ab[1][11] ), .IN2(\ab[0][12] ), .Q(\SUMB[1][11] ) );
  AND2X4 U1040 ( .IN1(n599), .IN2(n546), .Q(\ab[0][30] ) );
  NAND2X0 U1041 ( .IN1(\ab[22][2] ), .IN2(\CARRYB[21][2] ), .QN(n1132) );
  NAND3X1 U1042 ( .IN1(n1138), .IN2(n1139), .IN3(n1140), .QN(\CARRYB[5][7] )
         );
  NAND2X0 U1043 ( .IN1(\SUMB[9][24] ), .IN2(\ab[10][23] ), .QN(n1005) );
  NAND2X0 U1044 ( .IN1(\SUMB[20][21] ), .IN2(\ab[21][20] ), .QN(n573) );
  NAND2X0 U1045 ( .IN1(\ab[24][22] ), .IN2(\SUMB[23][23] ), .QN(n1536) );
  XOR3X1 U1046 ( .IN1(\ab[2][14] ), .IN2(n948), .IN3(\SUMB[1][15] ), .Q(
        \SUMB[2][14] ) );
  NAND2X1 U1047 ( .IN1(\ab[2][14] ), .IN2(n948), .QN(n350) );
  NAND2X0 U1048 ( .IN1(\ab[2][14] ), .IN2(\SUMB[1][15] ), .QN(n351) );
  NAND2X0 U1049 ( .IN1(n948), .IN2(\SUMB[1][15] ), .QN(n352) );
  NAND3X1 U1050 ( .IN1(n350), .IN2(n351), .IN3(n352), .QN(\CARRYB[2][14] ) );
  XOR2X1 U1051 ( .IN1(\ab[3][14] ), .IN2(\SUMB[2][15] ), .Q(n353) );
  NAND2X0 U1052 ( .IN1(\ab[3][14] ), .IN2(\SUMB[2][15] ), .QN(n354) );
  NAND2X0 U1053 ( .IN1(\ab[3][14] ), .IN2(\CARRYB[2][14] ), .QN(n355) );
  NAND2X0 U1054 ( .IN1(\SUMB[2][15] ), .IN2(\CARRYB[2][14] ), .QN(n356) );
  NAND3X1 U1055 ( .IN1(n1298), .IN2(n1299), .IN3(n1300), .QN(\CARRYB[11][9] )
         );
  XOR3X1 U1056 ( .IN1(\ab[15][6] ), .IN2(\CARRYB[14][6] ), .IN3(\SUMB[14][7] ), 
        .Q(\SUMB[15][6] ) );
  NAND2X0 U1057 ( .IN1(\ab[15][6] ), .IN2(\CARRYB[14][6] ), .QN(n357) );
  NAND2X0 U1058 ( .IN1(\ab[15][6] ), .IN2(\SUMB[14][7] ), .QN(n358) );
  NAND2X0 U1059 ( .IN1(\CARRYB[14][6] ), .IN2(\SUMB[14][7] ), .QN(n359) );
  NAND3X1 U1060 ( .IN1(n357), .IN2(n358), .IN3(n359), .QN(\CARRYB[15][6] ) );
  XOR2X1 U1061 ( .IN1(\ab[16][6] ), .IN2(\SUMB[15][7] ), .Q(n360) );
  NAND2X0 U1062 ( .IN1(\ab[16][6] ), .IN2(\SUMB[15][7] ), .QN(n361) );
  NAND2X0 U1063 ( .IN1(\ab[16][6] ), .IN2(\CARRYB[15][6] ), .QN(n362) );
  NAND2X0 U1064 ( .IN1(\SUMB[15][7] ), .IN2(\CARRYB[15][6] ), .QN(n363) );
  NAND3X1 U1065 ( .IN1(n361), .IN2(n362), .IN3(n363), .QN(\CARRYB[16][6] ) );
  XOR3X1 U1066 ( .IN1(\ab[10][9] ), .IN2(\CARRYB[9][9] ), .IN3(\SUMB[9][10] ), 
        .Q(\SUMB[10][9] ) );
  XOR2X1 U1067 ( .IN1(\ab[11][8] ), .IN2(\CARRYB[10][8] ), .Q(n364) );
  XOR2X2 U1068 ( .IN1(n364), .IN2(\SUMB[10][9] ), .Q(\SUMB[11][8] ) );
  NAND2X0 U1069 ( .IN1(\ab[10][9] ), .IN2(\CARRYB[9][9] ), .QN(n365) );
  NAND2X1 U1070 ( .IN1(\ab[10][9] ), .IN2(\SUMB[9][10] ), .QN(n366) );
  NAND2X0 U1071 ( .IN1(\CARRYB[9][9] ), .IN2(\SUMB[9][10] ), .QN(n367) );
  NAND3X1 U1072 ( .IN1(n365), .IN2(n366), .IN3(n367), .QN(\CARRYB[10][9] ) );
  NAND2X0 U1073 ( .IN1(\ab[11][8] ), .IN2(n22), .QN(n368) );
  NAND2X0 U1074 ( .IN1(\ab[11][8] ), .IN2(\SUMB[10][9] ), .QN(n369) );
  NAND2X0 U1075 ( .IN1(n22), .IN2(\SUMB[10][9] ), .QN(n370) );
  NAND3X1 U1076 ( .IN1(n368), .IN2(n369), .IN3(n370), .QN(\CARRYB[11][8] ) );
  XOR2X1 U1077 ( .IN1(\ab[9][9] ), .IN2(\CARRYB[8][9] ), .Q(n371) );
  XOR2X1 U1078 ( .IN1(n371), .IN2(\SUMB[8][10] ), .Q(\SUMB[9][9] ) );
  NAND2X0 U1079 ( .IN1(\SUMB[8][10] ), .IN2(\CARRYB[8][9] ), .QN(n372) );
  NAND2X0 U1080 ( .IN1(\SUMB[8][10] ), .IN2(\ab[9][9] ), .QN(n373) );
  NAND2X0 U1081 ( .IN1(\CARRYB[8][9] ), .IN2(\ab[9][9] ), .QN(n374) );
  NAND3X1 U1082 ( .IN1(n372), .IN2(n373), .IN3(n374), .QN(\CARRYB[9][9] ) );
  XNOR2X2 U1083 ( .IN1(n375), .IN2(\SUMB[6][15] ), .Q(\SUMB[7][14] ) );
  XNOR2X1 U1084 ( .IN1(\ab[7][14] ), .IN2(\CARRYB[6][14] ), .Q(n375) );
  XOR2X1 U1085 ( .IN1(n1644), .IN2(\SUMB[12][11] ), .Q(\SUMB[13][10] ) );
  NAND2X0 U1086 ( .IN1(\CARRYB[10][12] ), .IN2(\ab[11][12] ), .QN(n1322) );
  XOR2X1 U1087 ( .IN1(\ab[10][11] ), .IN2(\CARRYB[9][11] ), .Q(n376) );
  XOR2X1 U1088 ( .IN1(n376), .IN2(\SUMB[9][12] ), .Q(\SUMB[10][11] ) );
  NAND2X0 U1089 ( .IN1(\SUMB[9][12] ), .IN2(\CARRYB[9][11] ), .QN(n377) );
  NAND2X0 U1090 ( .IN1(\SUMB[9][12] ), .IN2(\ab[10][11] ), .QN(n378) );
  NAND2X1 U1091 ( .IN1(\CARRYB[9][11] ), .IN2(\ab[10][11] ), .QN(n379) );
  NAND3X1 U1092 ( .IN1(n377), .IN2(n378), .IN3(n379), .QN(\CARRYB[10][11] ) );
  XNOR2X2 U1093 ( .IN1(n380), .IN2(\CARRYB[11][10] ), .Q(\SUMB[12][10] ) );
  XNOR2X1 U1094 ( .IN1(\ab[12][10] ), .IN2(\SUMB[11][11] ), .Q(n380) );
  XNOR2X1 U1095 ( .IN1(\ab[21][4] ), .IN2(\SUMB[20][5] ), .Q(n381) );
  XOR2X1 U1096 ( .IN1(\ab[13][17] ), .IN2(\CARRYB[12][17] ), .Q(n382) );
  NAND2X0 U1097 ( .IN1(\SUMB[12][18] ), .IN2(\CARRYB[12][17] ), .QN(n383) );
  NAND2X0 U1098 ( .IN1(\SUMB[12][18] ), .IN2(\ab[13][17] ), .QN(n384) );
  NAND2X0 U1099 ( .IN1(\CARRYB[12][17] ), .IN2(\ab[13][17] ), .QN(n385) );
  NAND3X1 U1100 ( .IN1(n383), .IN2(n384), .IN3(n385), .QN(\CARRYB[13][17] ) );
  XOR3X1 U1101 ( .IN1(\ab[2][22] ), .IN2(n716), .IN3(\SUMB[1][23] ), .Q(
        \SUMB[2][22] ) );
  NAND2X0 U1102 ( .IN1(\ab[2][22] ), .IN2(n716), .QN(n386) );
  NAND2X0 U1103 ( .IN1(n716), .IN2(\SUMB[1][23] ), .QN(n388) );
  XOR2X1 U1104 ( .IN1(\ab[3][22] ), .IN2(\SUMB[2][23] ), .Q(n389) );
  XOR2X2 U1105 ( .IN1(n389), .IN2(\CARRYB[2][22] ), .Q(\SUMB[3][22] ) );
  NAND2X0 U1106 ( .IN1(\ab[3][22] ), .IN2(\SUMB[2][23] ), .QN(n390) );
  NAND2X0 U1107 ( .IN1(\ab[3][22] ), .IN2(\CARRYB[2][22] ), .QN(n391) );
  NAND2X0 U1108 ( .IN1(\SUMB[2][23] ), .IN2(\CARRYB[2][22] ), .QN(n392) );
  NAND3X1 U1109 ( .IN1(n391), .IN2(n390), .IN3(n392), .QN(\CARRYB[3][22] ) );
  XNOR2X2 U1110 ( .IN1(n393), .IN2(\SUMB[9][13] ), .Q(\SUMB[10][12] ) );
  XNOR2X1 U1111 ( .IN1(\ab[10][12] ), .IN2(\CARRYB[9][12] ), .Q(n393) );
  XNOR2X2 U1112 ( .IN1(n394), .IN2(\CARRYB[24][3] ), .Q(\SUMB[25][3] ) );
  XOR2X2 U1113 ( .IN1(n1706), .IN2(\CARRYB[17][6] ), .Q(\SUMB[18][6] ) );
  XOR3X1 U1114 ( .IN1(\ab[28][19] ), .IN2(\CARRYB[27][19] ), .IN3(
        \SUMB[27][20] ), .Q(\SUMB[28][19] ) );
  NAND2X0 U1115 ( .IN1(\ab[28][19] ), .IN2(\CARRYB[27][19] ), .QN(n395) );
  NAND2X1 U1116 ( .IN1(\ab[28][19] ), .IN2(\SUMB[27][20] ), .QN(n396) );
  NAND2X0 U1117 ( .IN1(\CARRYB[27][19] ), .IN2(\SUMB[27][20] ), .QN(n397) );
  NAND2X0 U1118 ( .IN1(\ab[29][19] ), .IN2(\SUMB[28][20] ), .QN(n398) );
  NAND2X0 U1119 ( .IN1(\ab[29][19] ), .IN2(\CARRYB[28][19] ), .QN(n399) );
  NAND2X0 U1120 ( .IN1(\SUMB[28][20] ), .IN2(\CARRYB[28][19] ), .QN(n400) );
  NAND3X1 U1121 ( .IN1(n398), .IN2(n399), .IN3(n400), .QN(\CARRYB[29][19] ) );
  XOR3X1 U1122 ( .IN1(n963), .IN2(\ab[2][27] ), .IN3(\SUMB[1][28] ), .Q(
        \SUMB[2][27] ) );
  NAND2X1 U1123 ( .IN1(n963), .IN2(\ab[2][27] ), .QN(n401) );
  NAND2X0 U1124 ( .IN1(n963), .IN2(\SUMB[1][28] ), .QN(n402) );
  NAND2X0 U1125 ( .IN1(\ab[2][27] ), .IN2(\SUMB[1][28] ), .QN(n403) );
  XOR2X1 U1126 ( .IN1(\ab[3][27] ), .IN2(\SUMB[2][28] ), .Q(n404) );
  NAND2X0 U1127 ( .IN1(\ab[3][27] ), .IN2(\SUMB[2][28] ), .QN(n405) );
  NAND2X0 U1128 ( .IN1(\ab[3][27] ), .IN2(\CARRYB[2][27] ), .QN(n406) );
  NAND2X0 U1129 ( .IN1(\SUMB[2][28] ), .IN2(\CARRYB[2][27] ), .QN(n407) );
  NAND3X1 U1130 ( .IN1(n405), .IN2(n406), .IN3(n407), .QN(\CARRYB[3][27] ) );
  XOR3X1 U1131 ( .IN1(\ab[4][27] ), .IN2(\CARRYB[3][27] ), .IN3(\SUMB[3][28] ), 
        .Q(\SUMB[4][27] ) );
  NAND2X1 U1132 ( .IN1(\ab[4][27] ), .IN2(\CARRYB[3][27] ), .QN(n408) );
  NAND2X0 U1133 ( .IN1(\ab[4][27] ), .IN2(\SUMB[3][28] ), .QN(n409) );
  NAND2X0 U1134 ( .IN1(\CARRYB[3][27] ), .IN2(\SUMB[3][28] ), .QN(n410) );
  NAND3X1 U1135 ( .IN1(n408), .IN2(n409), .IN3(n410), .QN(\CARRYB[4][27] ) );
  XOR2X1 U1136 ( .IN1(\ab[5][27] ), .IN2(\SUMB[4][28] ), .Q(n411) );
  NAND2X0 U1137 ( .IN1(\ab[5][27] ), .IN2(\SUMB[4][28] ), .QN(n412) );
  NAND2X0 U1138 ( .IN1(\ab[5][27] ), .IN2(\CARRYB[4][27] ), .QN(n413) );
  NAND2X0 U1139 ( .IN1(\SUMB[4][28] ), .IN2(\CARRYB[4][27] ), .QN(n414) );
  NAND3X1 U1140 ( .IN1(n412), .IN2(n413), .IN3(n414), .QN(\CARRYB[5][27] ) );
  NAND3X1 U1141 ( .IN1(n475), .IN2(n476), .IN3(n477), .QN(\CARRYB[15][16] ) );
  NAND2X0 U1142 ( .IN1(\CARRYB[14][16] ), .IN2(\ab[15][16] ), .QN(n477) );
  XOR3X1 U1143 ( .IN1(\ab[12][20] ), .IN2(\CARRYB[11][20] ), .IN3(
        \SUMB[11][21] ), .Q(\SUMB[12][20] ) );
  NAND2X1 U1144 ( .IN1(\ab[12][20] ), .IN2(\CARRYB[11][20] ), .QN(n415) );
  NAND2X0 U1145 ( .IN1(\ab[12][20] ), .IN2(\SUMB[11][21] ), .QN(n416) );
  NAND2X0 U1146 ( .IN1(\CARRYB[11][20] ), .IN2(\SUMB[11][21] ), .QN(n417) );
  NAND3X1 U1147 ( .IN1(n415), .IN2(n416), .IN3(n417), .QN(\CARRYB[12][20] ) );
  NAND2X0 U1148 ( .IN1(\ab[13][20] ), .IN2(\SUMB[12][21] ), .QN(n418) );
  NAND2X0 U1149 ( .IN1(\ab[13][20] ), .IN2(\CARRYB[12][20] ), .QN(n419) );
  NAND2X0 U1150 ( .IN1(\SUMB[12][21] ), .IN2(\CARRYB[12][20] ), .QN(n420) );
  XNOR3X1 U1151 ( .IN1(n421), .IN2(\CARRYB[14][19] ), .IN3(\SUMB[14][20] ), 
        .Q(\SUMB[15][19] ) );
  NAND2X0 U1152 ( .IN1(\SUMB[10][12] ), .IN2(\ab[11][11] ), .QN(n1653) );
  NAND2X0 U1153 ( .IN1(\SUMB[18][9] ), .IN2(\ab[19][8] ), .QN(n1297) );
  XOR3X1 U1154 ( .IN1(\ab[8][23] ), .IN2(\CARRYB[7][23] ), .IN3(\SUMB[7][24] ), 
        .Q(\SUMB[8][23] ) );
  XOR2X1 U1155 ( .IN1(\ab[9][22] ), .IN2(\CARRYB[8][22] ), .Q(n423) );
  XOR2X2 U1156 ( .IN1(n423), .IN2(\SUMB[8][23] ), .Q(\SUMB[9][22] ) );
  NAND2X1 U1157 ( .IN1(\ab[8][23] ), .IN2(\CARRYB[7][23] ), .QN(n424) );
  NAND2X0 U1158 ( .IN1(\ab[8][23] ), .IN2(\SUMB[7][24] ), .QN(n425) );
  NAND2X0 U1159 ( .IN1(\CARRYB[7][23] ), .IN2(\SUMB[7][24] ), .QN(n426) );
  NAND3X1 U1160 ( .IN1(n424), .IN2(n425), .IN3(n426), .QN(\CARRYB[8][23] ) );
  NAND2X0 U1161 ( .IN1(\ab[9][22] ), .IN2(\CARRYB[8][22] ), .QN(n427) );
  NAND2X0 U1162 ( .IN1(\ab[9][22] ), .IN2(\SUMB[8][23] ), .QN(n428) );
  NAND2X0 U1163 ( .IN1(\CARRYB[8][22] ), .IN2(\SUMB[8][23] ), .QN(n429) );
  NAND3X1 U1164 ( .IN1(n427), .IN2(n428), .IN3(n429), .QN(\CARRYB[9][22] ) );
  XOR3X1 U1165 ( .IN1(\ab[22][21] ), .IN2(\CARRYB[21][21] ), .IN3(
        \SUMB[21][22] ), .Q(\SUMB[22][21] ) );
  XOR2X1 U1166 ( .IN1(\ab[23][20] ), .IN2(\CARRYB[22][20] ), .Q(n430) );
  NAND2X1 U1167 ( .IN1(\ab[22][21] ), .IN2(\CARRYB[21][21] ), .QN(n431) );
  NAND2X0 U1168 ( .IN1(\ab[22][21] ), .IN2(\SUMB[21][22] ), .QN(n432) );
  NAND2X0 U1169 ( .IN1(\CARRYB[21][21] ), .IN2(\SUMB[21][22] ), .QN(n433) );
  NAND3X1 U1170 ( .IN1(n431), .IN2(n432), .IN3(n433), .QN(\CARRYB[22][21] ) );
  NAND2X0 U1171 ( .IN1(\ab[23][20] ), .IN2(\CARRYB[22][20] ), .QN(n434) );
  NAND2X0 U1172 ( .IN1(\ab[23][20] ), .IN2(\SUMB[22][21] ), .QN(n435) );
  NAND2X0 U1173 ( .IN1(\CARRYB[22][20] ), .IN2(\SUMB[22][21] ), .QN(n436) );
  XOR3X1 U1174 ( .IN1(\CARRYB[19][22] ), .IN2(\ab[20][22] ), .IN3(
        \SUMB[19][23] ), .Q(\SUMB[20][22] ) );
  NAND2X0 U1175 ( .IN1(\CARRYB[19][22] ), .IN2(\SUMB[19][23] ), .QN(n437) );
  NAND2X0 U1176 ( .IN1(\CARRYB[19][22] ), .IN2(\ab[20][22] ), .QN(n438) );
  NAND2X1 U1177 ( .IN1(\SUMB[19][23] ), .IN2(\ab[20][22] ), .QN(n439) );
  NAND3X0 U1178 ( .IN1(n437), .IN2(n438), .IN3(n439), .QN(\CARRYB[20][22] ) );
  XOR2X1 U1179 ( .IN1(\ab[14][18] ), .IN2(\CARRYB[13][18] ), .Q(n440) );
  NAND2X1 U1180 ( .IN1(\ab[13][19] ), .IN2(\CARRYB[12][19] ), .QN(n441) );
  NAND2X0 U1181 ( .IN1(\ab[13][19] ), .IN2(\SUMB[12][20] ), .QN(n442) );
  NAND2X0 U1182 ( .IN1(\CARRYB[12][19] ), .IN2(\SUMB[12][20] ), .QN(n443) );
  NAND2X0 U1183 ( .IN1(\ab[14][18] ), .IN2(\CARRYB[13][18] ), .QN(n444) );
  NAND2X0 U1184 ( .IN1(\ab[14][18] ), .IN2(\SUMB[13][19] ), .QN(n445) );
  NAND2X0 U1185 ( .IN1(\CARRYB[13][18] ), .IN2(\SUMB[13][19] ), .QN(n446) );
  XOR2X1 U1186 ( .IN1(\ab[16][17] ), .IN2(\CARRYB[15][17] ), .Q(n447) );
  XOR2X1 U1187 ( .IN1(n447), .IN2(\SUMB[15][18] ), .Q(\SUMB[16][17] ) );
  NAND2X1 U1188 ( .IN1(\ab[15][18] ), .IN2(\CARRYB[14][18] ), .QN(n448) );
  NAND2X0 U1189 ( .IN1(\ab[15][18] ), .IN2(\SUMB[14][19] ), .QN(n449) );
  NAND2X0 U1190 ( .IN1(\CARRYB[14][18] ), .IN2(\SUMB[14][19] ), .QN(n450) );
  NAND3X1 U1191 ( .IN1(n448), .IN2(n449), .IN3(n450), .QN(\CARRYB[15][18] ) );
  NAND2X0 U1192 ( .IN1(\ab[16][17] ), .IN2(\CARRYB[15][17] ), .QN(n451) );
  NAND2X0 U1193 ( .IN1(\ab[16][17] ), .IN2(\SUMB[15][18] ), .QN(n452) );
  NAND2X0 U1194 ( .IN1(\CARRYB[15][17] ), .IN2(\SUMB[15][18] ), .QN(n453) );
  XOR3X1 U1195 ( .IN1(\ab[11][20] ), .IN2(\CARRYB[10][20] ), .IN3(
        \SUMB[10][21] ), .Q(\SUMB[11][20] ) );
  XOR2X1 U1196 ( .IN1(\ab[12][19] ), .IN2(\CARRYB[11][19] ), .Q(n454) );
  XOR2X2 U1197 ( .IN1(n454), .IN2(\SUMB[11][20] ), .Q(\SUMB[12][19] ) );
  NAND2X1 U1198 ( .IN1(\ab[11][20] ), .IN2(\CARRYB[10][20] ), .QN(n455) );
  NAND2X0 U1199 ( .IN1(\ab[11][20] ), .IN2(\SUMB[10][21] ), .QN(n456) );
  NAND2X0 U1200 ( .IN1(\CARRYB[10][20] ), .IN2(\SUMB[10][21] ), .QN(n457) );
  NAND3X1 U1201 ( .IN1(n455), .IN2(n456), .IN3(n457), .QN(\CARRYB[11][20] ) );
  NAND2X0 U1202 ( .IN1(\ab[12][19] ), .IN2(\CARRYB[11][19] ), .QN(n458) );
  NAND2X0 U1203 ( .IN1(\ab[12][19] ), .IN2(\SUMB[11][20] ), .QN(n459) );
  NAND2X0 U1204 ( .IN1(\CARRYB[11][19] ), .IN2(\SUMB[11][20] ), .QN(n460) );
  NAND3X1 U1205 ( .IN1(n458), .IN2(n459), .IN3(n460), .QN(\CARRYB[12][19] ) );
  XOR3X1 U1206 ( .IN1(\ab[18][13] ), .IN2(\CARRYB[17][13] ), .IN3(
        \SUMB[17][14] ), .Q(\SUMB[18][13] ) );
  NAND2X0 U1207 ( .IN1(\ab[18][13] ), .IN2(\SUMB[17][14] ), .QN(n462) );
  NAND2X0 U1208 ( .IN1(\CARRYB[17][13] ), .IN2(\SUMB[17][14] ), .QN(n463) );
  NAND3X1 U1209 ( .IN1(n461), .IN2(n462), .IN3(n463), .QN(\CARRYB[18][13] ) );
  XOR2X1 U1210 ( .IN1(\ab[19][13] ), .IN2(\SUMB[18][14] ), .Q(n464) );
  NAND2X0 U1211 ( .IN1(\ab[19][13] ), .IN2(\SUMB[18][14] ), .QN(n465) );
  NAND2X0 U1212 ( .IN1(\ab[19][13] ), .IN2(\CARRYB[18][13] ), .QN(n466) );
  NAND2X0 U1213 ( .IN1(\SUMB[18][14] ), .IN2(\CARRYB[18][13] ), .QN(n467) );
  XOR3X1 U1214 ( .IN1(\ab[21][11] ), .IN2(\CARRYB[20][11] ), .IN3(
        \SUMB[20][12] ), .Q(\SUMB[21][11] ) );
  NAND2X0 U1215 ( .IN1(\ab[21][11] ), .IN2(\CARRYB[20][11] ), .QN(n468) );
  NAND2X1 U1216 ( .IN1(\ab[21][11] ), .IN2(\SUMB[20][12] ), .QN(n469) );
  NAND2X0 U1217 ( .IN1(\CARRYB[20][11] ), .IN2(\SUMB[20][12] ), .QN(n470) );
  NAND3X1 U1218 ( .IN1(n468), .IN2(n469), .IN3(n470), .QN(\CARRYB[21][11] ) );
  XOR2X1 U1219 ( .IN1(\ab[22][11] ), .IN2(\SUMB[21][12] ), .Q(n471) );
  XOR2X2 U1220 ( .IN1(n471), .IN2(\CARRYB[21][11] ), .Q(\SUMB[22][11] ) );
  NAND2X0 U1221 ( .IN1(\ab[22][11] ), .IN2(\SUMB[21][12] ), .QN(n472) );
  NAND2X0 U1222 ( .IN1(\ab[22][11] ), .IN2(\CARRYB[21][11] ), .QN(n473) );
  NAND2X0 U1223 ( .IN1(\SUMB[21][12] ), .IN2(\CARRYB[21][11] ), .QN(n474) );
  XOR3X1 U1224 ( .IN1(\SUMB[14][17] ), .IN2(\ab[15][16] ), .IN3(
        \CARRYB[14][16] ), .Q(\SUMB[15][16] ) );
  NAND2X0 U1225 ( .IN1(\SUMB[14][17] ), .IN2(\CARRYB[14][16] ), .QN(n475) );
  NAND2X0 U1226 ( .IN1(\SUMB[14][17] ), .IN2(\ab[15][16] ), .QN(n476) );
  XOR2X1 U1227 ( .IN1(\ab[14][17] ), .IN2(\CARRYB[13][17] ), .Q(n478) );
  NAND2X0 U1228 ( .IN1(\ab[13][18] ), .IN2(\SUMB[12][19] ), .QN(n480) );
  NAND2X0 U1229 ( .IN1(\CARRYB[12][18] ), .IN2(\SUMB[12][19] ), .QN(n481) );
  NAND3X1 U1230 ( .IN1(n479), .IN2(n480), .IN3(n481), .QN(\CARRYB[13][18] ) );
  NAND2X0 U1231 ( .IN1(\ab[14][17] ), .IN2(\CARRYB[13][17] ), .QN(n482) );
  NAND2X0 U1232 ( .IN1(\ab[14][17] ), .IN2(\SUMB[13][18] ), .QN(n483) );
  NAND2X0 U1233 ( .IN1(\CARRYB[13][17] ), .IN2(\SUMB[13][18] ), .QN(n484) );
  NAND3X1 U1234 ( .IN1(n482), .IN2(n483), .IN3(n484), .QN(\CARRYB[14][17] ) );
  NAND2X0 U1235 ( .IN1(\SUMB[30][9] ), .IN2(\ab[31][8] ), .QN(n1835) );
  DELLN1X2 U1236 ( .INP(n2205), .Z(n600) );
  DELLN1X2 U1237 ( .INP(n2205), .Z(n601) );
  XNOR2X2 U1238 ( .IN1(n485), .IN2(\CARRYB[30][10] ), .Q(\SUMB[31][10] ) );
  NAND2X0 U1239 ( .IN1(\CARRYB[19][13] ), .IN2(\ab[20][13] ), .QN(n1309) );
  NAND2X0 U1240 ( .IN1(\SUMB[19][14] ), .IN2(\CARRYB[19][13] ), .QN(n1307) );
  XOR3X1 U1241 ( .IN1(\ab[20][10] ), .IN2(\CARRYB[19][10] ), .IN3(
        \SUMB[19][11] ), .Q(\SUMB[20][10] ) );
  XOR2X1 U1242 ( .IN1(\ab[21][9] ), .IN2(\CARRYB[20][9] ), .Q(n486) );
  XOR2X2 U1243 ( .IN1(n486), .IN2(\SUMB[20][10] ), .Q(\SUMB[21][9] ) );
  NAND2X0 U1244 ( .IN1(\ab[20][10] ), .IN2(\CARRYB[19][10] ), .QN(n487) );
  NAND2X0 U1245 ( .IN1(\ab[20][10] ), .IN2(\SUMB[19][11] ), .QN(n488) );
  NAND2X0 U1246 ( .IN1(\CARRYB[19][10] ), .IN2(\SUMB[19][11] ), .QN(n489) );
  NAND3X1 U1247 ( .IN1(n487), .IN2(n488), .IN3(n489), .QN(\CARRYB[20][10] ) );
  NAND2X0 U1248 ( .IN1(\ab[21][9] ), .IN2(\CARRYB[20][9] ), .QN(n490) );
  NAND2X0 U1249 ( .IN1(\ab[21][9] ), .IN2(\SUMB[20][10] ), .QN(n491) );
  NAND2X0 U1250 ( .IN1(\CARRYB[20][9] ), .IN2(\SUMB[20][10] ), .QN(n492) );
  NAND3X1 U1251 ( .IN1(n490), .IN2(n491), .IN3(n492), .QN(\CARRYB[21][9] ) );
  XOR3X1 U1252 ( .IN1(\ab[10][13] ), .IN2(\CARRYB[9][13] ), .IN3(\SUMB[9][14] ), .Q(\SUMB[10][13] ) );
  NAND2X0 U1253 ( .IN1(\ab[10][13] ), .IN2(\CARRYB[9][13] ), .QN(n493) );
  NAND2X0 U1254 ( .IN1(\ab[10][13] ), .IN2(\SUMB[9][14] ), .QN(n494) );
  NAND2X0 U1255 ( .IN1(\CARRYB[9][13] ), .IN2(\SUMB[9][14] ), .QN(n495) );
  NAND3X1 U1256 ( .IN1(n493), .IN2(n494), .IN3(n495), .QN(\CARRYB[10][13] ) );
  XOR2X1 U1257 ( .IN1(\ab[11][13] ), .IN2(\SUMB[10][14] ), .Q(n496) );
  NAND2X0 U1258 ( .IN1(\ab[11][13] ), .IN2(\SUMB[10][14] ), .QN(n497) );
  NAND2X0 U1259 ( .IN1(\ab[11][13] ), .IN2(\CARRYB[10][13] ), .QN(n498) );
  NAND2X0 U1260 ( .IN1(\SUMB[10][14] ), .IN2(\CARRYB[10][13] ), .QN(n499) );
  NAND3X1 U1261 ( .IN1(n497), .IN2(n498), .IN3(n499), .QN(\CARRYB[11][13] ) );
  XOR2X1 U1262 ( .IN1(\ab[19][10] ), .IN2(\SUMB[18][11] ), .Q(n500) );
  XOR2X1 U1263 ( .IN1(n500), .IN2(\CARRYB[18][10] ), .Q(\SUMB[19][10] ) );
  NAND2X0 U1264 ( .IN1(\CARRYB[18][10] ), .IN2(\SUMB[18][11] ), .QN(n501) );
  NAND2X0 U1265 ( .IN1(\CARRYB[18][10] ), .IN2(\ab[19][10] ), .QN(n502) );
  NAND2X0 U1266 ( .IN1(\SUMB[18][11] ), .IN2(\ab[19][10] ), .QN(n503) );
  NAND3X1 U1267 ( .IN1(n501), .IN2(n502), .IN3(n503), .QN(\CARRYB[19][10] ) );
  XOR3X1 U1268 ( .IN1(\ab[28][7] ), .IN2(\CARRYB[27][7] ), .IN3(\SUMB[27][8] ), 
        .Q(\SUMB[28][7] ) );
  NAND2X0 U1269 ( .IN1(\ab[28][7] ), .IN2(\CARRYB[27][7] ), .QN(n504) );
  NAND2X1 U1270 ( .IN1(\ab[28][7] ), .IN2(\SUMB[27][8] ), .QN(n505) );
  NAND2X0 U1271 ( .IN1(\CARRYB[27][7] ), .IN2(\SUMB[27][8] ), .QN(n506) );
  XOR2X1 U1272 ( .IN1(\ab[29][7] ), .IN2(\SUMB[28][8] ), .Q(n507) );
  XOR2X2 U1273 ( .IN1(n507), .IN2(\CARRYB[28][7] ), .Q(\SUMB[29][7] ) );
  NAND2X0 U1274 ( .IN1(\ab[29][7] ), .IN2(\SUMB[28][8] ), .QN(n508) );
  NAND2X0 U1275 ( .IN1(\ab[29][7] ), .IN2(\CARRYB[28][7] ), .QN(n509) );
  NAND2X0 U1276 ( .IN1(\SUMB[28][8] ), .IN2(\CARRYB[28][7] ), .QN(n510) );
  XOR3X1 U1277 ( .IN1(\CARRYB[26][7] ), .IN2(\ab[27][7] ), .IN3(\SUMB[26][8] ), 
        .Q(\SUMB[27][7] ) );
  NAND2X0 U1278 ( .IN1(\CARRYB[26][7] ), .IN2(\SUMB[26][8] ), .QN(n511) );
  NAND2X0 U1279 ( .IN1(\CARRYB[26][7] ), .IN2(\ab[27][7] ), .QN(n512) );
  NAND2X0 U1280 ( .IN1(\SUMB[26][8] ), .IN2(\ab[27][7] ), .QN(n513) );
  XOR2X1 U1281 ( .IN1(n978), .IN2(\CARRYB[17][11] ), .Q(\SUMB[18][11] ) );
  XOR2X1 U1282 ( .IN1(\ab[15][20] ), .IN2(\SUMB[14][21] ), .Q(n514) );
  XOR2X1 U1283 ( .IN1(n514), .IN2(\CARRYB[14][20] ), .Q(\SUMB[15][20] ) );
  NAND2X0 U1284 ( .IN1(\CARRYB[14][20] ), .IN2(\SUMB[14][21] ), .QN(n515) );
  NAND2X0 U1285 ( .IN1(\CARRYB[14][20] ), .IN2(\ab[15][20] ), .QN(n516) );
  NAND2X1 U1286 ( .IN1(\SUMB[14][21] ), .IN2(\ab[15][20] ), .QN(n517) );
  XOR3X1 U1287 ( .IN1(\ab[17][18] ), .IN2(\CARRYB[16][18] ), .IN3(
        \SUMB[16][19] ), .Q(\SUMB[17][18] ) );
  XOR2X1 U1288 ( .IN1(\ab[18][17] ), .IN2(\CARRYB[17][17] ), .Q(n518) );
  NAND2X0 U1289 ( .IN1(\ab[17][18] ), .IN2(\CARRYB[16][18] ), .QN(n519) );
  NAND2X1 U1290 ( .IN1(\ab[17][18] ), .IN2(\SUMB[16][19] ), .QN(n520) );
  NAND2X0 U1291 ( .IN1(\CARRYB[16][18] ), .IN2(\SUMB[16][19] ), .QN(n521) );
  NAND2X0 U1292 ( .IN1(\ab[18][17] ), .IN2(\CARRYB[17][17] ), .QN(n522) );
  NAND2X0 U1293 ( .IN1(\ab[18][17] ), .IN2(\SUMB[17][18] ), .QN(n523) );
  NAND2X0 U1294 ( .IN1(\CARRYB[17][17] ), .IN2(\SUMB[17][18] ), .QN(n524) );
  XOR3X1 U1295 ( .IN1(\CARRYB[2][29] ), .IN2(\ab[3][29] ), .IN3(\SUMB[2][30] ), 
        .Q(\SUMB[3][29] ) );
  NAND2X1 U1296 ( .IN1(\CARRYB[2][29] ), .IN2(\ab[3][29] ), .QN(n525) );
  NAND2X0 U1297 ( .IN1(\CARRYB[2][29] ), .IN2(\SUMB[2][30] ), .QN(n526) );
  NAND2X0 U1298 ( .IN1(\ab[3][29] ), .IN2(\SUMB[2][30] ), .QN(n527) );
  NAND3X1 U1299 ( .IN1(n525), .IN2(n526), .IN3(n527), .QN(\CARRYB[3][29] ) );
  XOR2X1 U1300 ( .IN1(\ab[4][29] ), .IN2(\SUMB[3][30] ), .Q(n528) );
  XOR2X2 U1301 ( .IN1(n528), .IN2(\CARRYB[3][29] ), .Q(\SUMB[4][29] ) );
  NAND2X0 U1302 ( .IN1(\ab[4][29] ), .IN2(\SUMB[3][30] ), .QN(n529) );
  NAND2X0 U1303 ( .IN1(\ab[4][29] ), .IN2(\CARRYB[3][29] ), .QN(n530) );
  NAND2X0 U1304 ( .IN1(\SUMB[3][30] ), .IN2(\CARRYB[3][29] ), .QN(n531) );
  NAND3X1 U1305 ( .IN1(n529), .IN2(n530), .IN3(n531), .QN(\CARRYB[4][29] ) );
  NAND2X0 U1306 ( .IN1(\ab[19][19] ), .IN2(\CARRYB[18][19] ), .QN(n1156) );
  XOR3X1 U1307 ( .IN1(\ab[20][1] ), .IN2(\CARRYB[19][1] ), .IN3(\SUMB[19][2] ), 
        .Q(\SUMB[20][1] ) );
  NAND2X0 U1308 ( .IN1(\ab[20][1] ), .IN2(\SUMB[19][2] ), .QN(n533) );
  NAND2X0 U1309 ( .IN1(\CARRYB[19][1] ), .IN2(\SUMB[19][2] ), .QN(n534) );
  NAND3X1 U1310 ( .IN1(n532), .IN2(n533), .IN3(n534), .QN(\CARRYB[20][1] ) );
  XOR2X1 U1311 ( .IN1(\ab[21][1] ), .IN2(\SUMB[20][2] ), .Q(n535) );
  NAND2X0 U1312 ( .IN1(\ab[21][1] ), .IN2(\SUMB[20][2] ), .QN(n536) );
  NAND2X0 U1313 ( .IN1(\ab[21][1] ), .IN2(\CARRYB[20][1] ), .QN(n537) );
  NAND2X0 U1314 ( .IN1(\SUMB[20][2] ), .IN2(n18), .QN(n538) );
  NAND3X1 U1315 ( .IN1(n536), .IN2(n537), .IN3(n538), .QN(\CARRYB[21][1] ) );
  XOR3X1 U1316 ( .IN1(\ab[3][5] ), .IN2(\CARRYB[2][5] ), .IN3(\SUMB[2][6] ), 
        .Q(\SUMB[3][5] ) );
  NAND2X0 U1317 ( .IN1(\ab[3][5] ), .IN2(\CARRYB[2][5] ), .QN(n539) );
  NAND2X1 U1318 ( .IN1(\ab[3][5] ), .IN2(\SUMB[2][6] ), .QN(n540) );
  NAND2X0 U1319 ( .IN1(\CARRYB[2][5] ), .IN2(\SUMB[2][6] ), .QN(n541) );
  XOR2X1 U1320 ( .IN1(\ab[4][5] ), .IN2(\SUMB[3][6] ), .Q(n542) );
  NAND2X0 U1321 ( .IN1(\ab[4][5] ), .IN2(\SUMB[3][6] ), .QN(n543) );
  NAND2X0 U1322 ( .IN1(\ab[4][5] ), .IN2(\CARRYB[3][5] ), .QN(n544) );
  NAND2X0 U1323 ( .IN1(\SUMB[3][6] ), .IN2(\CARRYB[3][5] ), .QN(n545) );
  XOR3X1 U1324 ( .IN1(\ab[23][0] ), .IN2(\CARRYB[22][0] ), .IN3(\SUMB[22][1] ), 
        .Q(\A1[21] ) );
  NAND2X0 U1325 ( .IN1(\ab[23][0] ), .IN2(\CARRYB[22][0] ), .QN(n547) );
  NAND2X0 U1326 ( .IN1(\ab[23][0] ), .IN2(\SUMB[22][1] ), .QN(n548) );
  NAND2X0 U1327 ( .IN1(\SUMB[22][1] ), .IN2(\CARRYB[22][0] ), .QN(n549) );
  NAND3X1 U1328 ( .IN1(n549), .IN2(n548), .IN3(n547), .QN(\CARRYB[23][0] ) );
  XOR2X1 U1329 ( .IN1(\ab[24][0] ), .IN2(\SUMB[23][1] ), .Q(n550) );
  XOR2X1 U1330 ( .IN1(n550), .IN2(\CARRYB[23][0] ), .Q(\A1[22] ) );
  NAND2X0 U1331 ( .IN1(\ab[24][0] ), .IN2(\SUMB[23][1] ), .QN(n551) );
  NAND2X0 U1332 ( .IN1(\ab[24][0] ), .IN2(\CARRYB[23][0] ), .QN(n552) );
  NAND2X0 U1333 ( .IN1(\SUMB[23][1] ), .IN2(\CARRYB[23][0] ), .QN(n553) );
  NAND3X1 U1334 ( .IN1(n551), .IN2(n552), .IN3(n553), .QN(\CARRYB[24][0] ) );
  XOR3X1 U1335 ( .IN1(\CARRYB[16][0] ), .IN2(\ab[17][0] ), .IN3(\SUMB[16][1] ), 
        .Q(\A1[15] ) );
  NAND2X0 U1336 ( .IN1(\CARRYB[16][0] ), .IN2(\SUMB[16][1] ), .QN(n554) );
  NAND2X0 U1337 ( .IN1(\CARRYB[16][0] ), .IN2(\ab[17][0] ), .QN(n555) );
  NAND2X0 U1338 ( .IN1(\SUMB[16][1] ), .IN2(\ab[17][0] ), .QN(n556) );
  NAND3X1 U1339 ( .IN1(n554), .IN2(n555), .IN3(n556), .QN(\CARRYB[17][0] ) );
  XOR3X1 U1340 ( .IN1(\ab[12][24] ), .IN2(\CARRYB[11][24] ), .IN3(
        \SUMB[11][25] ), .Q(\SUMB[12][24] ) );
  NAND2X0 U1341 ( .IN1(\ab[12][24] ), .IN2(\CARRYB[11][24] ), .QN(n557) );
  NAND2X1 U1342 ( .IN1(\ab[12][24] ), .IN2(\SUMB[11][25] ), .QN(n558) );
  NAND2X0 U1343 ( .IN1(\CARRYB[11][24] ), .IN2(\SUMB[11][25] ), .QN(n559) );
  NAND3X1 U1344 ( .IN1(n557), .IN2(n558), .IN3(n559), .QN(\CARRYB[12][24] ) );
  XOR2X1 U1345 ( .IN1(\ab[13][24] ), .IN2(\SUMB[12][25] ), .Q(n560) );
  NAND2X0 U1346 ( .IN1(\ab[13][24] ), .IN2(\SUMB[12][25] ), .QN(n561) );
  NAND2X0 U1347 ( .IN1(\ab[13][24] ), .IN2(\CARRYB[12][24] ), .QN(n562) );
  NAND2X0 U1348 ( .IN1(\SUMB[12][25] ), .IN2(\CARRYB[12][24] ), .QN(n563) );
  XOR3X1 U1349 ( .IN1(\ab[5][28] ), .IN2(\CARRYB[4][28] ), .IN3(\SUMB[4][29] ), 
        .Q(\SUMB[5][28] ) );
  NAND2X0 U1350 ( .IN1(\ab[5][28] ), .IN2(\CARRYB[4][28] ), .QN(n564) );
  NAND2X1 U1351 ( .IN1(\ab[5][28] ), .IN2(\SUMB[4][29] ), .QN(n565) );
  NAND2X0 U1352 ( .IN1(\CARRYB[4][28] ), .IN2(\SUMB[4][29] ), .QN(n566) );
  XOR2X1 U1353 ( .IN1(\ab[6][28] ), .IN2(\SUMB[5][29] ), .Q(n567) );
  NAND2X0 U1354 ( .IN1(\ab[6][28] ), .IN2(\SUMB[5][29] ), .QN(n568) );
  NAND2X0 U1355 ( .IN1(\ab[6][28] ), .IN2(\CARRYB[5][28] ), .QN(n569) );
  NAND2X0 U1356 ( .IN1(\SUMB[5][29] ), .IN2(\CARRYB[5][28] ), .QN(n570) );
  XOR3X1 U1357 ( .IN1(\CARRYB[20][20] ), .IN2(\ab[21][20] ), .IN3(
        \SUMB[20][21] ), .Q(\SUMB[21][20] ) );
  NAND2X0 U1358 ( .IN1(\CARRYB[20][20] ), .IN2(\SUMB[20][21] ), .QN(n571) );
  NAND2X0 U1359 ( .IN1(\CARRYB[20][20] ), .IN2(\ab[21][20] ), .QN(n572) );
  XOR2X1 U1360 ( .IN1(\ab[20][20] ), .IN2(\CARRYB[19][20] ), .Q(n574) );
  XOR2X1 U1361 ( .IN1(n574), .IN2(\SUMB[19][21] ), .Q(\SUMB[20][20] ) );
  NAND2X0 U1362 ( .IN1(\SUMB[19][21] ), .IN2(\CARRYB[19][20] ), .QN(n575) );
  NAND2X0 U1363 ( .IN1(\SUMB[19][21] ), .IN2(\ab[20][20] ), .QN(n576) );
  NAND2X1 U1364 ( .IN1(\CARRYB[19][20] ), .IN2(\ab[20][20] ), .QN(n577) );
  DELLN1X2 U1365 ( .INP(n2210), .Z(n578) );
  DELLN1X2 U1366 ( .INP(n2210), .Z(n579) );
  DELLN2X2 U1367 ( .INP(n721), .Z(n2090) );
  DELLN1X2 U1368 ( .INP(n2210), .Z(n580) );
  XOR3X1 U1369 ( .IN1(\ab[21][6] ), .IN2(\CARRYB[20][6] ), .IN3(\SUMB[20][7] ), 
        .Q(\SUMB[21][6] ) );
  NAND2X0 U1370 ( .IN1(\ab[21][6] ), .IN2(\CARRYB[20][6] ), .QN(n581) );
  NAND2X1 U1371 ( .IN1(\ab[21][6] ), .IN2(\SUMB[20][7] ), .QN(n582) );
  NAND2X0 U1372 ( .IN1(\CARRYB[20][6] ), .IN2(\SUMB[20][7] ), .QN(n583) );
  XOR2X1 U1373 ( .IN1(\ab[22][6] ), .IN2(\SUMB[21][7] ), .Q(n584) );
  NAND2X0 U1374 ( .IN1(\ab[22][6] ), .IN2(\SUMB[21][7] ), .QN(n585) );
  NAND2X0 U1375 ( .IN1(\ab[22][6] ), .IN2(\CARRYB[21][6] ), .QN(n586) );
  NAND2X0 U1376 ( .IN1(\SUMB[21][7] ), .IN2(\CARRYB[21][6] ), .QN(n587) );
  XOR3X1 U1377 ( .IN1(\CARRYB[16][8] ), .IN2(\ab[17][8] ), .IN3(\SUMB[16][9] ), 
        .Q(\SUMB[17][8] ) );
  NAND2X0 U1378 ( .IN1(\CARRYB[16][8] ), .IN2(\SUMB[16][9] ), .QN(n588) );
  NAND2X1 U1379 ( .IN1(\CARRYB[16][8] ), .IN2(\ab[17][8] ), .QN(n589) );
  NAND2X0 U1380 ( .IN1(\SUMB[16][9] ), .IN2(\ab[17][8] ), .QN(n590) );
  XOR2X1 U1381 ( .IN1(\ab[20][6] ), .IN2(\CARRYB[19][6] ), .Q(n592) );
  NAND2X0 U1382 ( .IN1(\ab[19][7] ), .IN2(\CARRYB[18][7] ), .QN(n593) );
  NAND2X0 U1383 ( .IN1(\ab[19][7] ), .IN2(\SUMB[18][8] ), .QN(n594) );
  NAND2X0 U1384 ( .IN1(\CARRYB[18][7] ), .IN2(\SUMB[18][8] ), .QN(n595) );
  NAND2X0 U1385 ( .IN1(\ab[20][6] ), .IN2(\CARRYB[19][6] ), .QN(n596) );
  NAND2X0 U1386 ( .IN1(\ab[20][6] ), .IN2(\SUMB[19][7] ), .QN(n597) );
  NAND2X0 U1387 ( .IN1(\CARRYB[19][6] ), .IN2(\SUMB[19][7] ), .QN(n598) );
  INVX0 U1388 ( .INP(n1971), .ZN(n599) );
  XOR3X1 U1389 ( .IN1(\ab[23][16] ), .IN2(\CARRYB[22][16] ), .IN3(
        \SUMB[22][17] ), .Q(\SUMB[23][16] ) );
  NAND2X1 U1390 ( .IN1(\ab[23][16] ), .IN2(\CARRYB[22][16] ), .QN(n602) );
  NAND2X0 U1391 ( .IN1(\ab[23][16] ), .IN2(\SUMB[22][17] ), .QN(n603) );
  NAND2X0 U1392 ( .IN1(\CARRYB[22][16] ), .IN2(\SUMB[22][17] ), .QN(n604) );
  XOR2X1 U1393 ( .IN1(\ab[24][16] ), .IN2(\SUMB[23][17] ), .Q(n605) );
  NAND2X0 U1394 ( .IN1(\ab[24][16] ), .IN2(\SUMB[23][17] ), .QN(n606) );
  NAND2X0 U1395 ( .IN1(\ab[24][16] ), .IN2(\CARRYB[23][16] ), .QN(n607) );
  NAND2X0 U1396 ( .IN1(\SUMB[23][17] ), .IN2(\CARRYB[23][16] ), .QN(n608) );
  XOR2X1 U1397 ( .IN1(\ab[19][20] ), .IN2(\CARRYB[18][20] ), .Q(n609) );
  XOR2X1 U1398 ( .IN1(n609), .IN2(\SUMB[18][21] ), .Q(\SUMB[19][20] ) );
  NAND2X0 U1399 ( .IN1(\SUMB[18][21] ), .IN2(\CARRYB[18][20] ), .QN(n610) );
  NAND2X0 U1400 ( .IN1(\SUMB[18][21] ), .IN2(\ab[19][20] ), .QN(n611) );
  NAND2X1 U1401 ( .IN1(\CARRYB[18][20] ), .IN2(\ab[19][20] ), .QN(n612) );
  NAND3X0 U1402 ( .IN1(n610), .IN2(n611), .IN3(n612), .QN(\CARRYB[19][20] ) );
  XOR3X1 U1403 ( .IN1(\ab[9][23] ), .IN2(\CARRYB[8][23] ), .IN3(\SUMB[8][24] ), 
        .Q(\SUMB[9][23] ) );
  XOR2X1 U1404 ( .IN1(\ab[10][22] ), .IN2(\CARRYB[9][22] ), .Q(n613) );
  NAND2X0 U1405 ( .IN1(\ab[9][23] ), .IN2(\CARRYB[8][23] ), .QN(n614) );
  NAND2X0 U1406 ( .IN1(\ab[9][23] ), .IN2(\SUMB[8][24] ), .QN(n615) );
  NAND2X0 U1407 ( .IN1(\CARRYB[8][23] ), .IN2(\SUMB[8][24] ), .QN(n616) );
  NAND2X0 U1408 ( .IN1(\ab[10][22] ), .IN2(\CARRYB[9][22] ), .QN(n617) );
  NAND2X0 U1409 ( .IN1(\ab[10][22] ), .IN2(\SUMB[9][23] ), .QN(n618) );
  NAND2X0 U1410 ( .IN1(\CARRYB[9][22] ), .IN2(\SUMB[9][23] ), .QN(n619) );
  XOR3X1 U1411 ( .IN1(\SUMB[21][18] ), .IN2(\ab[22][17] ), .IN3(
        \CARRYB[21][17] ), .Q(\SUMB[22][17] ) );
  NAND2X0 U1412 ( .IN1(\SUMB[21][18] ), .IN2(\CARRYB[21][17] ), .QN(n620) );
  NAND2X0 U1413 ( .IN1(\SUMB[21][18] ), .IN2(\ab[22][17] ), .QN(n621) );
  NAND2X0 U1414 ( .IN1(\CARRYB[21][17] ), .IN2(\ab[22][17] ), .QN(n622) );
  NAND3X0 U1415 ( .IN1(n707), .IN2(n708), .IN3(n709), .QN(\CARRYB[18][20] ) );
  NAND3X0 U1416 ( .IN1(n1665), .IN2(n1666), .IN3(n1667), .QN(\CARRYB[21][17] )
         );
  XOR2X2 U1417 ( .IN1(n1056), .IN2(\CARRYB[18][18] ), .Q(\SUMB[19][18] ) );
  XNOR2X1 U1418 ( .IN1(\SUMB[20][22] ), .IN2(\ab[21][21] ), .Q(n623) );
  NAND2X0 U1419 ( .IN1(\ab[29][16] ), .IN2(\CARRYB[28][16] ), .QN(n865) );
  XNOR2X1 U1420 ( .IN1(\ab[16][20] ), .IN2(\CARRYB[15][20] ), .Q(n624) );
  NAND2X0 U1421 ( .IN1(\ab[20][3] ), .IN2(\CARRYB[19][3] ), .QN(n625) );
  NAND2X0 U1422 ( .IN1(\ab[20][3] ), .IN2(\SUMB[19][4] ), .QN(n626) );
  NAND2X0 U1423 ( .IN1(\CARRYB[19][3] ), .IN2(\SUMB[19][4] ), .QN(n627) );
  XOR2X1 U1424 ( .IN1(\ab[21][3] ), .IN2(\SUMB[20][4] ), .Q(n628) );
  NAND2X0 U1425 ( .IN1(\ab[21][3] ), .IN2(\SUMB[20][4] ), .QN(n629) );
  NAND2X0 U1426 ( .IN1(\ab[21][3] ), .IN2(\CARRYB[20][3] ), .QN(n630) );
  NAND2X0 U1427 ( .IN1(\SUMB[20][4] ), .IN2(\CARRYB[20][3] ), .QN(n631) );
  XOR3X1 U1428 ( .IN1(\ab[2][10] ), .IN2(n753), .IN3(\SUMB[1][11] ), .Q(
        \SUMB[2][10] ) );
  NAND2X1 U1429 ( .IN1(\ab[2][10] ), .IN2(n753), .QN(n632) );
  NAND2X0 U1430 ( .IN1(\ab[2][10] ), .IN2(\SUMB[1][11] ), .QN(n633) );
  NAND2X0 U1431 ( .IN1(n753), .IN2(\SUMB[1][11] ), .QN(n634) );
  NAND3X1 U1432 ( .IN1(n632), .IN2(n633), .IN3(n634), .QN(\CARRYB[2][10] ) );
  XOR2X1 U1433 ( .IN1(\ab[3][10] ), .IN2(\SUMB[2][11] ), .Q(n635) );
  XOR2X2 U1434 ( .IN1(n635), .IN2(\CARRYB[2][10] ), .Q(\SUMB[3][10] ) );
  NAND2X0 U1435 ( .IN1(\ab[3][10] ), .IN2(\SUMB[2][11] ), .QN(n636) );
  NAND2X0 U1436 ( .IN1(\ab[3][10] ), .IN2(\CARRYB[2][10] ), .QN(n637) );
  NAND2X0 U1437 ( .IN1(\SUMB[2][11] ), .IN2(\CARRYB[2][10] ), .QN(n638) );
  NAND3X1 U1438 ( .IN1(n636), .IN2(n637), .IN3(n638), .QN(\CARRYB[3][10] ) );
  XOR3X1 U1439 ( .IN1(\CARRYB[7][8] ), .IN2(\ab[8][8] ), .IN3(\SUMB[7][9] ), 
        .Q(\SUMB[8][8] ) );
  NAND2X0 U1440 ( .IN1(\CARRYB[7][8] ), .IN2(\ab[8][8] ), .QN(n639) );
  NAND2X0 U1441 ( .IN1(\CARRYB[7][8] ), .IN2(\SUMB[7][9] ), .QN(n640) );
  NAND2X0 U1442 ( .IN1(\ab[8][8] ), .IN2(\SUMB[7][9] ), .QN(n641) );
  XOR2X1 U1443 ( .IN1(\ab[9][8] ), .IN2(\SUMB[8][9] ), .Q(n642) );
  XOR2X2 U1444 ( .IN1(n642), .IN2(\CARRYB[8][8] ), .Q(\SUMB[9][8] ) );
  NAND2X0 U1445 ( .IN1(\ab[9][8] ), .IN2(\SUMB[8][9] ), .QN(n643) );
  NAND2X0 U1446 ( .IN1(\ab[9][8] ), .IN2(\CARRYB[8][8] ), .QN(n644) );
  NAND2X0 U1447 ( .IN1(\SUMB[8][9] ), .IN2(\CARRYB[8][8] ), .QN(n645) );
  DELLN1X2 U1448 ( .INP(n2217), .Z(n2117) );
  XOR3X1 U1449 ( .IN1(\CARRYB[30][22] ), .IN2(\ab[31][22] ), .IN3(
        \SUMB[30][23] ), .Q(\SUMB[31][22] ) );
  NAND2X0 U1450 ( .IN1(\CARRYB[30][22] ), .IN2(\SUMB[30][23] ), .QN(n646) );
  NAND2X0 U1451 ( .IN1(\CARRYB[30][22] ), .IN2(\ab[31][22] ), .QN(n647) );
  NAND2X1 U1452 ( .IN1(\SUMB[30][23] ), .IN2(\ab[31][22] ), .QN(n648) );
  NAND3X0 U1453 ( .IN1(n646), .IN2(n647), .IN3(n648), .QN(\CARRYB[31][22] ) );
  XOR3X1 U1454 ( .IN1(\CARRYB[22][25] ), .IN2(\ab[23][25] ), .IN3(
        \SUMB[22][26] ), .Q(\SUMB[23][25] ) );
  NAND2X0 U1455 ( .IN1(\CARRYB[22][25] ), .IN2(\SUMB[22][26] ), .QN(n649) );
  NAND2X0 U1456 ( .IN1(\CARRYB[22][25] ), .IN2(\ab[23][25] ), .QN(n650) );
  NAND2X0 U1457 ( .IN1(\SUMB[22][26] ), .IN2(\ab[23][25] ), .QN(n651) );
  XOR3X1 U1458 ( .IN1(\CARRYB[17][25] ), .IN2(\ab[18][25] ), .IN3(
        \SUMB[17][26] ), .Q(\SUMB[18][25] ) );
  NAND2X0 U1459 ( .IN1(\CARRYB[17][25] ), .IN2(\SUMB[17][26] ), .QN(n652) );
  NAND2X0 U1460 ( .IN1(\CARRYB[17][25] ), .IN2(\ab[18][25] ), .QN(n653) );
  NAND2X0 U1461 ( .IN1(\SUMB[17][26] ), .IN2(\ab[18][25] ), .QN(n654) );
  XOR2X1 U1462 ( .IN1(\ab[10][28] ), .IN2(\CARRYB[9][28] ), .Q(n655) );
  XOR2X1 U1463 ( .IN1(n655), .IN2(\SUMB[9][29] ), .Q(\SUMB[10][28] ) );
  NAND2X0 U1464 ( .IN1(\SUMB[9][29] ), .IN2(\CARRYB[9][28] ), .QN(n656) );
  NAND2X0 U1465 ( .IN1(\SUMB[9][29] ), .IN2(\ab[10][28] ), .QN(n657) );
  NAND2X0 U1466 ( .IN1(\CARRYB[9][28] ), .IN2(\ab[10][28] ), .QN(n658) );
  XOR3X1 U1467 ( .IN1(\ab[2][2] ), .IN2(n947), .IN3(\SUMB[1][3] ), .Q(
        \SUMB[2][2] ) );
  NAND2X0 U1468 ( .IN1(\ab[2][2] ), .IN2(n947), .QN(n660) );
  NAND2X1 U1469 ( .IN1(\ab[2][2] ), .IN2(\SUMB[1][3] ), .QN(n661) );
  NAND2X0 U1470 ( .IN1(n947), .IN2(\SUMB[1][3] ), .QN(n662) );
  XOR2X1 U1471 ( .IN1(\ab[3][2] ), .IN2(\SUMB[2][3] ), .Q(n663) );
  NAND2X0 U1472 ( .IN1(\ab[3][2] ), .IN2(\SUMB[2][3] ), .QN(n664) );
  NAND2X0 U1473 ( .IN1(\ab[3][2] ), .IN2(\CARRYB[2][2] ), .QN(n665) );
  NAND2X0 U1474 ( .IN1(\SUMB[2][3] ), .IN2(\CARRYB[2][2] ), .QN(n666) );
  XOR3X1 U1475 ( .IN1(\CARRYB[21][5] ), .IN2(\ab[22][5] ), .IN3(\SUMB[21][6] ), 
        .Q(\SUMB[22][5] ) );
  NAND2X1 U1476 ( .IN1(\CARRYB[21][5] ), .IN2(\SUMB[21][6] ), .QN(n667) );
  NAND2X1 U1477 ( .IN1(\CARRYB[21][5] ), .IN2(\ab[22][5] ), .QN(n668) );
  NAND2X0 U1478 ( .IN1(\SUMB[21][6] ), .IN2(\ab[22][5] ), .QN(n669) );
  NAND3X0 U1479 ( .IN1(n667), .IN2(n668), .IN3(n669), .QN(\CARRYB[22][5] ) );
  XOR3X1 U1480 ( .IN1(\ab[24][5] ), .IN2(\CARRYB[23][5] ), .IN3(\SUMB[23][6] ), 
        .Q(\SUMB[24][5] ) );
  NAND2X1 U1481 ( .IN1(\ab[24][5] ), .IN2(\CARRYB[23][5] ), .QN(n670) );
  NAND2X0 U1482 ( .IN1(\ab[24][5] ), .IN2(\SUMB[23][6] ), .QN(n671) );
  NAND2X0 U1483 ( .IN1(\CARRYB[23][5] ), .IN2(\SUMB[23][6] ), .QN(n672) );
  XOR2X1 U1484 ( .IN1(\ab[25][5] ), .IN2(\SUMB[24][6] ), .Q(n673) );
  NAND2X0 U1485 ( .IN1(\ab[25][5] ), .IN2(\SUMB[24][6] ), .QN(n674) );
  NAND2X0 U1486 ( .IN1(\ab[25][5] ), .IN2(\CARRYB[24][5] ), .QN(n675) );
  NAND2X0 U1487 ( .IN1(\SUMB[24][6] ), .IN2(\CARRYB[24][5] ), .QN(n676) );
  XOR3X1 U1488 ( .IN1(\CARRYB[8][6] ), .IN2(\ab[9][6] ), .IN3(\SUMB[8][7] ), 
        .Q(\SUMB[9][6] ) );
  NAND2X1 U1489 ( .IN1(\CARRYB[8][6] ), .IN2(\SUMB[8][7] ), .QN(n677) );
  NAND2X1 U1490 ( .IN1(\CARRYB[8][6] ), .IN2(\ab[9][6] ), .QN(n678) );
  NAND2X0 U1491 ( .IN1(\SUMB[8][7] ), .IN2(\ab[9][6] ), .QN(n679) );
  NAND3X0 U1492 ( .IN1(n677), .IN2(n678), .IN3(n679), .QN(\CARRYB[9][6] ) );
  XOR3X1 U1493 ( .IN1(\ab[10][6] ), .IN2(\CARRYB[9][6] ), .IN3(\SUMB[9][7] ), 
        .Q(\SUMB[10][6] ) );
  NAND2X1 U1494 ( .IN1(\ab[10][6] ), .IN2(\CARRYB[9][6] ), .QN(n680) );
  NAND2X0 U1495 ( .IN1(\ab[10][6] ), .IN2(\SUMB[9][7] ), .QN(n681) );
  NAND2X0 U1496 ( .IN1(\CARRYB[9][6] ), .IN2(\SUMB[9][7] ), .QN(n682) );
  NAND3X1 U1497 ( .IN1(n680), .IN2(n681), .IN3(n682), .QN(\CARRYB[10][6] ) );
  XOR2X1 U1498 ( .IN1(\ab[11][6] ), .IN2(\SUMB[10][7] ), .Q(n683) );
  XOR2X2 U1499 ( .IN1(n683), .IN2(\CARRYB[10][6] ), .Q(\SUMB[11][6] ) );
  NAND2X0 U1500 ( .IN1(\ab[11][6] ), .IN2(\SUMB[10][7] ), .QN(n684) );
  NAND2X0 U1501 ( .IN1(\ab[11][6] ), .IN2(\CARRYB[10][6] ), .QN(n685) );
  NAND2X0 U1502 ( .IN1(\SUMB[10][7] ), .IN2(\CARRYB[10][6] ), .QN(n686) );
  NAND3X1 U1503 ( .IN1(n684), .IN2(n685), .IN3(n686), .QN(\CARRYB[11][6] ) );
  XOR2X1 U1504 ( .IN1(\ab[15][1] ), .IN2(\SUMB[14][2] ), .Q(n1856) );
  XOR3X1 U1505 ( .IN1(\ab[25][21] ), .IN2(\CARRYB[24][21] ), .IN3(
        \SUMB[24][22] ), .Q(\SUMB[25][21] ) );
  NAND2X0 U1506 ( .IN1(\ab[25][21] ), .IN2(\CARRYB[24][21] ), .QN(n688) );
  NAND2X1 U1507 ( .IN1(\ab[25][21] ), .IN2(\SUMB[24][22] ), .QN(n689) );
  NAND2X0 U1508 ( .IN1(\CARRYB[24][21] ), .IN2(\SUMB[24][22] ), .QN(n690) );
  NAND3X1 U1509 ( .IN1(n688), .IN2(n689), .IN3(n690), .QN(\CARRYB[25][21] ) );
  XOR2X1 U1510 ( .IN1(\ab[26][21] ), .IN2(\SUMB[25][22] ), .Q(n691) );
  XOR2X2 U1511 ( .IN1(n691), .IN2(\CARRYB[25][21] ), .Q(\SUMB[26][21] ) );
  NAND2X0 U1512 ( .IN1(\ab[26][21] ), .IN2(\SUMB[25][22] ), .QN(n692) );
  NAND2X0 U1513 ( .IN1(\ab[26][21] ), .IN2(\CARRYB[25][21] ), .QN(n693) );
  NAND2X0 U1514 ( .IN1(\SUMB[25][22] ), .IN2(\CARRYB[25][21] ), .QN(n694) );
  XOR3X1 U1515 ( .IN1(\ab[11][10] ), .IN2(\CARRYB[10][10] ), .IN3(
        \SUMB[10][11] ), .Q(\SUMB[11][10] ) );
  NAND2X0 U1516 ( .IN1(\ab[11][10] ), .IN2(\SUMB[10][11] ), .QN(n696) );
  NAND2X0 U1517 ( .IN1(\CARRYB[10][10] ), .IN2(\SUMB[10][11] ), .QN(n697) );
  NAND2X0 U1518 ( .IN1(\ab[12][10] ), .IN2(n591), .QN(n698) );
  NAND2X0 U1519 ( .IN1(\ab[12][10] ), .IN2(\CARRYB[11][10] ), .QN(n699) );
  NAND2X0 U1520 ( .IN1(\CARRYB[11][10] ), .IN2(n591), .QN(n700) );
  DELLN1X2 U1521 ( .INP(n2225), .Z(n2142) );
  NAND2X0 U1522 ( .IN1(\CARRYB[14][22] ), .IN2(\ab[15][22] ), .QN(n1162) );
  XNOR2X2 U1523 ( .IN1(n701), .IN2(\CARRYB[6][7] ), .Q(\SUMB[7][7] ) );
  XNOR2X1 U1524 ( .IN1(\ab[7][7] ), .IN2(\SUMB[6][8] ), .Q(n701) );
  XNOR2X1 U1525 ( .IN1(\ab[18][8] ), .IN2(\CARRYB[17][8] ), .Q(n702) );
  NAND2X0 U1526 ( .IN1(\ab[6][6] ), .IN2(\CARRYB[5][6] ), .QN(n1347) );
  NAND2X0 U1527 ( .IN1(\ab[17][20] ), .IN2(\SUMB[16][21] ), .QN(n703) );
  NAND2X0 U1528 ( .IN1(\ab[17][20] ), .IN2(\CARRYB[16][20] ), .QN(n704) );
  NAND2X0 U1529 ( .IN1(\SUMB[16][21] ), .IN2(\CARRYB[16][20] ), .QN(n705) );
  XOR2X1 U1530 ( .IN1(n706), .IN2(\CARRYB[17][20] ), .Q(\SUMB[18][20] ) );
  NAND2X0 U1531 ( .IN1(\SUMB[17][21] ), .IN2(\ab[18][20] ), .QN(n707) );
  NAND2X0 U1532 ( .IN1(\SUMB[17][21] ), .IN2(\CARRYB[17][20] ), .QN(n708) );
  NAND2X0 U1533 ( .IN1(\ab[18][20] ), .IN2(\CARRYB[17][20] ), .QN(n709) );
  NAND2X0 U1534 ( .IN1(\ab[15][21] ), .IN2(\CARRYB[14][21] ), .QN(n710) );
  NAND2X0 U1535 ( .IN1(\ab[15][21] ), .IN2(\SUMB[14][22] ), .QN(n711) );
  NAND2X0 U1536 ( .IN1(\CARRYB[14][21] ), .IN2(\SUMB[14][22] ), .QN(n712) );
  NAND2X0 U1537 ( .IN1(\ab[16][20] ), .IN2(\CARRYB[15][20] ), .QN(n713) );
  NAND2X0 U1538 ( .IN1(\ab[16][20] ), .IN2(\SUMB[15][21] ), .QN(n714) );
  NAND2X0 U1539 ( .IN1(\CARRYB[15][20] ), .IN2(\SUMB[15][21] ), .QN(n715) );
  AND2X1 U1540 ( .IN1(\ab[0][23] ), .IN2(\ab[1][22] ), .Q(n716) );
  XOR2X1 U1541 ( .IN1(\ab[1][22] ), .IN2(\ab[0][23] ), .Q(\SUMB[1][22] ) );
  XOR2X1 U1542 ( .IN1(\ab[6][10] ), .IN2(\SUMB[5][11] ), .Q(n717) );
  XOR2X1 U1543 ( .IN1(n717), .IN2(\CARRYB[5][10] ), .Q(\SUMB[6][10] ) );
  NAND2X0 U1544 ( .IN1(\CARRYB[5][10] ), .IN2(\SUMB[5][11] ), .QN(n718) );
  NAND2X0 U1545 ( .IN1(\CARRYB[5][10] ), .IN2(\ab[6][10] ), .QN(n719) );
  NAND2X1 U1546 ( .IN1(\SUMB[5][11] ), .IN2(\ab[6][10] ), .QN(n720) );
  INVX0 U1547 ( .INP(A[1]), .ZN(n721) );
  XOR2X1 U1548 ( .IN1(\ab[5][10] ), .IN2(\SUMB[4][11] ), .Q(n722) );
  XOR2X1 U1549 ( .IN1(n722), .IN2(\CARRYB[4][10] ), .Q(\SUMB[5][10] ) );
  NAND2X0 U1550 ( .IN1(\CARRYB[4][10] ), .IN2(\SUMB[4][11] ), .QN(n723) );
  NAND2X0 U1551 ( .IN1(\CARRYB[4][10] ), .IN2(\ab[5][10] ), .QN(n724) );
  NAND2X1 U1552 ( .IN1(\SUMB[4][11] ), .IN2(\ab[5][10] ), .QN(n725) );
  XOR3X1 U1553 ( .IN1(\ab[4][8] ), .IN2(\CARRYB[3][8] ), .IN3(\SUMB[3][9] ), 
        .Q(\SUMB[4][8] ) );
  NAND2X0 U1554 ( .IN1(\ab[4][8] ), .IN2(\CARRYB[3][8] ), .QN(n726) );
  NAND2X0 U1555 ( .IN1(\ab[4][8] ), .IN2(\SUMB[3][9] ), .QN(n727) );
  NAND2X0 U1556 ( .IN1(\CARRYB[3][8] ), .IN2(\SUMB[3][9] ), .QN(n728) );
  NAND3X1 U1557 ( .IN1(n726), .IN2(n727), .IN3(n728), .QN(\CARRYB[4][8] ) );
  XOR2X1 U1558 ( .IN1(\ab[5][8] ), .IN2(\SUMB[4][9] ), .Q(n729) );
  XOR2X2 U1559 ( .IN1(n729), .IN2(\CARRYB[4][8] ), .Q(\SUMB[5][8] ) );
  NAND2X0 U1560 ( .IN1(\ab[5][8] ), .IN2(\SUMB[4][9] ), .QN(n730) );
  NAND2X0 U1561 ( .IN1(\ab[5][8] ), .IN2(\CARRYB[4][8] ), .QN(n731) );
  NAND2X0 U1562 ( .IN1(\SUMB[4][9] ), .IN2(\CARRYB[4][8] ), .QN(n732) );
  NAND3X1 U1563 ( .IN1(n730), .IN2(n731), .IN3(n732), .QN(\CARRYB[5][8] ) );
  AND2X1 U1564 ( .IN1(\ab[0][10] ), .IN2(\ab[1][9] ), .Q(n1782) );
  XOR3X1 U1565 ( .IN1(\ab[12][3] ), .IN2(\CARRYB[11][3] ), .IN3(\SUMB[11][4] ), 
        .Q(\SUMB[12][3] ) );
  NAND2X0 U1566 ( .IN1(\ab[12][3] ), .IN2(\CARRYB[11][3] ), .QN(n733) );
  NAND2X0 U1567 ( .IN1(\ab[12][3] ), .IN2(\SUMB[11][4] ), .QN(n734) );
  NAND2X0 U1568 ( .IN1(\CARRYB[11][3] ), .IN2(\SUMB[11][4] ), .QN(n735) );
  XOR2X1 U1569 ( .IN1(\ab[13][3] ), .IN2(\SUMB[12][4] ), .Q(n736) );
  NAND2X0 U1570 ( .IN1(\ab[13][3] ), .IN2(\SUMB[12][4] ), .QN(n737) );
  NAND2X0 U1571 ( .IN1(\ab[13][3] ), .IN2(\CARRYB[12][3] ), .QN(n738) );
  NAND2X0 U1572 ( .IN1(\SUMB[12][4] ), .IN2(\CARRYB[12][3] ), .QN(n739) );
  XOR3X1 U1573 ( .IN1(\ab[12][5] ), .IN2(\CARRYB[11][5] ), .IN3(\SUMB[11][6] ), 
        .Q(\SUMB[12][5] ) );
  XOR2X1 U1574 ( .IN1(\ab[13][4] ), .IN2(\CARRYB[12][4] ), .Q(n740) );
  NAND2X0 U1575 ( .IN1(\ab[12][5] ), .IN2(\CARRYB[11][5] ), .QN(n741) );
  NAND2X0 U1576 ( .IN1(\ab[12][5] ), .IN2(\SUMB[11][6] ), .QN(n742) );
  NAND2X0 U1577 ( .IN1(\CARRYB[11][5] ), .IN2(\SUMB[11][6] ), .QN(n743) );
  NAND3X1 U1578 ( .IN1(n741), .IN2(n742), .IN3(n743), .QN(\CARRYB[12][5] ) );
  NAND2X0 U1579 ( .IN1(\ab[13][4] ), .IN2(\CARRYB[12][4] ), .QN(n744) );
  NAND2X0 U1580 ( .IN1(\ab[13][4] ), .IN2(\SUMB[12][5] ), .QN(n745) );
  NAND2X0 U1581 ( .IN1(\CARRYB[12][4] ), .IN2(\SUMB[12][5] ), .QN(n746) );
  NAND3X1 U1582 ( .IN1(n744), .IN2(n745), .IN3(n746), .QN(\CARRYB[13][4] ) );
  XOR3X1 U1583 ( .IN1(\ab[13][5] ), .IN2(\CARRYB[12][5] ), .IN3(\SUMB[12][6] ), 
        .Q(\SUMB[13][5] ) );
  NAND2X0 U1584 ( .IN1(\ab[13][5] ), .IN2(\CARRYB[12][5] ), .QN(n747) );
  NAND2X1 U1585 ( .IN1(\ab[13][5] ), .IN2(\SUMB[12][6] ), .QN(n748) );
  NAND2X0 U1586 ( .IN1(\CARRYB[12][5] ), .IN2(\SUMB[12][6] ), .QN(n749) );
  NAND2X0 U1587 ( .IN1(\ab[14][5] ), .IN2(\SUMB[13][6] ), .QN(n750) );
  NAND2X0 U1588 ( .IN1(\ab[14][5] ), .IN2(\CARRYB[13][5] ), .QN(n751) );
  NAND2X0 U1589 ( .IN1(\SUMB[13][6] ), .IN2(\CARRYB[13][5] ), .QN(n752) );
  AND2X1 U1590 ( .IN1(\ab[0][11] ), .IN2(\ab[1][10] ), .Q(n753) );
  AND2X1 U1591 ( .IN1(\ab[0][6] ), .IN2(\ab[1][5] ), .Q(n754) );
  XNOR2X1 U1592 ( .IN1(\ab[16][2] ), .IN2(\SUMB[15][3] ), .Q(n755) );
  XOR3X1 U1593 ( .IN1(\ab[29][20] ), .IN2(\CARRYB[28][20] ), .IN3(
        \SUMB[28][21] ), .Q(\SUMB[29][20] ) );
  NAND2X1 U1594 ( .IN1(\ab[29][20] ), .IN2(\CARRYB[28][20] ), .QN(n756) );
  NAND2X0 U1595 ( .IN1(\ab[29][20] ), .IN2(\SUMB[28][21] ), .QN(n757) );
  NAND2X0 U1596 ( .IN1(\CARRYB[28][20] ), .IN2(\SUMB[28][21] ), .QN(n758) );
  NAND3X1 U1597 ( .IN1(n756), .IN2(n757), .IN3(n758), .QN(\CARRYB[29][20] ) );
  XOR2X1 U1598 ( .IN1(\ab[30][20] ), .IN2(\SUMB[29][21] ), .Q(n759) );
  NAND2X0 U1599 ( .IN1(\ab[30][20] ), .IN2(\SUMB[29][21] ), .QN(n760) );
  NAND2X0 U1600 ( .IN1(\ab[30][20] ), .IN2(\CARRYB[29][20] ), .QN(n761) );
  NAND2X0 U1601 ( .IN1(\SUMB[29][21] ), .IN2(\CARRYB[29][20] ), .QN(n762) );
  XOR2X1 U1602 ( .IN1(\ab[23][23] ), .IN2(\SUMB[22][24] ), .Q(n763) );
  NAND2X0 U1603 ( .IN1(\CARRYB[22][23] ), .IN2(\SUMB[22][24] ), .QN(n764) );
  NAND2X0 U1604 ( .IN1(\CARRYB[22][23] ), .IN2(\ab[23][23] ), .QN(n765) );
  XOR3X1 U1605 ( .IN1(\CARRYB[8][26] ), .IN2(\ab[9][26] ), .IN3(\SUMB[8][27] ), 
        .Q(\SUMB[9][26] ) );
  XOR2X1 U1606 ( .IN1(\ab[10][25] ), .IN2(\CARRYB[9][25] ), .Q(n767) );
  NAND2X0 U1607 ( .IN1(\ab[9][26] ), .IN2(\CARRYB[8][26] ), .QN(n768) );
  NAND2X0 U1608 ( .IN1(\ab[9][26] ), .IN2(\SUMB[8][27] ), .QN(n769) );
  NAND2X0 U1609 ( .IN1(\CARRYB[8][26] ), .IN2(\SUMB[8][27] ), .QN(n770) );
  NAND2X0 U1610 ( .IN1(\ab[10][25] ), .IN2(\CARRYB[9][25] ), .QN(n771) );
  NAND2X0 U1611 ( .IN1(\ab[10][25] ), .IN2(\SUMB[9][26] ), .QN(n772) );
  NAND2X0 U1612 ( .IN1(\CARRYB[9][25] ), .IN2(\SUMB[9][26] ), .QN(n773) );
  XOR3X1 U1613 ( .IN1(\CARRYB[26][20] ), .IN2(\ab[27][20] ), .IN3(
        \SUMB[26][21] ), .Q(\SUMB[27][20] ) );
  NAND2X0 U1614 ( .IN1(\CARRYB[26][20] ), .IN2(\SUMB[26][21] ), .QN(n774) );
  NAND2X0 U1615 ( .IN1(\SUMB[26][21] ), .IN2(\ab[27][20] ), .QN(n776) );
  XOR3X1 U1616 ( .IN1(\CARRYB[21][23] ), .IN2(\ab[22][23] ), .IN3(
        \SUMB[21][24] ), .Q(\SUMB[22][23] ) );
  NAND2X0 U1617 ( .IN1(\CARRYB[21][23] ), .IN2(\SUMB[21][24] ), .QN(n777) );
  NAND2X0 U1618 ( .IN1(\CARRYB[21][23] ), .IN2(\ab[22][23] ), .QN(n778) );
  NAND2X0 U1619 ( .IN1(\SUMB[21][24] ), .IN2(\ab[22][23] ), .QN(n779) );
  NAND2X0 U1620 ( .IN1(\CARRYB[7][26] ), .IN2(\SUMB[7][27] ), .QN(n780) );
  NAND2X0 U1621 ( .IN1(\SUMB[7][27] ), .IN2(\ab[8][26] ), .QN(n782) );
  XNOR3X1 U1622 ( .IN1(n1027), .IN2(\CARRYB[23][22] ), .IN3(\SUMB[23][23] ), 
        .Q(\SUMB[24][22] ) );
  XOR2X1 U1623 ( .IN1(\ab[1][27] ), .IN2(\ab[0][28] ), .Q(\SUMB[1][27] ) );
  NAND2X0 U1624 ( .IN1(\ab[18][5] ), .IN2(\SUMB[17][6] ), .QN(n1913) );
  XOR3X1 U1625 ( .IN1(\ab[28][15] ), .IN2(\CARRYB[27][15] ), .IN3(
        \SUMB[27][16] ), .Q(\SUMB[28][15] ) );
  NAND2X1 U1626 ( .IN1(\ab[28][15] ), .IN2(\CARRYB[27][15] ), .QN(n783) );
  NAND2X0 U1627 ( .IN1(\ab[28][15] ), .IN2(\SUMB[27][16] ), .QN(n784) );
  NAND2X0 U1628 ( .IN1(\CARRYB[27][15] ), .IN2(\SUMB[27][16] ), .QN(n785) );
  NAND3X1 U1629 ( .IN1(n783), .IN2(n784), .IN3(n785), .QN(\CARRYB[28][15] ) );
  XOR2X1 U1630 ( .IN1(\ab[29][15] ), .IN2(\SUMB[28][16] ), .Q(n786) );
  NAND2X0 U1631 ( .IN1(\ab[29][15] ), .IN2(\SUMB[28][16] ), .QN(n787) );
  NAND2X0 U1632 ( .IN1(\ab[29][15] ), .IN2(\CARRYB[28][15] ), .QN(n788) );
  NAND2X0 U1633 ( .IN1(\SUMB[28][16] ), .IN2(\CARRYB[28][15] ), .QN(n789) );
  XOR3X1 U1634 ( .IN1(\CARRYB[25][17] ), .IN2(\ab[26][17] ), .IN3(
        \SUMB[25][18] ), .Q(\SUMB[26][17] ) );
  NAND2X0 U1635 ( .IN1(\CARRYB[25][17] ), .IN2(\SUMB[25][18] ), .QN(n790) );
  NAND2X1 U1636 ( .IN1(\CARRYB[25][17] ), .IN2(\ab[26][17] ), .QN(n791) );
  NAND2X0 U1637 ( .IN1(\SUMB[25][18] ), .IN2(\ab[26][17] ), .QN(n792) );
  NAND3X0 U1638 ( .IN1(n790), .IN2(n791), .IN3(n792), .QN(\CARRYB[26][17] ) );
  XOR3X1 U1639 ( .IN1(\CARRYB[3][20] ), .IN2(\ab[4][20] ), .IN3(\SUMB[3][21] ), 
        .Q(\SUMB[4][20] ) );
  NAND2X0 U1640 ( .IN1(\CARRYB[3][20] ), .IN2(\SUMB[3][21] ), .QN(n793) );
  NAND2X0 U1641 ( .IN1(\CARRYB[3][20] ), .IN2(\ab[4][20] ), .QN(n794) );
  NAND2X1 U1642 ( .IN1(\SUMB[3][21] ), .IN2(\ab[4][20] ), .QN(n795) );
  NAND3X1 U1643 ( .IN1(n793), .IN2(n794), .IN3(n795), .QN(\CARRYB[4][20] ) );
  XOR3X1 U1644 ( .IN1(\ab[10][19] ), .IN2(\CARRYB[9][19] ), .IN3(\SUMB[9][20] ), .Q(\SUMB[10][19] ) );
  NAND2X0 U1645 ( .IN1(\ab[10][19] ), .IN2(\CARRYB[9][19] ), .QN(n796) );
  NAND2X1 U1646 ( .IN1(\ab[10][19] ), .IN2(\SUMB[9][20] ), .QN(n797) );
  NAND2X0 U1647 ( .IN1(\CARRYB[9][19] ), .IN2(\SUMB[9][20] ), .QN(n798) );
  NAND3X1 U1648 ( .IN1(n796), .IN2(n797), .IN3(n798), .QN(\CARRYB[10][19] ) );
  NAND2X0 U1649 ( .IN1(\ab[11][18] ), .IN2(\CARRYB[10][18] ), .QN(n799) );
  NAND2X0 U1650 ( .IN1(\ab[11][18] ), .IN2(\SUMB[10][19] ), .QN(n800) );
  NAND2X0 U1651 ( .IN1(\CARRYB[10][18] ), .IN2(\SUMB[10][19] ), .QN(n801) );
  XOR3X1 U1652 ( .IN1(\CARRYB[30][9] ), .IN2(\ab[31][9] ), .IN3(\SUMB[30][10] ), .Q(\SUMB[31][9] ) );
  NAND2X0 U1653 ( .IN1(\CARRYB[30][9] ), .IN2(\SUMB[30][10] ), .QN(n802) );
  NAND2X0 U1654 ( .IN1(\CARRYB[30][9] ), .IN2(\ab[31][9] ), .QN(n803) );
  NAND2X1 U1655 ( .IN1(\SUMB[30][10] ), .IN2(\ab[31][9] ), .QN(n804) );
  NAND3X0 U1656 ( .IN1(n802), .IN2(n803), .IN3(n804), .QN(\CARRYB[31][9] ) );
  XOR2X1 U1657 ( .IN1(\ab[27][9] ), .IN2(\CARRYB[26][9] ), .Q(n805) );
  NAND2X1 U1658 ( .IN1(\ab[26][10] ), .IN2(\CARRYB[25][10] ), .QN(n806) );
  NAND2X0 U1659 ( .IN1(\ab[26][10] ), .IN2(\SUMB[25][11] ), .QN(n807) );
  NAND2X0 U1660 ( .IN1(\CARRYB[25][10] ), .IN2(\SUMB[25][11] ), .QN(n808) );
  NAND2X0 U1661 ( .IN1(\ab[27][9] ), .IN2(\CARRYB[26][9] ), .QN(n809) );
  NAND2X0 U1662 ( .IN1(\ab[27][9] ), .IN2(\SUMB[26][10] ), .QN(n810) );
  NAND2X0 U1663 ( .IN1(\CARRYB[26][9] ), .IN2(\SUMB[26][10] ), .QN(n811) );
  XOR3X1 U1664 ( .IN1(\SUMB[22][11] ), .IN2(\ab[23][10] ), .IN3(
        \CARRYB[22][10] ), .Q(\SUMB[23][10] ) );
  NAND2X0 U1665 ( .IN1(\SUMB[22][11] ), .IN2(\CARRYB[22][10] ), .QN(n812) );
  NAND2X0 U1666 ( .IN1(\SUMB[22][11] ), .IN2(\ab[23][10] ), .QN(n813) );
  NAND2X0 U1667 ( .IN1(\CARRYB[22][10] ), .IN2(\ab[23][10] ), .QN(n814) );
  NAND3X0 U1668 ( .IN1(n812), .IN2(n813), .IN3(n814), .QN(\CARRYB[23][10] ) );
  XOR3X1 U1669 ( .IN1(\ab[3][17] ), .IN2(\CARRYB[2][17] ), .IN3(\SUMB[2][18] ), 
        .Q(\SUMB[3][17] ) );
  NAND2X0 U1670 ( .IN1(\ab[3][17] ), .IN2(\CARRYB[2][17] ), .QN(n815) );
  NAND2X1 U1671 ( .IN1(\ab[3][17] ), .IN2(\SUMB[2][18] ), .QN(n816) );
  NAND2X0 U1672 ( .IN1(\CARRYB[2][17] ), .IN2(\SUMB[2][18] ), .QN(n817) );
  NAND3X1 U1673 ( .IN1(n815), .IN2(n816), .IN3(n817), .QN(\CARRYB[3][17] ) );
  XOR2X1 U1674 ( .IN1(\ab[4][17] ), .IN2(\SUMB[3][18] ), .Q(n818) );
  NAND2X0 U1675 ( .IN1(\ab[4][17] ), .IN2(\SUMB[3][18] ), .QN(n819) );
  NAND2X0 U1676 ( .IN1(\ab[4][17] ), .IN2(\CARRYB[3][17] ), .QN(n820) );
  NAND2X0 U1677 ( .IN1(\SUMB[3][18] ), .IN2(\CARRYB[3][17] ), .QN(n821) );
  XOR3X1 U1678 ( .IN1(\ab[9][16] ), .IN2(\CARRYB[8][16] ), .IN3(\SUMB[8][17] ), 
        .Q(\SUMB[9][16] ) );
  NAND2X0 U1679 ( .IN1(\ab[9][16] ), .IN2(\CARRYB[8][16] ), .QN(n822) );
  NAND2X1 U1680 ( .IN1(\ab[9][16] ), .IN2(\SUMB[8][17] ), .QN(n823) );
  NAND2X0 U1681 ( .IN1(\CARRYB[8][16] ), .IN2(\SUMB[8][17] ), .QN(n824) );
  XOR2X1 U1682 ( .IN1(\ab[10][16] ), .IN2(\SUMB[9][17] ), .Q(n825) );
  XOR2X2 U1683 ( .IN1(n825), .IN2(\CARRYB[9][16] ), .Q(\SUMB[10][16] ) );
  NAND2X0 U1684 ( .IN1(\ab[10][16] ), .IN2(\SUMB[9][17] ), .QN(n826) );
  NAND2X0 U1685 ( .IN1(\ab[10][16] ), .IN2(\CARRYB[9][16] ), .QN(n827) );
  NAND2X0 U1686 ( .IN1(\SUMB[9][17] ), .IN2(\CARRYB[9][16] ), .QN(n828) );
  XOR3X1 U1687 ( .IN1(\ab[15][15] ), .IN2(\CARRYB[14][15] ), .IN3(
        \SUMB[14][16] ), .Q(\SUMB[15][15] ) );
  NAND2X0 U1688 ( .IN1(\ab[15][15] ), .IN2(\CARRYB[14][15] ), .QN(n829) );
  NAND2X1 U1689 ( .IN1(\ab[15][15] ), .IN2(\SUMB[14][16] ), .QN(n830) );
  NAND2X0 U1690 ( .IN1(\CARRYB[14][15] ), .IN2(\SUMB[14][16] ), .QN(n831) );
  NAND3X1 U1691 ( .IN1(n829), .IN2(n830), .IN3(n831), .QN(\CARRYB[15][15] ) );
  XOR2X1 U1692 ( .IN1(\ab[16][15] ), .IN2(\SUMB[15][16] ), .Q(n832) );
  NAND2X0 U1693 ( .IN1(\ab[16][15] ), .IN2(\SUMB[15][16] ), .QN(n833) );
  NAND2X0 U1694 ( .IN1(\ab[16][15] ), .IN2(\CARRYB[15][15] ), .QN(n834) );
  NAND2X0 U1695 ( .IN1(\SUMB[15][16] ), .IN2(\CARRYB[15][15] ), .QN(n835) );
  NAND3X1 U1696 ( .IN1(n833), .IN2(n834), .IN3(n835), .QN(\CARRYB[16][15] ) );
  XOR2X1 U1697 ( .IN1(\CARRYB[31][9] ), .IN2(\SUMB[31][10] ), .Q(\A1[39] ) );
  XOR3X1 U1698 ( .IN1(\ab[22][27] ), .IN2(\CARRYB[21][27] ), .IN3(
        \SUMB[21][28] ), .Q(\SUMB[22][27] ) );
  NAND2X1 U1699 ( .IN1(\ab[22][27] ), .IN2(\CARRYB[21][27] ), .QN(n837) );
  NAND2X0 U1700 ( .IN1(\ab[22][27] ), .IN2(\SUMB[21][28] ), .QN(n838) );
  NAND2X0 U1701 ( .IN1(\CARRYB[21][27] ), .IN2(\SUMB[21][28] ), .QN(n839) );
  NAND3X1 U1702 ( .IN1(n837), .IN2(n838), .IN3(n839), .QN(\CARRYB[22][27] ) );
  XOR2X1 U1703 ( .IN1(\ab[23][27] ), .IN2(\SUMB[22][28] ), .Q(n840) );
  XOR2X2 U1704 ( .IN1(n840), .IN2(\CARRYB[22][27] ), .Q(\SUMB[23][27] ) );
  NAND2X0 U1705 ( .IN1(\ab[23][27] ), .IN2(\SUMB[22][28] ), .QN(n841) );
  NAND2X0 U1706 ( .IN1(\ab[23][27] ), .IN2(\CARRYB[22][27] ), .QN(n842) );
  NAND2X0 U1707 ( .IN1(\SUMB[22][28] ), .IN2(\CARRYB[22][27] ), .QN(n843) );
  NAND3X1 U1708 ( .IN1(n841), .IN2(n842), .IN3(n843), .QN(\CARRYB[23][27] ) );
  XOR3X1 U1709 ( .IN1(\ab[13][30] ), .IN2(\CARRYB[12][30] ), .IN3(\ab[12][31] ), .Q(\SUMB[13][30] ) );
  NAND2X0 U1710 ( .IN1(\ab[13][30] ), .IN2(\CARRYB[12][30] ), .QN(n844) );
  NAND2X1 U1711 ( .IN1(\ab[13][30] ), .IN2(\ab[12][31] ), .QN(n845) );
  NAND2X0 U1712 ( .IN1(\CARRYB[12][30] ), .IN2(\ab[12][31] ), .QN(n846) );
  XOR2X1 U1713 ( .IN1(\ab[14][30] ), .IN2(\ab[13][31] ), .Q(n847) );
  XOR2X1 U1714 ( .IN1(n847), .IN2(\CARRYB[13][30] ), .Q(\SUMB[14][30] ) );
  NAND2X0 U1715 ( .IN1(\ab[14][30] ), .IN2(\ab[13][31] ), .QN(n848) );
  NAND2X0 U1716 ( .IN1(\ab[14][30] ), .IN2(\CARRYB[13][30] ), .QN(n849) );
  NAND2X0 U1717 ( .IN1(\ab[13][31] ), .IN2(\CARRYB[13][30] ), .QN(n850) );
  XOR3X1 U1718 ( .IN1(\ab[7][30] ), .IN2(\CARRYB[6][30] ), .IN3(\ab[6][31] ), 
        .Q(\SUMB[7][30] ) );
  NAND2X0 U1719 ( .IN1(\ab[7][30] ), .IN2(\CARRYB[6][30] ), .QN(n851) );
  NAND2X0 U1720 ( .IN1(\ab[7][30] ), .IN2(\ab[6][31] ), .QN(n852) );
  NAND2X0 U1721 ( .IN1(\CARRYB[6][30] ), .IN2(\ab[6][31] ), .QN(n853) );
  NAND3X1 U1722 ( .IN1(n851), .IN2(n852), .IN3(n853), .QN(\CARRYB[7][30] ) );
  XOR2X1 U1723 ( .IN1(n854), .IN2(\CARRYB[7][30] ), .Q(\SUMB[8][30] ) );
  NAND2X0 U1724 ( .IN1(\ab[8][30] ), .IN2(\ab[7][31] ), .QN(n855) );
  NAND2X0 U1725 ( .IN1(\ab[8][30] ), .IN2(\CARRYB[7][30] ), .QN(n856) );
  NAND2X0 U1726 ( .IN1(\ab[7][31] ), .IN2(\CARRYB[7][30] ), .QN(n857) );
  NAND3X1 U1727 ( .IN1(n855), .IN2(n856), .IN3(n857), .QN(\CARRYB[8][30] ) );
  XOR3X1 U1728 ( .IN1(\ab[5][3] ), .IN2(\CARRYB[4][3] ), .IN3(\SUMB[4][4] ), 
        .Q(\SUMB[5][3] ) );
  NAND2X0 U1729 ( .IN1(\ab[5][3] ), .IN2(\CARRYB[4][3] ), .QN(n858) );
  NAND2X1 U1730 ( .IN1(\ab[5][3] ), .IN2(\SUMB[4][4] ), .QN(n859) );
  NAND2X0 U1731 ( .IN1(\CARRYB[4][3] ), .IN2(\SUMB[4][4] ), .QN(n860) );
  XOR2X1 U1732 ( .IN1(\ab[6][3] ), .IN2(\SUMB[5][4] ), .Q(n861) );
  NAND2X0 U1733 ( .IN1(\ab[6][3] ), .IN2(\SUMB[5][4] ), .QN(n862) );
  NAND2X0 U1734 ( .IN1(\ab[6][3] ), .IN2(\CARRYB[5][3] ), .QN(n863) );
  NAND2X0 U1735 ( .IN1(\SUMB[5][4] ), .IN2(\CARRYB[5][3] ), .QN(n864) );
  DELLN1X2 U1736 ( .INP(n2209), .Z(n2095) );
  XOR3X1 U1737 ( .IN1(\ab[29][16] ), .IN2(\CARRYB[28][16] ), .IN3(
        \SUMB[28][17] ), .Q(\SUMB[29][16] ) );
  NAND2X0 U1738 ( .IN1(\ab[29][16] ), .IN2(\SUMB[28][17] ), .QN(n866) );
  NAND2X0 U1739 ( .IN1(\CARRYB[28][16] ), .IN2(\SUMB[28][17] ), .QN(n867) );
  XOR2X1 U1740 ( .IN1(\ab[30][16] ), .IN2(\SUMB[29][17] ), .Q(n868) );
  NAND2X0 U1741 ( .IN1(\ab[30][16] ), .IN2(\SUMB[29][17] ), .QN(n869) );
  NAND2X0 U1742 ( .IN1(\ab[30][16] ), .IN2(\CARRYB[29][16] ), .QN(n870) );
  NAND2X0 U1743 ( .IN1(\SUMB[29][17] ), .IN2(\CARRYB[29][16] ), .QN(n871) );
  XOR3X1 U1744 ( .IN1(\CARRYB[27][17] ), .IN2(\ab[28][17] ), .IN3(
        \SUMB[27][18] ), .Q(\SUMB[28][17] ) );
  NAND2X0 U1745 ( .IN1(\CARRYB[27][17] ), .IN2(\SUMB[27][18] ), .QN(n872) );
  NAND2X1 U1746 ( .IN1(\CARRYB[27][17] ), .IN2(\ab[28][17] ), .QN(n873) );
  NAND2X0 U1747 ( .IN1(\SUMB[27][18] ), .IN2(\ab[28][17] ), .QN(n874) );
  XOR3X1 U1748 ( .IN1(\CARRYB[9][18] ), .IN2(\ab[10][18] ), .IN3(\SUMB[9][19] ), .Q(\SUMB[10][18] ) );
  NAND2X0 U1749 ( .IN1(\CARRYB[9][18] ), .IN2(\SUMB[9][19] ), .QN(n875) );
  NAND2X0 U1750 ( .IN1(\CARRYB[9][18] ), .IN2(\ab[10][18] ), .QN(n876) );
  NAND2X0 U1751 ( .IN1(\SUMB[9][19] ), .IN2(\ab[10][18] ), .QN(n877) );
  XOR3X1 U1752 ( .IN1(\CARRYB[8][18] ), .IN2(\ab[9][18] ), .IN3(\SUMB[8][19] ), 
        .Q(\SUMB[9][18] ) );
  NAND2X0 U1753 ( .IN1(\CARRYB[8][18] ), .IN2(\SUMB[8][19] ), .QN(n878) );
  NAND2X1 U1754 ( .IN1(\CARRYB[8][18] ), .IN2(\ab[9][18] ), .QN(n879) );
  NAND2X0 U1755 ( .IN1(\SUMB[8][19] ), .IN2(\ab[9][18] ), .QN(n880) );
  NAND3X1 U1756 ( .IN1(n878), .IN2(n879), .IN3(n880), .QN(\CARRYB[9][18] ) );
  DELLN1X2 U1757 ( .INP(n2209), .Z(n2096) );
  XOR3X1 U1758 ( .IN1(\ab[30][21] ), .IN2(\CARRYB[29][21] ), .IN3(
        \SUMB[29][22] ), .Q(\SUMB[30][21] ) );
  NAND2X0 U1759 ( .IN1(\ab[30][21] ), .IN2(\CARRYB[29][21] ), .QN(n881) );
  NAND2X1 U1760 ( .IN1(\ab[30][21] ), .IN2(\SUMB[29][22] ), .QN(n882) );
  NAND2X0 U1761 ( .IN1(\CARRYB[29][21] ), .IN2(\SUMB[29][22] ), .QN(n883) );
  XOR2X1 U1762 ( .IN1(\ab[31][21] ), .IN2(\SUMB[30][22] ), .Q(n884) );
  NAND2X0 U1763 ( .IN1(\ab[31][21] ), .IN2(\SUMB[30][22] ), .QN(n885) );
  NAND2X0 U1764 ( .IN1(\ab[31][21] ), .IN2(\CARRYB[30][21] ), .QN(n886) );
  NAND2X0 U1765 ( .IN1(\SUMB[30][22] ), .IN2(\CARRYB[30][21] ), .QN(n887) );
  XOR3X1 U1766 ( .IN1(\ab[22][24] ), .IN2(\CARRYB[21][24] ), .IN3(
        \SUMB[21][25] ), .Q(\SUMB[22][24] ) );
  NAND2X0 U1767 ( .IN1(\ab[22][24] ), .IN2(\CARRYB[21][24] ), .QN(n888) );
  NAND2X1 U1768 ( .IN1(\ab[22][24] ), .IN2(\SUMB[21][25] ), .QN(n889) );
  NAND2X0 U1769 ( .IN1(\CARRYB[21][24] ), .IN2(\SUMB[21][25] ), .QN(n890) );
  XOR2X1 U1770 ( .IN1(\ab[23][24] ), .IN2(\SUMB[22][25] ), .Q(n891) );
  XOR2X2 U1771 ( .IN1(n891), .IN2(\CARRYB[22][24] ), .Q(\SUMB[23][24] ) );
  NAND2X0 U1772 ( .IN1(\ab[23][24] ), .IN2(\SUMB[22][25] ), .QN(n892) );
  NAND2X0 U1773 ( .IN1(\ab[23][24] ), .IN2(\CARRYB[22][24] ), .QN(n893) );
  NAND2X0 U1774 ( .IN1(\SUMB[22][25] ), .IN2(\CARRYB[22][24] ), .QN(n894) );
  XOR3X1 U1775 ( .IN1(\CARRYB[28][21] ), .IN2(\ab[29][21] ), .IN3(
        \SUMB[28][22] ), .Q(\SUMB[29][21] ) );
  NAND2X0 U1776 ( .IN1(\CARRYB[28][21] ), .IN2(\SUMB[28][22] ), .QN(n895) );
  NAND2X0 U1777 ( .IN1(\CARRYB[28][21] ), .IN2(\ab[29][21] ), .QN(n896) );
  NAND2X0 U1778 ( .IN1(\SUMB[28][22] ), .IN2(\ab[29][21] ), .QN(n897) );
  XOR3X1 U1779 ( .IN1(\ab[16][24] ), .IN2(\CARRYB[15][24] ), .IN3(
        \SUMB[15][25] ), .Q(\SUMB[16][24] ) );
  NAND2X1 U1780 ( .IN1(\ab[16][24] ), .IN2(\CARRYB[15][24] ), .QN(n898) );
  NAND2X0 U1781 ( .IN1(\ab[16][24] ), .IN2(\SUMB[15][25] ), .QN(n899) );
  NAND2X0 U1782 ( .IN1(\CARRYB[15][24] ), .IN2(\SUMB[15][25] ), .QN(n900) );
  XOR2X1 U1783 ( .IN1(\ab[17][24] ), .IN2(\SUMB[16][25] ), .Q(n901) );
  NAND2X0 U1784 ( .IN1(\ab[17][24] ), .IN2(\SUMB[16][25] ), .QN(n902) );
  NAND2X0 U1785 ( .IN1(\ab[17][24] ), .IN2(\CARRYB[16][24] ), .QN(n903) );
  NAND2X0 U1786 ( .IN1(\SUMB[16][25] ), .IN2(\CARRYB[16][24] ), .QN(n904) );
  XOR3X1 U1787 ( .IN1(\ab[11][26] ), .IN2(\CARRYB[10][26] ), .IN3(
        \SUMB[10][27] ), .Q(\SUMB[11][26] ) );
  NAND2X0 U1788 ( .IN1(\ab[11][26] ), .IN2(\CARRYB[10][26] ), .QN(n905) );
  NAND2X1 U1789 ( .IN1(\ab[11][26] ), .IN2(\SUMB[10][27] ), .QN(n906) );
  NAND2X0 U1790 ( .IN1(\CARRYB[10][26] ), .IN2(\SUMB[10][27] ), .QN(n907) );
  XOR2X1 U1791 ( .IN1(\ab[12][26] ), .IN2(\SUMB[11][27] ), .Q(n908) );
  NAND2X0 U1792 ( .IN1(\ab[12][26] ), .IN2(\SUMB[11][27] ), .QN(n909) );
  NAND2X0 U1793 ( .IN1(\ab[12][26] ), .IN2(\CARRYB[11][26] ), .QN(n910) );
  NAND2X0 U1794 ( .IN1(\SUMB[11][27] ), .IN2(\CARRYB[11][26] ), .QN(n911) );
  XOR3X1 U1795 ( .IN1(\CARRYB[9][26] ), .IN2(\ab[10][26] ), .IN3(\SUMB[9][27] ), .Q(\SUMB[10][26] ) );
  NAND2X0 U1796 ( .IN1(\CARRYB[9][26] ), .IN2(\SUMB[9][27] ), .QN(n912) );
  NAND2X0 U1797 ( .IN1(\CARRYB[9][26] ), .IN2(\ab[10][26] ), .QN(n913) );
  NAND2X1 U1798 ( .IN1(\SUMB[9][27] ), .IN2(\ab[10][26] ), .QN(n914) );
  XOR3X1 U1799 ( .IN1(\CARRYB[5][27] ), .IN2(\ab[6][27] ), .IN3(\SUMB[5][28] ), 
        .Q(\SUMB[6][27] ) );
  NAND2X0 U1800 ( .IN1(\CARRYB[5][27] ), .IN2(\SUMB[5][28] ), .QN(n915) );
  NAND2X1 U1801 ( .IN1(\CARRYB[5][27] ), .IN2(\ab[6][27] ), .QN(n916) );
  NAND2X0 U1802 ( .IN1(\SUMB[5][28] ), .IN2(\ab[6][27] ), .QN(n917) );
  XOR3X1 U1803 ( .IN1(\ab[18][0] ), .IN2(\CARRYB[17][0] ), .IN3(\SUMB[17][1] ), 
        .Q(\A1[16] ) );
  NAND2X0 U1804 ( .IN1(\ab[18][0] ), .IN2(\CARRYB[17][0] ), .QN(n918) );
  NAND2X0 U1805 ( .IN1(\ab[18][0] ), .IN2(\SUMB[17][1] ), .QN(n919) );
  NAND2X0 U1806 ( .IN1(\CARRYB[17][0] ), .IN2(\SUMB[17][1] ), .QN(n920) );
  XOR2X1 U1807 ( .IN1(n921), .IN2(n62), .Q(\A1[17] ) );
  NAND2X0 U1808 ( .IN1(\ab[19][0] ), .IN2(\SUMB[18][1] ), .QN(n922) );
  NAND2X0 U1809 ( .IN1(\ab[19][0] ), .IN2(\CARRYB[18][0] ), .QN(n923) );
  NAND2X0 U1810 ( .IN1(\SUMB[18][1] ), .IN2(n62), .QN(n924) );
  XOR3X1 U1811 ( .IN1(\ab[12][2] ), .IN2(\CARRYB[11][2] ), .IN3(\SUMB[11][3] ), 
        .Q(\SUMB[12][2] ) );
  XOR2X1 U1812 ( .IN1(\ab[13][1] ), .IN2(\CARRYB[12][1] ), .Q(n925) );
  NAND2X0 U1813 ( .IN1(\ab[12][2] ), .IN2(\CARRYB[11][2] ), .QN(n926) );
  NAND2X0 U1814 ( .IN1(\ab[12][2] ), .IN2(\SUMB[11][3] ), .QN(n927) );
  NAND2X0 U1815 ( .IN1(\CARRYB[11][2] ), .IN2(\SUMB[11][3] ), .QN(n928) );
  NAND3X1 U1816 ( .IN1(n926), .IN2(n927), .IN3(n928), .QN(\CARRYB[12][2] ) );
  NAND2X0 U1817 ( .IN1(\ab[13][1] ), .IN2(\CARRYB[12][1] ), .QN(n929) );
  NAND2X0 U1818 ( .IN1(\ab[13][1] ), .IN2(\SUMB[12][2] ), .QN(n930) );
  NAND2X0 U1819 ( .IN1(\CARRYB[12][1] ), .IN2(\SUMB[12][2] ), .QN(n931) );
  NAND3X1 U1820 ( .IN1(n929), .IN2(n930), .IN3(n931), .QN(\CARRYB[13][1] ) );
  AND2X1 U1821 ( .IN1(\ab[0][28] ), .IN2(\ab[1][27] ), .Q(n963) );
  XOR2X1 U1822 ( .IN1(\ab[15][3] ), .IN2(\SUMB[14][4] ), .Q(n932) );
  XOR2X1 U1823 ( .IN1(n932), .IN2(\CARRYB[14][3] ), .Q(\SUMB[15][3] ) );
  NOR2X0 U1824 ( .IN1(n2099), .IN2(n2003), .QN(n933) );
  DELLN1X2 U1825 ( .INP(n2211), .Z(n2099) );
  XOR3X1 U1826 ( .IN1(\ab[6][15] ), .IN2(\CARRYB[5][15] ), .IN3(\SUMB[5][16] ), 
        .Q(\SUMB[6][15] ) );
  NAND2X0 U1827 ( .IN1(\ab[6][15] ), .IN2(\CARRYB[5][15] ), .QN(n934) );
  NAND2X1 U1828 ( .IN1(\ab[6][15] ), .IN2(\SUMB[5][16] ), .QN(n935) );
  NAND2X0 U1829 ( .IN1(\CARRYB[5][15] ), .IN2(\SUMB[5][16] ), .QN(n936) );
  NAND2X0 U1830 ( .IN1(\ab[7][14] ), .IN2(\CARRYB[6][14] ), .QN(n937) );
  NAND2X0 U1831 ( .IN1(\ab[7][14] ), .IN2(\SUMB[6][15] ), .QN(n938) );
  NAND2X0 U1832 ( .IN1(\CARRYB[6][14] ), .IN2(\SUMB[6][15] ), .QN(n939) );
  XOR3X1 U1833 ( .IN1(\ab[2][15] ), .IN2(n15), .IN3(\SUMB[1][16] ), .Q(
        \SUMB[2][15] ) );
  NAND2X0 U1834 ( .IN1(\ab[2][15] ), .IN2(n15), .QN(n940) );
  NAND2X1 U1835 ( .IN1(\ab[2][15] ), .IN2(\SUMB[1][16] ), .QN(n941) );
  NAND2X0 U1836 ( .IN1(n15), .IN2(\SUMB[1][16] ), .QN(n942) );
  NAND3X1 U1837 ( .IN1(n940), .IN2(n941), .IN3(n942), .QN(\CARRYB[2][15] ) );
  XOR2X1 U1838 ( .IN1(\ab[3][15] ), .IN2(\SUMB[2][16] ), .Q(n943) );
  NAND2X0 U1839 ( .IN1(\ab[3][15] ), .IN2(\SUMB[2][16] ), .QN(n944) );
  NAND2X0 U1840 ( .IN1(\ab[3][15] ), .IN2(\CARRYB[2][15] ), .QN(n945) );
  NAND2X0 U1841 ( .IN1(\SUMB[2][16] ), .IN2(\CARRYB[2][15] ), .QN(n946) );
  NAND3X1 U1842 ( .IN1(n944), .IN2(n945), .IN3(n946), .QN(\CARRYB[3][15] ) );
  DELLN1X2 U1843 ( .INP(n2224), .Z(n2137) );
  DELLN1X2 U1844 ( .INP(n2224), .Z(n2139) );
  NAND2X0 U1845 ( .IN1(\ab[17][1] ), .IN2(\SUMB[16][2] ), .QN(n1433) );
  AND2X1 U1846 ( .IN1(\ab[0][3] ), .IN2(\ab[1][2] ), .Q(n947) );
  XOR3X1 U1847 ( .IN1(\ab[16][5] ), .IN2(\CARRYB[15][5] ), .IN3(\SUMB[15][6] ), 
        .Q(\SUMB[16][5] ) );
  NAND2X0 U1848 ( .IN1(\ab[16][5] ), .IN2(\CARRYB[15][5] ), .QN(n949) );
  NAND2X1 U1849 ( .IN1(\ab[16][5] ), .IN2(\SUMB[15][6] ), .QN(n950) );
  NAND2X0 U1850 ( .IN1(\CARRYB[15][5] ), .IN2(\SUMB[15][6] ), .QN(n951) );
  NAND3X1 U1851 ( .IN1(n949), .IN2(n950), .IN3(n951), .QN(\CARRYB[16][5] ) );
  XOR2X1 U1852 ( .IN1(\ab[17][5] ), .IN2(\SUMB[16][6] ), .Q(n952) );
  NAND2X0 U1853 ( .IN1(\ab[17][5] ), .IN2(\SUMB[16][6] ), .QN(n953) );
  NAND2X0 U1854 ( .IN1(\ab[17][5] ), .IN2(\CARRYB[16][5] ), .QN(n954) );
  NAND2X0 U1855 ( .IN1(\SUMB[16][6] ), .IN2(\CARRYB[16][5] ), .QN(n955) );
  NAND3X1 U1856 ( .IN1(n953), .IN2(n954), .IN3(n955), .QN(\CARRYB[17][5] ) );
  XOR3X1 U1857 ( .IN1(\ab[6][18] ), .IN2(\CARRYB[5][18] ), .IN3(\SUMB[5][19] ), 
        .Q(\SUMB[6][18] ) );
  NAND2X1 U1858 ( .IN1(\ab[6][18] ), .IN2(\CARRYB[5][18] ), .QN(n956) );
  NAND2X0 U1859 ( .IN1(\ab[6][18] ), .IN2(\SUMB[5][19] ), .QN(n957) );
  NAND2X0 U1860 ( .IN1(\CARRYB[5][18] ), .IN2(\SUMB[5][19] ), .QN(n958) );
  NAND3X1 U1861 ( .IN1(n956), .IN2(n957), .IN3(n958), .QN(\CARRYB[6][18] ) );
  XOR2X1 U1862 ( .IN1(\ab[7][18] ), .IN2(\SUMB[6][19] ), .Q(n959) );
  NAND2X0 U1863 ( .IN1(\ab[7][18] ), .IN2(\SUMB[6][19] ), .QN(n960) );
  NAND2X0 U1864 ( .IN1(\ab[7][18] ), .IN2(\CARRYB[6][18] ), .QN(n961) );
  NAND2X0 U1865 ( .IN1(\SUMB[6][19] ), .IN2(\CARRYB[6][18] ), .QN(n962) );
  NAND2X0 U1866 ( .IN1(\ab[21][0] ), .IN2(\CARRYB[20][0] ), .QN(n1954) );
  NAND2X0 U1867 ( .IN1(\CARRYB[20][0] ), .IN2(\SUMB[20][1] ), .QN(n1956) );
  XOR3X1 U1868 ( .IN1(\CARRYB[29][0] ), .IN2(\ab[30][0] ), .IN3(\SUMB[29][1] ), 
        .Q(\A1[28] ) );
  DELLN1X2 U1869 ( .INP(n2219), .Z(n2123) );
  NAND2X0 U1870 ( .IN1(\SUMB[15][15] ), .IN2(\CARRYB[15][14] ), .QN(n964) );
  NAND2X0 U1871 ( .IN1(\SUMB[15][15] ), .IN2(\ab[16][14] ), .QN(n965) );
  NAND2X0 U1872 ( .IN1(\CARRYB[15][14] ), .IN2(\ab[16][14] ), .QN(n966) );
  NAND2X0 U1873 ( .IN1(\CARRYB[29][0] ), .IN2(\ab[30][0] ), .QN(n1969) );
  XOR3X1 U1874 ( .IN1(\ab[10][29] ), .IN2(\CARRYB[9][29] ), .IN3(\SUMB[9][30] ), .Q(\SUMB[10][29] ) );
  NAND2X0 U1875 ( .IN1(\ab[10][29] ), .IN2(\CARRYB[9][29] ), .QN(n967) );
  NAND2X1 U1876 ( .IN1(\ab[10][29] ), .IN2(\SUMB[9][30] ), .QN(n968) );
  NAND2X0 U1877 ( .IN1(\CARRYB[9][29] ), .IN2(\SUMB[9][30] ), .QN(n969) );
  NAND3X1 U1878 ( .IN1(n967), .IN2(n968), .IN3(n969), .QN(\CARRYB[10][29] ) );
  XOR2X1 U1879 ( .IN1(\ab[11][29] ), .IN2(\SUMB[10][30] ), .Q(n970) );
  NAND2X0 U1880 ( .IN1(\ab[11][29] ), .IN2(\SUMB[10][30] ), .QN(n971) );
  NAND2X0 U1881 ( .IN1(\ab[11][29] ), .IN2(\CARRYB[10][29] ), .QN(n972) );
  NAND2X0 U1882 ( .IN1(\SUMB[10][30] ), .IN2(n349), .QN(n973) );
  NAND3X1 U1883 ( .IN1(n971), .IN2(n972), .IN3(n973), .QN(\CARRYB[11][29] ) );
  XOR3X1 U1884 ( .IN1(\ab[31][0] ), .IN2(\SUMB[30][1] ), .IN3(\CARRYB[30][0] ), 
        .Q(\SUMB[31][0] ) );
  XNOR2X2 U1885 ( .IN1(n974), .IN2(\CARRYB[24][26] ), .Q(\SUMB[25][26] ) );
  XNOR2X1 U1886 ( .IN1(\ab[25][26] ), .IN2(\SUMB[24][27] ), .Q(n974) );
  DELLN1X2 U1887 ( .INP(n2210), .Z(n2097) );
  XOR3X1 U1888 ( .IN1(\ab[17][11] ), .IN2(\CARRYB[16][11] ), .IN3(
        \SUMB[16][12] ), .Q(\SUMB[17][11] ) );
  NAND2X1 U1889 ( .IN1(\ab[17][11] ), .IN2(\CARRYB[16][11] ), .QN(n975) );
  NAND2X0 U1890 ( .IN1(\ab[17][11] ), .IN2(\SUMB[16][12] ), .QN(n976) );
  NAND2X0 U1891 ( .IN1(\CARRYB[16][11] ), .IN2(\SUMB[16][12] ), .QN(n977) );
  NAND3X1 U1892 ( .IN1(n975), .IN2(n976), .IN3(n977), .QN(\CARRYB[17][11] ) );
  XOR2X1 U1893 ( .IN1(\ab[18][11] ), .IN2(\SUMB[17][12] ), .Q(n978) );
  NAND2X0 U1894 ( .IN1(\ab[18][11] ), .IN2(\SUMB[17][12] ), .QN(n979) );
  NAND2X0 U1895 ( .IN1(\ab[18][11] ), .IN2(\CARRYB[17][11] ), .QN(n980) );
  NAND2X0 U1896 ( .IN1(\SUMB[17][12] ), .IN2(\CARRYB[17][11] ), .QN(n981) );
  XOR3X1 U1897 ( .IN1(\CARRYB[4][16] ), .IN2(\ab[5][16] ), .IN3(\SUMB[4][17] ), 
        .Q(\SUMB[5][16] ) );
  NAND2X1 U1898 ( .IN1(\CARRYB[4][16] ), .IN2(\ab[5][16] ), .QN(n982) );
  NAND2X0 U1899 ( .IN1(\CARRYB[4][16] ), .IN2(\SUMB[4][17] ), .QN(n983) );
  NAND2X0 U1900 ( .IN1(\ab[5][16] ), .IN2(\SUMB[4][17] ), .QN(n984) );
  XOR2X1 U1901 ( .IN1(\ab[6][16] ), .IN2(\SUMB[5][17] ), .Q(n985) );
  NAND2X0 U1902 ( .IN1(\ab[6][16] ), .IN2(\SUMB[5][17] ), .QN(n986) );
  NAND2X0 U1903 ( .IN1(\ab[6][16] ), .IN2(\CARRYB[5][16] ), .QN(n987) );
  NAND2X0 U1904 ( .IN1(\SUMB[5][17] ), .IN2(\CARRYB[5][16] ), .QN(n988) );
  XOR3X1 U1905 ( .IN1(\ab[3][16] ), .IN2(\CARRYB[2][16] ), .IN3(\SUMB[2][17] ), 
        .Q(\SUMB[3][16] ) );
  NAND2X0 U1906 ( .IN1(\ab[3][16] ), .IN2(\CARRYB[2][16] ), .QN(n989) );
  NAND2X1 U1907 ( .IN1(\ab[3][16] ), .IN2(\SUMB[2][17] ), .QN(n990) );
  NAND2X0 U1908 ( .IN1(\CARRYB[2][16] ), .IN2(\SUMB[2][17] ), .QN(n991) );
  XOR2X1 U1909 ( .IN1(\ab[4][16] ), .IN2(\SUMB[3][17] ), .Q(n992) );
  NAND2X0 U1910 ( .IN1(\ab[4][16] ), .IN2(\SUMB[3][17] ), .QN(n993) );
  NAND2X0 U1911 ( .IN1(\ab[4][16] ), .IN2(\CARRYB[3][16] ), .QN(n994) );
  NAND2X0 U1912 ( .IN1(\SUMB[3][17] ), .IN2(\CARRYB[3][16] ), .QN(n995) );
  XOR3X1 U1913 ( .IN1(\ab[28][18] ), .IN2(\CARRYB[27][18] ), .IN3(
        \SUMB[27][19] ), .Q(\SUMB[28][18] ) );
  NAND2X0 U1914 ( .IN1(\ab[28][18] ), .IN2(\CARRYB[27][18] ), .QN(n996) );
  NAND2X1 U1915 ( .IN1(\ab[28][18] ), .IN2(\SUMB[27][19] ), .QN(n997) );
  NAND2X0 U1916 ( .IN1(\CARRYB[27][18] ), .IN2(\SUMB[27][19] ), .QN(n998) );
  NAND3X1 U1917 ( .IN1(n996), .IN2(n997), .IN3(n998), .QN(\CARRYB[28][18] ) );
  XOR2X1 U1918 ( .IN1(\ab[29][18] ), .IN2(\SUMB[28][19] ), .Q(n999) );
  NAND2X0 U1919 ( .IN1(\ab[29][18] ), .IN2(\SUMB[28][19] ), .QN(n1000) );
  NAND2X0 U1920 ( .IN1(\ab[29][18] ), .IN2(\CARRYB[28][18] ), .QN(n1001) );
  NAND2X0 U1921 ( .IN1(\SUMB[28][19] ), .IN2(\CARRYB[28][18] ), .QN(n1002) );
  XOR3X1 U1922 ( .IN1(\CARRYB[9][23] ), .IN2(\ab[10][23] ), .IN3(\SUMB[9][24] ), .Q(\SUMB[10][23] ) );
  NAND2X0 U1923 ( .IN1(\CARRYB[9][23] ), .IN2(\SUMB[9][24] ), .QN(n1003) );
  NAND2X0 U1924 ( .IN1(\CARRYB[9][23] ), .IN2(\ab[10][23] ), .QN(n1004) );
  XOR3X1 U1925 ( .IN1(\ab[12][23] ), .IN2(\CARRYB[11][23] ), .IN3(
        \SUMB[11][24] ), .Q(\SUMB[12][23] ) );
  NAND2X1 U1926 ( .IN1(\ab[12][23] ), .IN2(\CARRYB[11][23] ), .QN(n1006) );
  NAND2X0 U1927 ( .IN1(\ab[12][23] ), .IN2(\SUMB[11][24] ), .QN(n1007) );
  NAND2X0 U1928 ( .IN1(\CARRYB[11][23] ), .IN2(\SUMB[11][24] ), .QN(n1008) );
  XOR2X1 U1929 ( .IN1(\ab[13][23] ), .IN2(\SUMB[12][24] ), .Q(n1009) );
  NAND2X0 U1930 ( .IN1(\ab[13][23] ), .IN2(\SUMB[12][24] ), .QN(n1010) );
  NAND2X0 U1931 ( .IN1(\ab[13][23] ), .IN2(\CARRYB[12][23] ), .QN(n1011) );
  NAND2X0 U1932 ( .IN1(\SUMB[12][24] ), .IN2(\CARRYB[12][23] ), .QN(n1012) );
  XOR2X1 U1933 ( .IN1(\ab[21][19] ), .IN2(\CARRYB[20][19] ), .Q(n1013) );
  NAND2X0 U1934 ( .IN1(\SUMB[20][20] ), .IN2(\CARRYB[20][19] ), .QN(n1014) );
  NAND2X0 U1935 ( .IN1(\SUMB[20][20] ), .IN2(\ab[21][19] ), .QN(n1015) );
  NAND2X1 U1936 ( .IN1(\CARRYB[20][19] ), .IN2(\ab[21][19] ), .QN(n1016) );
  XOR2X1 U1937 ( .IN1(n1494), .IN2(\CARRYB[8][24] ), .Q(\SUMB[9][24] ) );
  XOR2X2 U1938 ( .IN1(\ab[1][16] ), .IN2(\ab[0][17] ), .Q(\SUMB[1][16] ) );
  XOR3X1 U1939 ( .IN1(\ab[4][26] ), .IN2(\CARRYB[3][26] ), .IN3(\SUMB[3][27] ), 
        .Q(\SUMB[4][26] ) );
  NAND2X0 U1940 ( .IN1(\ab[4][26] ), .IN2(\CARRYB[3][26] ), .QN(n1017) );
  NAND2X1 U1941 ( .IN1(\ab[4][26] ), .IN2(\SUMB[3][27] ), .QN(n1018) );
  NAND2X0 U1942 ( .IN1(\CARRYB[3][26] ), .IN2(\SUMB[3][27] ), .QN(n1019) );
  NAND3X1 U1943 ( .IN1(n1017), .IN2(n1018), .IN3(n1019), .QN(\CARRYB[4][26] )
         );
  XOR2X1 U1944 ( .IN1(\ab[5][26] ), .IN2(\SUMB[4][27] ), .Q(n1020) );
  NAND2X0 U1945 ( .IN1(\ab[5][26] ), .IN2(\SUMB[4][27] ), .QN(n1021) );
  NAND2X0 U1946 ( .IN1(\ab[5][26] ), .IN2(\CARRYB[4][26] ), .QN(n1022) );
  NAND2X0 U1947 ( .IN1(\SUMB[4][27] ), .IN2(\CARRYB[4][26] ), .QN(n1023) );
  XOR3X1 U1948 ( .IN1(\CARRYB[2][26] ), .IN2(\ab[3][26] ), .IN3(\SUMB[2][27] ), 
        .Q(\SUMB[3][26] ) );
  NAND2X0 U1949 ( .IN1(\CARRYB[2][26] ), .IN2(\SUMB[2][27] ), .QN(n1024) );
  NAND2X0 U1950 ( .IN1(\CARRYB[2][26] ), .IN2(\ab[3][26] ), .QN(n1025) );
  NAND2X0 U1951 ( .IN1(\SUMB[2][27] ), .IN2(\ab[3][26] ), .QN(n1026) );
  DELLN1X2 U1952 ( .INP(n2213), .Z(n2104) );
  XOR3X1 U1953 ( .IN1(\ab[18][26] ), .IN2(\CARRYB[17][26] ), .IN3(
        \SUMB[17][27] ), .Q(\SUMB[18][26] ) );
  XOR2X1 U1954 ( .IN1(\ab[19][25] ), .IN2(\CARRYB[18][25] ), .Q(n1028) );
  NAND2X0 U1955 ( .IN1(\ab[18][26] ), .IN2(\CARRYB[17][26] ), .QN(n1029) );
  NAND2X1 U1956 ( .IN1(\ab[18][26] ), .IN2(\SUMB[17][27] ), .QN(n1030) );
  NAND2X0 U1957 ( .IN1(\CARRYB[17][26] ), .IN2(\SUMB[17][27] ), .QN(n1031) );
  NAND2X0 U1958 ( .IN1(\ab[19][25] ), .IN2(\CARRYB[18][25] ), .QN(n1032) );
  NAND2X0 U1959 ( .IN1(\ab[19][25] ), .IN2(\SUMB[18][26] ), .QN(n1033) );
  NAND2X0 U1960 ( .IN1(\CARRYB[18][25] ), .IN2(\SUMB[18][26] ), .QN(n1034) );
  XOR3X1 U1961 ( .IN1(\ab[13][26] ), .IN2(\CARRYB[12][26] ), .IN3(
        \SUMB[12][27] ), .Q(\SUMB[13][26] ) );
  NAND2X0 U1962 ( .IN1(\ab[13][26] ), .IN2(\CARRYB[12][26] ), .QN(n1035) );
  NAND2X1 U1963 ( .IN1(\ab[13][26] ), .IN2(\SUMB[12][27] ), .QN(n1036) );
  NAND2X0 U1964 ( .IN1(\CARRYB[12][26] ), .IN2(\SUMB[12][27] ), .QN(n1037) );
  XOR2X1 U1965 ( .IN1(\ab[14][26] ), .IN2(\SUMB[13][27] ), .Q(n1038) );
  NAND2X0 U1966 ( .IN1(\ab[14][26] ), .IN2(\SUMB[13][27] ), .QN(n1039) );
  NAND2X0 U1967 ( .IN1(\ab[14][26] ), .IN2(\CARRYB[13][26] ), .QN(n1040) );
  NAND2X0 U1968 ( .IN1(\SUMB[13][27] ), .IN2(\CARRYB[13][26] ), .QN(n1041) );
  XOR3X1 U1969 ( .IN1(\ab[14][7] ), .IN2(\CARRYB[13][7] ), .IN3(\SUMB[13][8] ), 
        .Q(\SUMB[14][7] ) );
  NAND2X0 U1970 ( .IN1(\ab[14][7] ), .IN2(\CARRYB[13][7] ), .QN(n1042) );
  NAND2X0 U1971 ( .IN1(\ab[14][7] ), .IN2(\SUMB[13][8] ), .QN(n1043) );
  NAND2X0 U1972 ( .IN1(\CARRYB[13][7] ), .IN2(\SUMB[13][8] ), .QN(n1044) );
  NAND3X1 U1973 ( .IN1(n1042), .IN2(n1043), .IN3(n1044), .QN(\CARRYB[14][7] )
         );
  XOR2X1 U1974 ( .IN1(n1045), .IN2(\CARRYB[14][7] ), .Q(\SUMB[15][7] ) );
  NAND2X0 U1975 ( .IN1(\ab[15][7] ), .IN2(\SUMB[14][8] ), .QN(n1046) );
  NAND2X0 U1976 ( .IN1(\ab[15][7] ), .IN2(\CARRYB[14][7] ), .QN(n1047) );
  NAND2X0 U1977 ( .IN1(\SUMB[14][8] ), .IN2(\CARRYB[14][7] ), .QN(n1048) );
  NAND3X1 U1978 ( .IN1(n1046), .IN2(n1047), .IN3(n1048), .QN(\CARRYB[15][7] )
         );
  XOR3X1 U1979 ( .IN1(\ab[3][9] ), .IN2(\CARRYB[2][9] ), .IN3(\SUMB[2][10] ), 
        .Q(\SUMB[3][9] ) );
  NAND2X0 U1980 ( .IN1(\ab[3][9] ), .IN2(\CARRYB[2][9] ), .QN(n1049) );
  NAND2X1 U1981 ( .IN1(\ab[3][9] ), .IN2(\SUMB[2][10] ), .QN(n1050) );
  NAND2X0 U1982 ( .IN1(\CARRYB[2][9] ), .IN2(\SUMB[2][10] ), .QN(n1051) );
  NAND3X1 U1983 ( .IN1(n1049), .IN2(n1050), .IN3(n1051), .QN(\CARRYB[3][9] )
         );
  XOR2X1 U1984 ( .IN1(\ab[4][9] ), .IN2(\SUMB[3][10] ), .Q(n1052) );
  XOR2X2 U1985 ( .IN1(n1052), .IN2(\CARRYB[3][9] ), .Q(\SUMB[4][9] ) );
  NAND2X0 U1986 ( .IN1(\ab[4][9] ), .IN2(\SUMB[3][10] ), .QN(n1053) );
  NAND2X0 U1987 ( .IN1(\ab[4][9] ), .IN2(\CARRYB[3][9] ), .QN(n1054) );
  NAND2X0 U1988 ( .IN1(\SUMB[3][10] ), .IN2(\CARRYB[3][9] ), .QN(n1055) );
  NAND3X1 U1989 ( .IN1(n1053), .IN2(n1054), .IN3(n1055), .QN(\CARRYB[4][9] )
         );
  DELLN1X2 U1990 ( .INP(n2206), .Z(n2091) );
  DELLN1X2 U1991 ( .INP(n2228), .Z(n2147) );
  DELLN1X2 U1992 ( .INP(n2213), .Z(n2105) );
  XOR2X1 U1993 ( .IN1(\ab[19][18] ), .IN2(\SUMB[18][19] ), .Q(n1056) );
  NAND2X0 U1994 ( .IN1(\CARRYB[18][18] ), .IN2(\SUMB[18][19] ), .QN(n1057) );
  NAND2X0 U1995 ( .IN1(\CARRYB[18][18] ), .IN2(\ab[19][18] ), .QN(n1058) );
  NAND2X1 U1996 ( .IN1(\SUMB[18][19] ), .IN2(\ab[19][18] ), .QN(n1059) );
  NAND3X1 U1997 ( .IN1(n1057), .IN2(n1058), .IN3(n1059), .QN(\CARRYB[19][18] )
         );
  NAND2X0 U1998 ( .IN1(\ab[20][17] ), .IN2(\SUMB[19][18] ), .QN(n1662) );
  XOR3X1 U1999 ( .IN1(\ab[8][11] ), .IN2(\SUMB[7][12] ), .IN3(\CARRYB[7][11] ), 
        .Q(\SUMB[8][11] ) );
  NAND2X1 U2000 ( .IN1(\ab[8][11] ), .IN2(\SUMB[7][12] ), .QN(n1060) );
  NAND2X0 U2001 ( .IN1(\ab[8][11] ), .IN2(\CARRYB[7][11] ), .QN(n1061) );
  NAND2X0 U2002 ( .IN1(\SUMB[7][12] ), .IN2(\CARRYB[7][11] ), .QN(n1062) );
  NAND3X1 U2003 ( .IN1(n1060), .IN2(n1061), .IN3(n1062), .QN(\CARRYB[8][11] )
         );
  NAND2X0 U2004 ( .IN1(\ab[9][11] ), .IN2(\SUMB[8][12] ), .QN(n1063) );
  NAND2X0 U2005 ( .IN1(\ab[9][11] ), .IN2(\CARRYB[8][11] ), .QN(n1064) );
  NAND2X0 U2006 ( .IN1(\SUMB[8][12] ), .IN2(\CARRYB[8][11] ), .QN(n1065) );
  XOR3X1 U2007 ( .IN1(\ab[21][10] ), .IN2(\CARRYB[20][10] ), .IN3(
        \SUMB[20][11] ), .Q(\SUMB[21][10] ) );
  XOR2X1 U2008 ( .IN1(\ab[22][9] ), .IN2(\CARRYB[21][9] ), .Q(n1066) );
  XOR2X2 U2009 ( .IN1(n1066), .IN2(\SUMB[21][10] ), .Q(\SUMB[22][9] ) );
  NAND2X0 U2010 ( .IN1(\ab[21][10] ), .IN2(\CARRYB[20][10] ), .QN(n1067) );
  NAND2X0 U2011 ( .IN1(\ab[21][10] ), .IN2(\SUMB[20][11] ), .QN(n1068) );
  NAND2X0 U2012 ( .IN1(\CARRYB[20][10] ), .IN2(\SUMB[20][11] ), .QN(n1069) );
  NAND2X0 U2013 ( .IN1(\ab[22][9] ), .IN2(\CARRYB[21][9] ), .QN(n1070) );
  NAND2X0 U2014 ( .IN1(\ab[22][9] ), .IN2(\SUMB[21][10] ), .QN(n1071) );
  NAND2X0 U2015 ( .IN1(\CARRYB[21][9] ), .IN2(\SUMB[21][10] ), .QN(n1072) );
  NAND2X0 U2016 ( .IN1(\CARRYB[2][11] ), .IN2(\ab[3][11] ), .QN(n1073) );
  NAND2X0 U2017 ( .IN1(\CARRYB[2][11] ), .IN2(\SUMB[2][12] ), .QN(n1074) );
  NAND2X0 U2018 ( .IN1(\ab[3][11] ), .IN2(\SUMB[2][12] ), .QN(n1075) );
  NAND3X1 U2019 ( .IN1(n1073), .IN2(n1074), .IN3(n1075), .QN(\CARRYB[3][11] )
         );
  XOR2X1 U2020 ( .IN1(n1076), .IN2(\CARRYB[3][11] ), .Q(\SUMB[4][11] ) );
  NAND2X0 U2021 ( .IN1(\ab[4][11] ), .IN2(\SUMB[3][12] ), .QN(n1077) );
  NAND2X0 U2022 ( .IN1(\ab[4][11] ), .IN2(\CARRYB[3][11] ), .QN(n1078) );
  NAND2X0 U2023 ( .IN1(\SUMB[3][12] ), .IN2(\CARRYB[3][11] ), .QN(n1079) );
  NAND3X1 U2024 ( .IN1(n1077), .IN2(n1078), .IN3(n1079), .QN(\CARRYB[4][11] )
         );
  XOR3X1 U2025 ( .IN1(\ab[23][22] ), .IN2(\CARRYB[22][22] ), .IN3(
        \SUMB[22][23] ), .Q(\SUMB[23][22] ) );
  NAND2X1 U2026 ( .IN1(\ab[23][22] ), .IN2(\CARRYB[22][22] ), .QN(n1080) );
  NAND2X0 U2027 ( .IN1(\ab[23][22] ), .IN2(\SUMB[22][23] ), .QN(n1081) );
  NAND2X0 U2028 ( .IN1(\CARRYB[22][22] ), .IN2(\SUMB[22][23] ), .QN(n1082) );
  NAND2X0 U2029 ( .IN1(\ab[24][21] ), .IN2(\CARRYB[23][21] ), .QN(n1083) );
  NAND2X0 U2030 ( .IN1(\ab[24][21] ), .IN2(\SUMB[23][22] ), .QN(n1084) );
  NAND2X0 U2031 ( .IN1(\CARRYB[23][21] ), .IN2(\SUMB[23][22] ), .QN(n1085) );
  XOR3X1 U2032 ( .IN1(\ab[20][21] ), .IN2(\CARRYB[19][21] ), .IN3(
        \SUMB[19][22] ), .Q(\SUMB[20][21] ) );
  NAND2X1 U2033 ( .IN1(\ab[20][21] ), .IN2(\CARRYB[19][21] ), .QN(n1086) );
  NAND2X0 U2034 ( .IN1(\ab[20][21] ), .IN2(\SUMB[19][22] ), .QN(n1087) );
  NAND2X0 U2035 ( .IN1(\CARRYB[19][21] ), .IN2(\SUMB[19][22] ), .QN(n1088) );
  NAND2X0 U2036 ( .IN1(\ab[21][21] ), .IN2(\SUMB[20][22] ), .QN(n1089) );
  NAND2X0 U2037 ( .IN1(\ab[21][21] ), .IN2(\CARRYB[20][21] ), .QN(n1090) );
  NAND2X0 U2038 ( .IN1(\SUMB[20][22] ), .IN2(\CARRYB[20][21] ), .QN(n1091) );
  XOR3X1 U2039 ( .IN1(\ab[22][14] ), .IN2(\CARRYB[21][14] ), .IN3(
        \SUMB[21][15] ), .Q(\SUMB[22][14] ) );
  NAND2X0 U2040 ( .IN1(\ab[22][14] ), .IN2(\CARRYB[21][14] ), .QN(n1092) );
  NAND2X1 U2041 ( .IN1(\ab[22][14] ), .IN2(\SUMB[21][15] ), .QN(n1093) );
  NAND2X0 U2042 ( .IN1(\CARRYB[21][14] ), .IN2(\SUMB[21][15] ), .QN(n1094) );
  XOR2X1 U2043 ( .IN1(\ab[23][14] ), .IN2(\SUMB[22][15] ), .Q(n1095) );
  NAND2X0 U2044 ( .IN1(\ab[23][14] ), .IN2(\SUMB[22][15] ), .QN(n1096) );
  NAND2X0 U2045 ( .IN1(\ab[23][14] ), .IN2(\CARRYB[22][14] ), .QN(n1097) );
  NAND2X0 U2046 ( .IN1(\SUMB[22][15] ), .IN2(\CARRYB[22][14] ), .QN(n1098) );
  XOR3X1 U2047 ( .IN1(\CARRYB[23][14] ), .IN2(\ab[24][14] ), .IN3(
        \SUMB[23][15] ), .Q(\SUMB[24][14] ) );
  NAND2X1 U2048 ( .IN1(\CARRYB[23][14] ), .IN2(\ab[24][14] ), .QN(n1099) );
  NAND2X0 U2049 ( .IN1(\CARRYB[23][14] ), .IN2(\SUMB[23][15] ), .QN(n1100) );
  NAND2X0 U2050 ( .IN1(\ab[24][14] ), .IN2(\SUMB[23][15] ), .QN(n1101) );
  XOR2X1 U2051 ( .IN1(\ab[25][14] ), .IN2(\SUMB[24][15] ), .Q(n1102) );
  NAND2X0 U2052 ( .IN1(\ab[25][14] ), .IN2(\SUMB[24][15] ), .QN(n1103) );
  NAND2X0 U2053 ( .IN1(\ab[25][14] ), .IN2(\CARRYB[24][14] ), .QN(n1104) );
  NAND2X0 U2054 ( .IN1(\SUMB[24][15] ), .IN2(\CARRYB[24][14] ), .QN(n1105) );
  NAND2X0 U2055 ( .IN1(\ab[10][15] ), .IN2(\CARRYB[9][15] ), .QN(n1106) );
  NAND2X0 U2056 ( .IN1(\ab[10][15] ), .IN2(\SUMB[9][16] ), .QN(n1107) );
  NAND2X0 U2057 ( .IN1(\CARRYB[9][15] ), .IN2(\SUMB[9][16] ), .QN(n1108) );
  NAND3X1 U2058 ( .IN1(n1106), .IN2(n1107), .IN3(n1108), .QN(\CARRYB[10][15] )
         );
  XOR2X1 U2059 ( .IN1(\ab[11][15] ), .IN2(\SUMB[10][16] ), .Q(n1109) );
  XOR2X2 U2060 ( .IN1(n1109), .IN2(\CARRYB[10][15] ), .Q(\SUMB[11][15] ) );
  NAND2X0 U2061 ( .IN1(\ab[11][15] ), .IN2(\SUMB[10][16] ), .QN(n1110) );
  NAND2X0 U2062 ( .IN1(\ab[11][15] ), .IN2(\CARRYB[10][15] ), .QN(n1111) );
  NAND2X0 U2063 ( .IN1(\SUMB[10][16] ), .IN2(\CARRYB[10][15] ), .QN(n1112) );
  XOR3X1 U2064 ( .IN1(\CARRYB[8][15] ), .IN2(\ab[9][15] ), .IN3(\SUMB[8][16] ), 
        .Q(\SUMB[9][15] ) );
  NAND2X0 U2065 ( .IN1(\CARRYB[8][15] ), .IN2(\SUMB[8][16] ), .QN(n1113) );
  NAND2X0 U2066 ( .IN1(\CARRYB[8][15] ), .IN2(\ab[9][15] ), .QN(n1114) );
  NAND2X0 U2067 ( .IN1(\SUMB[8][16] ), .IN2(\ab[9][15] ), .QN(n1115) );
  NAND3X1 U2068 ( .IN1(n1113), .IN2(n1114), .IN3(n1115), .QN(\CARRYB[9][15] )
         );
  XOR3X1 U2069 ( .IN1(\ab[27][27] ), .IN2(\CARRYB[26][27] ), .IN3(
        \SUMB[26][28] ), .Q(\SUMB[27][27] ) );
  XOR2X1 U2070 ( .IN1(\ab[28][26] ), .IN2(\CARRYB[27][26] ), .Q(n1116) );
  NAND2X0 U2071 ( .IN1(\ab[27][27] ), .IN2(\CARRYB[26][27] ), .QN(n1117) );
  NAND2X1 U2072 ( .IN1(\ab[27][27] ), .IN2(\SUMB[26][28] ), .QN(n1118) );
  NAND2X0 U2073 ( .IN1(\CARRYB[26][27] ), .IN2(\SUMB[26][28] ), .QN(n1119) );
  NAND2X0 U2074 ( .IN1(\ab[28][26] ), .IN2(\CARRYB[27][26] ), .QN(n1120) );
  NAND2X0 U2075 ( .IN1(\ab[28][26] ), .IN2(\SUMB[27][27] ), .QN(n1121) );
  NAND2X0 U2076 ( .IN1(\CARRYB[27][26] ), .IN2(\SUMB[27][27] ), .QN(n1122) );
  NAND3X1 U2077 ( .IN1(n1120), .IN2(n1121), .IN3(n1122), .QN(\CARRYB[28][26] )
         );
  XOR3X1 U2078 ( .IN1(\ab[18][4] ), .IN2(\CARRYB[17][4] ), .IN3(\SUMB[17][5] ), 
        .Q(\SUMB[18][4] ) );
  XOR2X1 U2079 ( .IN1(\ab[19][3] ), .IN2(\CARRYB[18][3] ), .Q(n1124) );
  XOR2X2 U2080 ( .IN1(n1124), .IN2(\SUMB[18][4] ), .Q(\SUMB[19][3] ) );
  NAND2X0 U2081 ( .IN1(\ab[18][4] ), .IN2(\SUMB[17][5] ), .QN(n1126) );
  NAND2X0 U2082 ( .IN1(\CARRYB[17][4] ), .IN2(\SUMB[17][5] ), .QN(n1127) );
  NAND3X1 U2083 ( .IN1(n1125), .IN2(n1126), .IN3(n1127), .QN(\CARRYB[18][4] )
         );
  NAND2X0 U2084 ( .IN1(\ab[19][3] ), .IN2(\CARRYB[18][3] ), .QN(n1128) );
  NAND2X0 U2085 ( .IN1(\ab[19][3] ), .IN2(\SUMB[18][4] ), .QN(n1129) );
  NAND2X0 U2086 ( .IN1(\CARRYB[18][3] ), .IN2(\SUMB[18][4] ), .QN(n1130) );
  XOR3X1 U2087 ( .IN1(\ab[22][2] ), .IN2(\CARRYB[21][2] ), .IN3(\SUMB[21][3] ), 
        .Q(\SUMB[22][2] ) );
  XOR2X1 U2088 ( .IN1(\ab[23][1] ), .IN2(\CARRYB[22][1] ), .Q(n1131) );
  XOR2X2 U2089 ( .IN1(n1131), .IN2(\SUMB[22][2] ), .Q(\SUMB[23][1] ) );
  NAND2X0 U2090 ( .IN1(\ab[22][2] ), .IN2(\SUMB[21][3] ), .QN(n1133) );
  NAND2X0 U2091 ( .IN1(\CARRYB[21][2] ), .IN2(\SUMB[21][3] ), .QN(n1134) );
  NAND2X0 U2092 ( .IN1(\ab[23][1] ), .IN2(\CARRYB[22][1] ), .QN(n1135) );
  NAND2X0 U2093 ( .IN1(\ab[23][1] ), .IN2(\SUMB[22][2] ), .QN(n1136) );
  NAND2X0 U2094 ( .IN1(\CARRYB[22][1] ), .IN2(\SUMB[22][2] ), .QN(n1137) );
  XOR3X1 U2095 ( .IN1(\CARRYB[4][7] ), .IN2(\ab[5][7] ), .IN3(\SUMB[4][8] ), 
        .Q(\SUMB[5][7] ) );
  NAND2X0 U2096 ( .IN1(\CARRYB[4][7] ), .IN2(\SUMB[4][8] ), .QN(n1138) );
  NAND2X0 U2097 ( .IN1(\CARRYB[4][7] ), .IN2(\ab[5][7] ), .QN(n1139) );
  NAND2X1 U2098 ( .IN1(\SUMB[4][8] ), .IN2(\ab[5][7] ), .QN(n1140) );
  XOR3X1 U2099 ( .IN1(\ab[6][7] ), .IN2(\CARRYB[5][7] ), .IN3(\SUMB[5][8] ), 
        .Q(\SUMB[6][7] ) );
  NAND2X1 U2100 ( .IN1(\ab[6][7] ), .IN2(\CARRYB[5][7] ), .QN(n1141) );
  NAND2X0 U2101 ( .IN1(\ab[6][7] ), .IN2(\SUMB[5][8] ), .QN(n1142) );
  NAND2X0 U2102 ( .IN1(\CARRYB[5][7] ), .IN2(\SUMB[5][8] ), .QN(n1143) );
  NAND3X1 U2103 ( .IN1(n1141), .IN2(n1142), .IN3(n1143), .QN(\CARRYB[6][7] )
         );
  NAND2X0 U2104 ( .IN1(\ab[7][7] ), .IN2(\SUMB[6][8] ), .QN(n1144) );
  NAND2X0 U2105 ( .IN1(\ab[7][7] ), .IN2(\CARRYB[6][7] ), .QN(n1145) );
  NAND2X0 U2106 ( .IN1(\SUMB[6][8] ), .IN2(\CARRYB[6][7] ), .QN(n1146) );
  XOR3X1 U2107 ( .IN1(\ab[26][19] ), .IN2(\CARRYB[25][19] ), .IN3(
        \SUMB[25][20] ), .Q(\SUMB[26][19] ) );
  NAND2X0 U2108 ( .IN1(\ab[26][19] ), .IN2(\CARRYB[25][19] ), .QN(n1147) );
  NAND2X1 U2109 ( .IN1(\ab[26][19] ), .IN2(\SUMB[25][20] ), .QN(n1148) );
  NAND2X0 U2110 ( .IN1(\CARRYB[25][19] ), .IN2(\SUMB[25][20] ), .QN(n1149) );
  XOR2X1 U2111 ( .IN1(\ab[27][19] ), .IN2(\SUMB[26][20] ), .Q(n1150) );
  XOR2X2 U2112 ( .IN1(n1150), .IN2(\CARRYB[26][19] ), .Q(\SUMB[27][19] ) );
  NAND2X0 U2113 ( .IN1(\ab[27][19] ), .IN2(\SUMB[26][20] ), .QN(n1151) );
  NAND2X0 U2114 ( .IN1(\ab[27][19] ), .IN2(\CARRYB[26][19] ), .QN(n1152) );
  NAND2X0 U2115 ( .IN1(\SUMB[26][20] ), .IN2(\CARRYB[26][19] ), .QN(n1153) );
  XOR3X1 U2116 ( .IN1(\SUMB[18][20] ), .IN2(\ab[19][19] ), .IN3(
        \CARRYB[18][19] ), .Q(\SUMB[19][19] ) );
  NAND2X0 U2117 ( .IN1(\SUMB[18][20] ), .IN2(\ab[19][19] ), .QN(n1154) );
  NAND2X0 U2118 ( .IN1(\SUMB[18][20] ), .IN2(\CARRYB[18][19] ), .QN(n1155) );
  NAND3X1 U2119 ( .IN1(n1154), .IN2(n1155), .IN3(n1156), .QN(\CARRYB[19][19] )
         );
  XOR2X1 U2120 ( .IN1(\ab[20][19] ), .IN2(\SUMB[19][20] ), .Q(n1157) );
  NAND2X0 U2121 ( .IN1(\ab[20][19] ), .IN2(\SUMB[19][20] ), .QN(n1158) );
  NAND2X0 U2122 ( .IN1(\ab[20][19] ), .IN2(\CARRYB[19][19] ), .QN(n1159) );
  NAND2X0 U2123 ( .IN1(\SUMB[19][20] ), .IN2(\CARRYB[19][19] ), .QN(n1160) );
  XOR3X1 U2124 ( .IN1(\CARRYB[14][22] ), .IN2(\ab[15][22] ), .IN3(
        \SUMB[14][23] ), .Q(\SUMB[15][22] ) );
  NAND2X0 U2125 ( .IN1(\CARRYB[14][22] ), .IN2(\SUMB[14][23] ), .QN(n1161) );
  NAND2X0 U2126 ( .IN1(\SUMB[14][23] ), .IN2(\ab[15][22] ), .QN(n1163) );
  XNOR2X2 U2127 ( .IN1(n1164), .IN2(\CARRYB[19][2] ), .Q(\SUMB[20][2] ) );
  XNOR2X1 U2128 ( .IN1(\ab[20][2] ), .IN2(\SUMB[19][3] ), .Q(n1164) );
  NAND2X0 U2129 ( .IN1(\CARRYB[30][10] ), .IN2(\SUMB[30][11] ), .QN(n1165) );
  NAND2X0 U2130 ( .IN1(\CARRYB[30][10] ), .IN2(\ab[31][10] ), .QN(n1166) );
  NAND2X1 U2131 ( .IN1(\SUMB[30][11] ), .IN2(\ab[31][10] ), .QN(n1167) );
  NAND3X1 U2132 ( .IN1(n1165), .IN2(n1166), .IN3(n1167), .QN(\CARRYB[31][10] )
         );
  XOR3X1 U2133 ( .IN1(\ab[8][14] ), .IN2(\CARRYB[7][14] ), .IN3(\SUMB[7][15] ), 
        .Q(\SUMB[8][14] ) );
  NAND2X1 U2134 ( .IN1(\ab[8][14] ), .IN2(\CARRYB[7][14] ), .QN(n1168) );
  NAND2X0 U2135 ( .IN1(\ab[8][14] ), .IN2(\SUMB[7][15] ), .QN(n1169) );
  NAND2X0 U2136 ( .IN1(\CARRYB[7][14] ), .IN2(\SUMB[7][15] ), .QN(n1170) );
  XOR2X1 U2137 ( .IN1(\ab[9][14] ), .IN2(\SUMB[8][15] ), .Q(n1171) );
  XOR2X2 U2138 ( .IN1(n1171), .IN2(\CARRYB[8][14] ), .Q(\SUMB[9][14] ) );
  NAND2X0 U2139 ( .IN1(\ab[9][14] ), .IN2(\SUMB[8][15] ), .QN(n1172) );
  NAND2X0 U2140 ( .IN1(\ab[9][14] ), .IN2(\CARRYB[8][14] ), .QN(n1173) );
  NAND2X0 U2141 ( .IN1(\SUMB[8][15] ), .IN2(\CARRYB[8][14] ), .QN(n1174) );
  NAND3X1 U2142 ( .IN1(n1172), .IN2(n1173), .IN3(n1174), .QN(\CARRYB[9][14] )
         );
  XOR3X1 U2143 ( .IN1(\CARRYB[29][10] ), .IN2(\ab[30][10] ), .IN3(
        \SUMB[29][11] ), .Q(\SUMB[30][10] ) );
  NAND2X0 U2144 ( .IN1(\CARRYB[29][10] ), .IN2(\SUMB[29][11] ), .QN(n1175) );
  NAND2X0 U2145 ( .IN1(\CARRYB[29][10] ), .IN2(\ab[30][10] ), .QN(n1176) );
  NAND2X0 U2146 ( .IN1(\SUMB[29][11] ), .IN2(\ab[30][10] ), .QN(n1177) );
  NAND3X1 U2147 ( .IN1(n1175), .IN2(n1176), .IN3(n1177), .QN(\CARRYB[30][10] )
         );
  XOR3X1 U2148 ( .IN1(\CARRYB[27][10] ), .IN2(\ab[28][10] ), .IN3(
        \SUMB[27][11] ), .Q(\SUMB[28][10] ) );
  NAND2X0 U2149 ( .IN1(\CARRYB[27][10] ), .IN2(\SUMB[27][11] ), .QN(n1178) );
  NAND2X1 U2150 ( .IN1(\CARRYB[27][10] ), .IN2(\ab[28][10] ), .QN(n1179) );
  NAND2X0 U2151 ( .IN1(\SUMB[27][11] ), .IN2(\ab[28][10] ), .QN(n1180) );
  NAND3X0 U2152 ( .IN1(n1178), .IN2(n1179), .IN3(n1180), .QN(\CARRYB[28][10] )
         );
  NAND2X1 U2153 ( .IN1(\CARRYB[15][21] ), .IN2(\ab[16][21] ), .QN(n1181) );
  NAND2X0 U2154 ( .IN1(\CARRYB[15][21] ), .IN2(\SUMB[15][22] ), .QN(n1182) );
  NAND2X0 U2155 ( .IN1(\ab[16][21] ), .IN2(\SUMB[15][22] ), .QN(n1183) );
  XOR2X1 U2156 ( .IN1(\ab[17][21] ), .IN2(\SUMB[16][22] ), .Q(n1184) );
  XOR2X2 U2157 ( .IN1(n1184), .IN2(\CARRYB[16][21] ), .Q(\SUMB[17][21] ) );
  NAND2X0 U2158 ( .IN1(\ab[17][21] ), .IN2(\SUMB[16][22] ), .QN(n1185) );
  NAND2X0 U2159 ( .IN1(\ab[17][21] ), .IN2(\CARRYB[16][21] ), .QN(n1186) );
  NAND2X0 U2160 ( .IN1(\SUMB[16][22] ), .IN2(\CARRYB[16][21] ), .QN(n1187) );
  XOR3X1 U2161 ( .IN1(\ab[4][21] ), .IN2(\CARRYB[3][21] ), .IN3(\SUMB[3][22] ), 
        .Q(\SUMB[4][21] ) );
  NAND2X0 U2162 ( .IN1(\ab[4][21] ), .IN2(\SUMB[3][22] ), .QN(n1189) );
  NAND2X0 U2163 ( .IN1(\CARRYB[3][21] ), .IN2(\SUMB[3][22] ), .QN(n1190) );
  NAND2X0 U2164 ( .IN1(\ab[5][21] ), .IN2(\SUMB[4][22] ), .QN(n1191) );
  NAND2X0 U2165 ( .IN1(\ab[5][21] ), .IN2(\CARRYB[4][21] ), .QN(n1192) );
  NAND2X0 U2166 ( .IN1(\SUMB[4][22] ), .IN2(\CARRYB[4][21] ), .QN(n1193) );
  NAND3X1 U2167 ( .IN1(n1191), .IN2(n1192), .IN3(n1193), .QN(\CARRYB[5][21] )
         );
  XOR3X1 U2168 ( .IN1(\CARRYB[17][2] ), .IN2(\ab[18][2] ), .IN3(\SUMB[17][3] ), 
        .Q(\SUMB[18][2] ) );
  NAND2X0 U2169 ( .IN1(\CARRYB[17][2] ), .IN2(\SUMB[17][3] ), .QN(n1194) );
  NAND2X0 U2170 ( .IN1(\CARRYB[17][2] ), .IN2(\ab[18][2] ), .QN(n1195) );
  NAND2X1 U2171 ( .IN1(\SUMB[17][3] ), .IN2(\ab[18][2] ), .QN(n1196) );
  NAND3X0 U2172 ( .IN1(n1194), .IN2(n1195), .IN3(n1196), .QN(\CARRYB[18][2] )
         );
  XOR3X1 U2173 ( .IN1(\ab[3][4] ), .IN2(\CARRYB[2][4] ), .IN3(\SUMB[2][5] ), 
        .Q(\SUMB[3][4] ) );
  NAND2X1 U2174 ( .IN1(\ab[3][4] ), .IN2(\CARRYB[2][4] ), .QN(n1197) );
  NAND2X0 U2175 ( .IN1(\ab[3][4] ), .IN2(\SUMB[2][5] ), .QN(n1198) );
  NAND2X0 U2176 ( .IN1(\CARRYB[2][4] ), .IN2(\SUMB[2][5] ), .QN(n1199) );
  XOR2X1 U2177 ( .IN1(\ab[4][4] ), .IN2(\SUMB[3][5] ), .Q(n1200) );
  NAND2X0 U2178 ( .IN1(\ab[4][4] ), .IN2(\SUMB[3][5] ), .QN(n1201) );
  NAND2X0 U2179 ( .IN1(\ab[4][4] ), .IN2(\CARRYB[3][4] ), .QN(n1202) );
  NAND2X0 U2180 ( .IN1(\SUMB[3][5] ), .IN2(\CARRYB[3][4] ), .QN(n1203) );
  XOR3X1 U2181 ( .IN1(\ab[19][2] ), .IN2(\CARRYB[18][2] ), .IN3(\SUMB[18][3] ), 
        .Q(\SUMB[19][2] ) );
  NAND2X1 U2182 ( .IN1(\ab[19][2] ), .IN2(\CARRYB[18][2] ), .QN(n1204) );
  NAND2X0 U2183 ( .IN1(\ab[19][2] ), .IN2(\SUMB[18][3] ), .QN(n1205) );
  NAND2X0 U2184 ( .IN1(\CARRYB[18][2] ), .IN2(\SUMB[18][3] ), .QN(n1206) );
  NAND2X0 U2185 ( .IN1(\ab[20][2] ), .IN2(\SUMB[19][3] ), .QN(n1207) );
  NAND2X0 U2186 ( .IN1(\ab[20][2] ), .IN2(\CARRYB[19][2] ), .QN(n1208) );
  NAND2X0 U2187 ( .IN1(\SUMB[19][3] ), .IN2(\CARRYB[19][2] ), .QN(n1209) );
  XOR3X1 U2188 ( .IN1(\CARRYB[16][2] ), .IN2(\ab[17][2] ), .IN3(\SUMB[16][3] ), 
        .Q(\SUMB[17][2] ) );
  NAND2X0 U2189 ( .IN1(\CARRYB[16][2] ), .IN2(\SUMB[16][3] ), .QN(n1210) );
  NAND2X1 U2190 ( .IN1(\CARRYB[16][2] ), .IN2(\ab[17][2] ), .QN(n1211) );
  NAND2X0 U2191 ( .IN1(\SUMB[16][3] ), .IN2(\ab[17][2] ), .QN(n1212) );
  NAND3X0 U2192 ( .IN1(n1942), .IN2(n1943), .IN3(n1944), .QN(\CARRYB[16][2] )
         );
  DELLN1X2 U2193 ( .INP(n2216), .Z(n2114) );
  NBUFFX4 U2194 ( .INP(n2218), .Z(n2119) );
  DELLN1X2 U2195 ( .INP(n2218), .Z(n2121) );
  XOR3X1 U2196 ( .IN1(\ab[18][7] ), .IN2(\CARRYB[17][7] ), .IN3(\SUMB[17][8] ), 
        .Q(\SUMB[18][7] ) );
  NAND2X0 U2197 ( .IN1(\ab[18][7] ), .IN2(\CARRYB[17][7] ), .QN(n1213) );
  NAND2X0 U2198 ( .IN1(\ab[18][7] ), .IN2(\SUMB[17][8] ), .QN(n1214) );
  NAND2X0 U2199 ( .IN1(\CARRYB[17][7] ), .IN2(\SUMB[17][8] ), .QN(n1215) );
  NAND2X0 U2200 ( .IN1(\ab[19][6] ), .IN2(\CARRYB[18][6] ), .QN(n1216) );
  NAND2X0 U2201 ( .IN1(\ab[19][6] ), .IN2(\SUMB[18][7] ), .QN(n1217) );
  NAND2X0 U2202 ( .IN1(\CARRYB[18][6] ), .IN2(\SUMB[18][7] ), .QN(n1218) );
  XOR3X1 U2203 ( .IN1(\ab[2][8] ), .IN2(n1354), .IN3(\SUMB[1][9] ), .Q(
        \SUMB[2][8] ) );
  NAND2X1 U2204 ( .IN1(\ab[2][8] ), .IN2(n1354), .QN(n1219) );
  NAND2X0 U2205 ( .IN1(\ab[2][8] ), .IN2(\SUMB[1][9] ), .QN(n1220) );
  NAND2X0 U2206 ( .IN1(n1354), .IN2(\SUMB[1][9] ), .QN(n1221) );
  XOR2X1 U2207 ( .IN1(\ab[3][8] ), .IN2(\SUMB[2][9] ), .Q(n1222) );
  NAND2X0 U2208 ( .IN1(\ab[3][8] ), .IN2(\SUMB[2][9] ), .QN(n1223) );
  NAND2X0 U2209 ( .IN1(\ab[3][8] ), .IN2(\CARRYB[2][8] ), .QN(n1224) );
  NAND2X0 U2210 ( .IN1(\SUMB[2][9] ), .IN2(\CARRYB[2][8] ), .QN(n1225) );
  XOR2X2 U2211 ( .IN1(\CARRYB[31][1] ), .IN2(\SUMB[31][2] ), .Q(\A1[31] ) );
  DELLN1X2 U2212 ( .INP(n2231), .Z(n2157) );
  DELLN1X2 U2213 ( .INP(n2228), .Z(n2148) );
  XOR2X1 U2214 ( .IN1(\ab[31][11] ), .IN2(\SUMB[30][12] ), .Q(n1226) );
  XOR2X1 U2215 ( .IN1(n1226), .IN2(\CARRYB[30][11] ), .Q(\SUMB[31][11] ) );
  NAND2X0 U2216 ( .IN1(\CARRYB[30][11] ), .IN2(\SUMB[30][12] ), .QN(n1227) );
  NAND2X0 U2217 ( .IN1(\CARRYB[30][11] ), .IN2(\ab[31][11] ), .QN(n1228) );
  NAND2X1 U2218 ( .IN1(\SUMB[30][12] ), .IN2(\ab[31][11] ), .QN(n1229) );
  NAND2X0 U2219 ( .IN1(\ab[10][17] ), .IN2(\CARRYB[9][17] ), .QN(n1230) );
  NAND2X1 U2220 ( .IN1(\ab[10][17] ), .IN2(\SUMB[9][18] ), .QN(n1231) );
  NAND2X0 U2221 ( .IN1(\CARRYB[9][17] ), .IN2(\SUMB[9][18] ), .QN(n1232) );
  NAND3X1 U2222 ( .IN1(n1230), .IN2(n1231), .IN3(n1232), .QN(\CARRYB[10][17] )
         );
  XOR2X1 U2223 ( .IN1(\ab[11][17] ), .IN2(\SUMB[10][18] ), .Q(n1233) );
  NAND2X0 U2224 ( .IN1(\ab[11][17] ), .IN2(\SUMB[10][18] ), .QN(n1234) );
  NAND2X0 U2225 ( .IN1(\ab[11][17] ), .IN2(\CARRYB[10][17] ), .QN(n1235) );
  NAND2X0 U2226 ( .IN1(\SUMB[10][18] ), .IN2(\CARRYB[10][17] ), .QN(n1236) );
  NAND3X1 U2227 ( .IN1(n1234), .IN2(n1235), .IN3(n1236), .QN(\CARRYB[11][17] )
         );
  XOR3X1 U2228 ( .IN1(\ab[7][17] ), .IN2(\CARRYB[6][17] ), .IN3(\SUMB[6][18] ), 
        .Q(\SUMB[7][17] ) );
  NAND2X0 U2229 ( .IN1(\ab[7][17] ), .IN2(\CARRYB[6][17] ), .QN(n1237) );
  NAND2X1 U2230 ( .IN1(\ab[7][17] ), .IN2(\SUMB[6][18] ), .QN(n1238) );
  NAND2X0 U2231 ( .IN1(\CARRYB[6][17] ), .IN2(\SUMB[6][18] ), .QN(n1239) );
  NAND3X1 U2232 ( .IN1(n1237), .IN2(n1238), .IN3(n1239), .QN(\CARRYB[7][17] )
         );
  XOR2X1 U2233 ( .IN1(\ab[8][17] ), .IN2(\SUMB[7][18] ), .Q(n1240) );
  NAND2X0 U2234 ( .IN1(\ab[8][17] ), .IN2(\SUMB[7][18] ), .QN(n1241) );
  NAND2X0 U2235 ( .IN1(\ab[8][17] ), .IN2(\CARRYB[7][17] ), .QN(n1242) );
  NAND2X0 U2236 ( .IN1(\SUMB[7][18] ), .IN2(\CARRYB[7][17] ), .QN(n1243) );
  XOR3X1 U2237 ( .IN1(\ab[21][15] ), .IN2(\CARRYB[20][15] ), .IN3(
        \SUMB[20][16] ), .Q(\SUMB[21][15] ) );
  NAND2X0 U2238 ( .IN1(\ab[21][15] ), .IN2(\CARRYB[20][15] ), .QN(n1244) );
  NAND2X0 U2239 ( .IN1(\ab[21][15] ), .IN2(\SUMB[20][16] ), .QN(n1245) );
  NAND2X0 U2240 ( .IN1(\CARRYB[20][15] ), .IN2(\SUMB[20][16] ), .QN(n1246) );
  XOR2X1 U2241 ( .IN1(\ab[22][15] ), .IN2(\SUMB[21][16] ), .Q(n1247) );
  XOR2X2 U2242 ( .IN1(n1247), .IN2(\CARRYB[21][15] ), .Q(\SUMB[22][15] ) );
  NAND2X0 U2243 ( .IN1(\ab[22][15] ), .IN2(\SUMB[21][16] ), .QN(n1248) );
  NAND2X0 U2244 ( .IN1(\ab[22][15] ), .IN2(\CARRYB[21][15] ), .QN(n1249) );
  NAND2X0 U2245 ( .IN1(\SUMB[21][16] ), .IN2(\CARRYB[21][15] ), .QN(n1250) );
  XOR3X1 U2246 ( .IN1(\CARRYB[19][15] ), .IN2(\ab[20][15] ), .IN3(
        \SUMB[19][16] ), .Q(\SUMB[20][15] ) );
  NAND2X0 U2247 ( .IN1(\CARRYB[19][15] ), .IN2(\SUMB[19][16] ), .QN(n1251) );
  NAND2X1 U2248 ( .IN1(\CARRYB[19][15] ), .IN2(\ab[20][15] ), .QN(n1252) );
  NAND2X0 U2249 ( .IN1(\SUMB[19][16] ), .IN2(\ab[20][15] ), .QN(n1253) );
  XOR2X1 U2250 ( .IN1(\ab[30][11] ), .IN2(\SUMB[29][12] ), .Q(n1254) );
  XOR2X1 U2251 ( .IN1(n1254), .IN2(\CARRYB[29][11] ), .Q(\SUMB[30][11] ) );
  NAND2X0 U2252 ( .IN1(\CARRYB[29][11] ), .IN2(\SUMB[29][12] ), .QN(n1255) );
  NAND2X0 U2253 ( .IN1(\CARRYB[29][11] ), .IN2(\ab[30][11] ), .QN(n1256) );
  NAND2X1 U2254 ( .IN1(\SUMB[29][12] ), .IN2(\ab[30][11] ), .QN(n1257) );
  NAND3X1 U2255 ( .IN1(n1255), .IN2(n1256), .IN3(n1257), .QN(\CARRYB[30][11] )
         );
  XOR2X1 U2256 ( .IN1(n1886), .IN2(\CARRYB[29][12] ), .Q(\SUMB[30][12] ) );
  XOR2X1 U2257 ( .IN1(\CARRYB[31][11] ), .IN2(\SUMB[31][12] ), .Q(\A1[41] ) );
  XOR3X1 U2258 ( .IN1(\ab[25][15] ), .IN2(\CARRYB[24][15] ), .IN3(
        \SUMB[24][16] ), .Q(\SUMB[25][15] ) );
  NAND2X0 U2259 ( .IN1(\ab[25][15] ), .IN2(\CARRYB[24][15] ), .QN(n1471) );
  NBUFFX4 U2260 ( .INP(n2222), .Z(n2131) );
  NBUFFX4 U2261 ( .INP(n2222), .Z(n2133) );
  NBUFFX4 U2262 ( .INP(n2235), .Z(n2164) );
  NBUFFX4 U2263 ( .INP(n2235), .Z(n2166) );
  NBUFFX4 U2264 ( .INP(n2235), .Z(n2165) );
  NAND2X0 U2265 ( .IN1(\CARRYB[21][12] ), .IN2(\ab[22][12] ), .QN(n1306) );
  XOR3X1 U2266 ( .IN1(\ab[23][29] ), .IN2(\CARRYB[22][29] ), .IN3(
        \SUMB[22][30] ), .Q(\SUMB[23][29] ) );
  XOR2X1 U2267 ( .IN1(\ab[24][28] ), .IN2(\CARRYB[23][28] ), .Q(n1258) );
  NAND2X0 U2268 ( .IN1(\ab[23][29] ), .IN2(\CARRYB[22][29] ), .QN(n1259) );
  NAND2X1 U2269 ( .IN1(\ab[23][29] ), .IN2(\SUMB[22][30] ), .QN(n1260) );
  NAND2X0 U2270 ( .IN1(\CARRYB[22][29] ), .IN2(\SUMB[22][30] ), .QN(n1261) );
  NAND2X0 U2271 ( .IN1(\ab[24][28] ), .IN2(\CARRYB[23][28] ), .QN(n1262) );
  NAND2X0 U2272 ( .IN1(\ab[24][28] ), .IN2(\SUMB[23][29] ), .QN(n1263) );
  NAND2X0 U2273 ( .IN1(\CARRYB[23][28] ), .IN2(\SUMB[23][29] ), .QN(n1264) );
  XOR3X1 U2274 ( .IN1(\ab[21][29] ), .IN2(\CARRYB[20][29] ), .IN3(
        \SUMB[20][30] ), .Q(\SUMB[21][29] ) );
  NAND2X0 U2275 ( .IN1(\ab[21][29] ), .IN2(\CARRYB[20][29] ), .QN(n1265) );
  NAND2X1 U2276 ( .IN1(\ab[21][29] ), .IN2(\SUMB[20][30] ), .QN(n1266) );
  NAND2X0 U2277 ( .IN1(\CARRYB[20][29] ), .IN2(\SUMB[20][30] ), .QN(n1267) );
  XOR2X1 U2278 ( .IN1(\ab[22][29] ), .IN2(\SUMB[21][30] ), .Q(n1268) );
  XOR2X1 U2279 ( .IN1(n1268), .IN2(\CARRYB[21][29] ), .Q(\SUMB[22][29] ) );
  NAND2X0 U2280 ( .IN1(\ab[22][29] ), .IN2(\SUMB[21][30] ), .QN(n1269) );
  NAND2X0 U2281 ( .IN1(\ab[22][29] ), .IN2(\CARRYB[21][29] ), .QN(n1270) );
  NAND2X0 U2282 ( .IN1(\SUMB[21][30] ), .IN2(\CARRYB[21][29] ), .QN(n1271) );
  NBUFFX4 U2283 ( .INP(n2231), .Z(n2155) );
  XOR3X1 U2284 ( .IN1(\SUMB[23][13] ), .IN2(\ab[24][12] ), .IN3(
        \CARRYB[23][12] ), .Q(\SUMB[24][12] ) );
  NAND2X0 U2285 ( .IN1(\SUMB[23][13] ), .IN2(\CARRYB[23][12] ), .QN(n1272) );
  NAND2X0 U2286 ( .IN1(\SUMB[23][13] ), .IN2(\ab[24][12] ), .QN(n1273) );
  NAND2X1 U2287 ( .IN1(\CARRYB[23][12] ), .IN2(\ab[24][12] ), .QN(n1274) );
  NAND3X0 U2288 ( .IN1(n1272), .IN2(n1273), .IN3(n1274), .QN(\CARRYB[24][12] )
         );
  XOR3X1 U2289 ( .IN1(\ab[22][13] ), .IN2(\CARRYB[21][13] ), .IN3(
        \SUMB[21][14] ), .Q(\SUMB[22][13] ) );
  NAND2X1 U2290 ( .IN1(\ab[22][13] ), .IN2(\CARRYB[21][13] ), .QN(n1275) );
  NAND2X0 U2291 ( .IN1(\ab[22][13] ), .IN2(\SUMB[21][14] ), .QN(n1276) );
  NAND2X0 U2292 ( .IN1(\CARRYB[21][13] ), .IN2(\SUMB[21][14] ), .QN(n1277) );
  NAND3X0 U2293 ( .IN1(n1275), .IN2(n1276), .IN3(n1277), .QN(\CARRYB[22][13] )
         );
  XOR2X1 U2294 ( .IN1(\ab[23][13] ), .IN2(\SUMB[22][14] ), .Q(n1278) );
  XOR2X2 U2295 ( .IN1(n1278), .IN2(\CARRYB[22][13] ), .Q(\SUMB[23][13] ) );
  NAND2X0 U2296 ( .IN1(\ab[23][13] ), .IN2(\SUMB[22][14] ), .QN(n1279) );
  NAND2X0 U2297 ( .IN1(\ab[23][13] ), .IN2(\CARRYB[22][13] ), .QN(n1280) );
  NAND2X0 U2298 ( .IN1(\SUMB[22][14] ), .IN2(\CARRYB[22][13] ), .QN(n1281) );
  XOR3X1 U2299 ( .IN1(\ab[21][8] ), .IN2(\CARRYB[20][8] ), .IN3(\SUMB[20][9] ), 
        .Q(\SUMB[21][8] ) );
  XOR2X1 U2300 ( .IN1(\ab[22][7] ), .IN2(\CARRYB[21][7] ), .Q(n1282) );
  NAND2X0 U2301 ( .IN1(\ab[21][8] ), .IN2(\CARRYB[20][8] ), .QN(n1283) );
  NAND2X0 U2302 ( .IN1(\ab[21][8] ), .IN2(\SUMB[20][9] ), .QN(n1284) );
  NAND2X0 U2303 ( .IN1(\CARRYB[20][8] ), .IN2(\SUMB[20][9] ), .QN(n1285) );
  NAND3X1 U2304 ( .IN1(n1283), .IN2(n1284), .IN3(n1285), .QN(\CARRYB[21][8] )
         );
  NAND2X0 U2305 ( .IN1(\ab[22][7] ), .IN2(\CARRYB[21][7] ), .QN(n1286) );
  NAND2X0 U2306 ( .IN1(\ab[22][7] ), .IN2(\SUMB[21][8] ), .QN(n1287) );
  NAND2X0 U2307 ( .IN1(\CARRYB[21][7] ), .IN2(\SUMB[21][8] ), .QN(n1288) );
  XOR3X1 U2308 ( .IN1(\ab[17][9] ), .IN2(\CARRYB[16][9] ), .IN3(\SUMB[16][10] ), .Q(\SUMB[17][9] ) );
  NAND2X0 U2309 ( .IN1(\ab[17][9] ), .IN2(\CARRYB[16][9] ), .QN(n1289) );
  NAND2X1 U2310 ( .IN1(\ab[17][9] ), .IN2(\SUMB[16][10] ), .QN(n1290) );
  NAND2X0 U2311 ( .IN1(\CARRYB[16][9] ), .IN2(\SUMB[16][10] ), .QN(n1291) );
  NAND2X0 U2312 ( .IN1(\ab[18][8] ), .IN2(\CARRYB[17][8] ), .QN(n1292) );
  NAND2X0 U2313 ( .IN1(\ab[18][8] ), .IN2(\SUMB[17][9] ), .QN(n1293) );
  NAND2X0 U2314 ( .IN1(\CARRYB[17][8] ), .IN2(\SUMB[17][9] ), .QN(n1294) );
  XOR3X1 U2315 ( .IN1(\CARRYB[18][8] ), .IN2(\ab[19][8] ), .IN3(\SUMB[18][9] ), 
        .Q(\SUMB[19][8] ) );
  NAND2X0 U2316 ( .IN1(\CARRYB[18][8] ), .IN2(\SUMB[18][9] ), .QN(n1295) );
  NAND2X0 U2317 ( .IN1(\CARRYB[18][8] ), .IN2(\ab[19][8] ), .QN(n1296) );
  XOR3X1 U2318 ( .IN1(\ab[11][9] ), .IN2(\CARRYB[10][9] ), .IN3(\SUMB[10][10] ), .Q(\SUMB[11][9] ) );
  NAND2X0 U2319 ( .IN1(\ab[11][9] ), .IN2(\CARRYB[10][9] ), .QN(n1298) );
  NAND2X0 U2320 ( .IN1(\CARRYB[10][9] ), .IN2(\SUMB[10][10] ), .QN(n1300) );
  NAND2X0 U2321 ( .IN1(\ab[12][9] ), .IN2(\SUMB[11][10] ), .QN(n1301) );
  NAND2X0 U2322 ( .IN1(\ab[12][9] ), .IN2(\CARRYB[11][9] ), .QN(n1302) );
  NAND2X0 U2323 ( .IN1(\CARRYB[11][9] ), .IN2(\SUMB[11][10] ), .QN(n1303) );
  XOR3X1 U2324 ( .IN1(\SUMB[21][13] ), .IN2(\ab[22][12] ), .IN3(
        \CARRYB[21][12] ), .Q(\SUMB[22][12] ) );
  NAND2X0 U2325 ( .IN1(\SUMB[21][13] ), .IN2(\CARRYB[21][12] ), .QN(n1304) );
  NAND2X0 U2326 ( .IN1(\SUMB[21][13] ), .IN2(\ab[22][12] ), .QN(n1305) );
  XOR3X1 U2327 ( .IN1(\SUMB[19][14] ), .IN2(\ab[20][13] ), .IN3(
        \CARRYB[19][13] ), .Q(\SUMB[20][13] ) );
  NAND2X0 U2328 ( .IN1(\SUMB[19][14] ), .IN2(\ab[20][13] ), .QN(n1308) );
  NAND3X0 U2329 ( .IN1(n1307), .IN2(n1308), .IN3(n1309), .QN(\CARRYB[20][13] )
         );
  XOR2X1 U2330 ( .IN1(n1685), .IN2(\CARRYB[18][14] ), .Q(\SUMB[19][14] ) );
  XNOR2X1 U2331 ( .IN1(\ab[19][12] ), .IN2(\SUMB[18][13] ), .Q(n1310) );
  NAND2X0 U2332 ( .IN1(\CARRYB[4][23] ), .IN2(\ab[5][23] ), .QN(n1523) );
  XNOR2X1 U2333 ( .IN1(\ab[30][6] ), .IN2(\SUMB[29][7] ), .Q(n1311) );
  XOR3X1 U2334 ( .IN1(\CARRYB[10][16] ), .IN2(\ab[11][16] ), .IN3(
        \SUMB[10][17] ), .Q(\SUMB[11][16] ) );
  NAND2X0 U2335 ( .IN1(\CARRYB[10][16] ), .IN2(\SUMB[10][17] ), .QN(n1312) );
  NAND2X0 U2336 ( .IN1(\SUMB[10][17] ), .IN2(\ab[11][16] ), .QN(n1314) );
  XOR3X1 U2337 ( .IN1(\CARRYB[16][13] ), .IN2(\ab[17][13] ), .IN3(
        \SUMB[16][14] ), .Q(\SUMB[17][13] ) );
  NAND2X0 U2338 ( .IN1(\CARRYB[16][13] ), .IN2(\SUMB[16][14] ), .QN(n1315) );
  NAND2X0 U2339 ( .IN1(\SUMB[16][14] ), .IN2(\ab[17][13] ), .QN(n1317) );
  NAND3X0 U2340 ( .IN1(n1315), .IN2(n1316), .IN3(n1317), .QN(\CARRYB[17][13] )
         );
  XOR3X1 U2341 ( .IN1(\CARRYB[12][14] ), .IN2(\ab[13][14] ), .IN3(
        \SUMB[12][15] ), .Q(\SUMB[13][14] ) );
  NAND2X0 U2342 ( .IN1(\SUMB[12][15] ), .IN2(\ab[13][14] ), .QN(n1320) );
  NAND3X0 U2343 ( .IN1(n1318), .IN2(n1319), .IN3(n1320), .QN(\CARRYB[13][14] )
         );
  XOR3X1 U2344 ( .IN1(\CARRYB[10][12] ), .IN2(\ab[11][12] ), .IN3(
        \SUMB[10][13] ), .Q(\SUMB[11][12] ) );
  NAND2X0 U2345 ( .IN1(\CARRYB[10][12] ), .IN2(\SUMB[10][13] ), .QN(n1321) );
  NAND2X0 U2346 ( .IN1(\SUMB[10][13] ), .IN2(\ab[11][12] ), .QN(n1323) );
  NAND2X0 U2347 ( .IN1(\ab[9][13] ), .IN2(\CARRYB[8][13] ), .QN(n1324) );
  NAND2X0 U2348 ( .IN1(\ab[9][13] ), .IN2(\SUMB[8][14] ), .QN(n1325) );
  NAND2X0 U2349 ( .IN1(\CARRYB[8][13] ), .IN2(\SUMB[8][14] ), .QN(n1326) );
  NAND2X0 U2350 ( .IN1(\ab[10][12] ), .IN2(\CARRYB[9][12] ), .QN(n1327) );
  NAND2X0 U2351 ( .IN1(\ab[10][12] ), .IN2(\SUMB[9][13] ), .QN(n1328) );
  NAND2X0 U2352 ( .IN1(\CARRYB[9][12] ), .IN2(\SUMB[9][13] ), .QN(n1329) );
  XOR3X1 U2353 ( .IN1(\ab[29][2] ), .IN2(\CARRYB[28][2] ), .IN3(\SUMB[28][3] ), 
        .Q(\SUMB[29][2] ) );
  NAND2X0 U2354 ( .IN1(\ab[29][2] ), .IN2(\CARRYB[28][2] ), .QN(n1330) );
  NAND2X1 U2355 ( .IN1(\ab[29][2] ), .IN2(\SUMB[28][3] ), .QN(n1331) );
  NAND2X0 U2356 ( .IN1(\CARRYB[28][2] ), .IN2(\SUMB[28][3] ), .QN(n1332) );
  NAND3X1 U2357 ( .IN1(n1330), .IN2(n1331), .IN3(n1332), .QN(\CARRYB[29][2] )
         );
  XOR2X1 U2358 ( .IN1(\ab[30][2] ), .IN2(\SUMB[29][3] ), .Q(n1333) );
  NAND2X0 U2359 ( .IN1(\ab[30][2] ), .IN2(\SUMB[29][3] ), .QN(n1334) );
  NAND2X0 U2360 ( .IN1(\ab[30][2] ), .IN2(\CARRYB[29][2] ), .QN(n1335) );
  NAND2X0 U2361 ( .IN1(\SUMB[29][3] ), .IN2(\CARRYB[29][2] ), .QN(n1336) );
  XOR3X1 U2362 ( .IN1(\ab[24][3] ), .IN2(\CARRYB[23][3] ), .IN3(\SUMB[23][4] ), 
        .Q(\SUMB[24][3] ) );
  NAND2X0 U2363 ( .IN1(\ab[24][3] ), .IN2(\CARRYB[23][3] ), .QN(n1337) );
  NAND2X1 U2364 ( .IN1(\ab[24][3] ), .IN2(\SUMB[23][4] ), .QN(n1338) );
  NAND2X0 U2365 ( .IN1(\CARRYB[23][3] ), .IN2(\SUMB[23][4] ), .QN(n1339) );
  NAND2X0 U2366 ( .IN1(\ab[25][3] ), .IN2(\SUMB[24][4] ), .QN(n1340) );
  NAND2X0 U2367 ( .IN1(\ab[25][3] ), .IN2(\CARRYB[24][3] ), .QN(n1341) );
  NAND2X0 U2368 ( .IN1(\SUMB[24][4] ), .IN2(\CARRYB[24][3] ), .QN(n1342) );
  XOR2X1 U2369 ( .IN1(\ab[23][3] ), .IN2(\SUMB[22][4] ), .Q(n1343) );
  XOR2X1 U2370 ( .IN1(n1343), .IN2(\CARRYB[22][3] ), .Q(\SUMB[23][3] ) );
  NAND2X0 U2371 ( .IN1(\CARRYB[22][3] ), .IN2(\SUMB[22][4] ), .QN(n1344) );
  NAND2X0 U2372 ( .IN1(\CARRYB[22][3] ), .IN2(\ab[23][3] ), .QN(n1345) );
  NAND2X1 U2373 ( .IN1(\SUMB[22][4] ), .IN2(\ab[23][3] ), .QN(n1346) );
  XOR3X1 U2374 ( .IN1(\ab[6][6] ), .IN2(\CARRYB[5][6] ), .IN3(\SUMB[5][7] ), 
        .Q(\SUMB[6][6] ) );
  NAND2X0 U2375 ( .IN1(\ab[6][6] ), .IN2(\SUMB[5][7] ), .QN(n1348) );
  NAND2X0 U2376 ( .IN1(\CARRYB[5][6] ), .IN2(\SUMB[5][7] ), .QN(n1349) );
  NAND3X1 U2377 ( .IN1(n1347), .IN2(n1348), .IN3(n1349), .QN(\CARRYB[6][6] )
         );
  XOR2X1 U2378 ( .IN1(\ab[7][6] ), .IN2(\SUMB[6][7] ), .Q(n1350) );
  XOR2X2 U2379 ( .IN1(n1350), .IN2(\CARRYB[6][6] ), .Q(\SUMB[7][6] ) );
  NAND2X0 U2380 ( .IN1(\ab[7][6] ), .IN2(\SUMB[6][7] ), .QN(n1351) );
  NAND2X0 U2381 ( .IN1(\ab[7][6] ), .IN2(\CARRYB[6][6] ), .QN(n1352) );
  NAND2X0 U2382 ( .IN1(\SUMB[6][7] ), .IN2(\CARRYB[6][6] ), .QN(n1353) );
  NAND3X1 U2383 ( .IN1(n1351), .IN2(n1352), .IN3(n1353), .QN(\CARRYB[7][6] )
         );
  XOR3X1 U2384 ( .IN1(\ab[7][12] ), .IN2(\CARRYB[6][12] ), .IN3(\SUMB[6][13] ), 
        .Q(\SUMB[7][12] ) );
  NAND2X1 U2385 ( .IN1(\ab[7][12] ), .IN2(\CARRYB[6][12] ), .QN(n1355) );
  NAND2X0 U2386 ( .IN1(\ab[7][12] ), .IN2(\SUMB[6][13] ), .QN(n1356) );
  NAND2X0 U2387 ( .IN1(\CARRYB[6][12] ), .IN2(\SUMB[6][13] ), .QN(n1357) );
  NAND3X1 U2388 ( .IN1(n1355), .IN2(n1356), .IN3(n1357), .QN(\CARRYB[7][12] )
         );
  NAND2X0 U2389 ( .IN1(\ab[8][12] ), .IN2(\SUMB[7][13] ), .QN(n1358) );
  NAND2X0 U2390 ( .IN1(\ab[8][12] ), .IN2(\CARRYB[7][12] ), .QN(n1359) );
  NAND2X0 U2391 ( .IN1(\SUMB[7][13] ), .IN2(\CARRYB[7][12] ), .QN(n1360) );
  NAND3X1 U2392 ( .IN1(n1358), .IN2(n1359), .IN3(n1360), .QN(\CARRYB[8][12] )
         );
  XOR3X1 U2393 ( .IN1(\CARRYB[5][13] ), .IN2(\ab[6][13] ), .IN3(\SUMB[5][14] ), 
        .Q(\SUMB[6][13] ) );
  NAND2X0 U2394 ( .IN1(\CARRYB[5][13] ), .IN2(\SUMB[5][14] ), .QN(n1361) );
  NAND2X1 U2395 ( .IN1(\CARRYB[5][13] ), .IN2(\ab[6][13] ), .QN(n1362) );
  NAND2X0 U2396 ( .IN1(\SUMB[5][14] ), .IN2(\ab[6][13] ), .QN(n1363) );
  DELLN1X2 U2397 ( .INP(n2230), .Z(n2152) );
  XOR3X1 U2398 ( .IN1(\ab[24][29] ), .IN2(\CARRYB[23][29] ), .IN3(
        \SUMB[23][30] ), .Q(\SUMB[24][29] ) );
  NAND2X0 U2399 ( .IN1(\ab[24][29] ), .IN2(\CARRYB[23][29] ), .QN(n1364) );
  NAND2X1 U2400 ( .IN1(\ab[24][29] ), .IN2(\SUMB[23][30] ), .QN(n1365) );
  NAND2X0 U2401 ( .IN1(\CARRYB[23][29] ), .IN2(\SUMB[23][30] ), .QN(n1366) );
  XOR2X1 U2402 ( .IN1(\ab[25][29] ), .IN2(\SUMB[24][30] ), .Q(n1367) );
  XOR2X1 U2403 ( .IN1(n1367), .IN2(\CARRYB[24][29] ), .Q(\SUMB[25][29] ) );
  NAND2X1 U2404 ( .IN1(\ab[25][29] ), .IN2(\SUMB[24][30] ), .QN(n1368) );
  NAND2X0 U2405 ( .IN1(\ab[25][29] ), .IN2(\CARRYB[24][29] ), .QN(n1369) );
  NAND2X0 U2406 ( .IN1(\SUMB[24][30] ), .IN2(\CARRYB[24][29] ), .QN(n1370) );
  XOR3X1 U2407 ( .IN1(\ab[3][12] ), .IN2(\CARRYB[2][12] ), .IN3(\SUMB[2][13] ), 
        .Q(\SUMB[3][12] ) );
  NAND2X1 U2408 ( .IN1(\ab[3][12] ), .IN2(\CARRYB[2][12] ), .QN(n1371) );
  NAND2X0 U2409 ( .IN1(\ab[3][12] ), .IN2(\SUMB[2][13] ), .QN(n1372) );
  NAND2X0 U2410 ( .IN1(\CARRYB[2][12] ), .IN2(\SUMB[2][13] ), .QN(n1373) );
  NAND3X1 U2411 ( .IN1(n1371), .IN2(n1372), .IN3(n1373), .QN(\CARRYB[3][12] )
         );
  XOR2X1 U2412 ( .IN1(\ab[4][12] ), .IN2(\SUMB[3][13] ), .Q(n1374) );
  XOR2X2 U2413 ( .IN1(n1374), .IN2(\CARRYB[3][12] ), .Q(\SUMB[4][12] ) );
  NAND2X0 U2414 ( .IN1(\ab[4][12] ), .IN2(\SUMB[3][13] ), .QN(n1375) );
  NAND2X0 U2415 ( .IN1(\ab[4][12] ), .IN2(\CARRYB[3][12] ), .QN(n1376) );
  NAND2X0 U2416 ( .IN1(\SUMB[3][13] ), .IN2(\CARRYB[3][12] ), .QN(n1377) );
  XOR3X1 U2417 ( .IN1(n1425), .IN2(\ab[2][13] ), .IN3(\SUMB[1][14] ), .Q(
        \SUMB[2][13] ) );
  NAND2X0 U2418 ( .IN1(n1425), .IN2(\SUMB[1][14] ), .QN(n1378) );
  NAND2X0 U2419 ( .IN1(\SUMB[1][14] ), .IN2(\ab[2][13] ), .QN(n1380) );
  NAND3X1 U2420 ( .IN1(n1900), .IN2(n1901), .IN3(n1902), .QN(\CARRYB[2][12] )
         );
  NAND2X0 U2421 ( .IN1(n9), .IN2(\SUMB[1][13] ), .QN(n1902) );
  XOR3X1 U2422 ( .IN1(\ab[11][28] ), .IN2(\CARRYB[10][28] ), .IN3(
        \SUMB[10][29] ), .Q(\SUMB[11][28] ) );
  NAND2X0 U2423 ( .IN1(\ab[11][28] ), .IN2(\CARRYB[10][28] ), .QN(n1381) );
  NAND2X1 U2424 ( .IN1(\ab[11][28] ), .IN2(\SUMB[10][29] ), .QN(n1382) );
  NAND2X0 U2425 ( .IN1(\CARRYB[10][28] ), .IN2(\SUMB[10][29] ), .QN(n1383) );
  NAND3X1 U2426 ( .IN1(n1381), .IN2(n1382), .IN3(n1383), .QN(\CARRYB[11][28] )
         );
  XOR2X1 U2427 ( .IN1(\ab[12][28] ), .IN2(\SUMB[11][29] ), .Q(n1384) );
  NAND2X0 U2428 ( .IN1(\ab[12][28] ), .IN2(\SUMB[11][29] ), .QN(n1385) );
  NAND2X0 U2429 ( .IN1(\ab[12][28] ), .IN2(\CARRYB[11][28] ), .QN(n1386) );
  NAND2X0 U2430 ( .IN1(\SUMB[11][29] ), .IN2(\CARRYB[11][28] ), .QN(n1387) );
  XOR3X1 U2431 ( .IN1(\ab[20][28] ), .IN2(\CARRYB[19][28] ), .IN3(
        \SUMB[19][29] ), .Q(\SUMB[20][28] ) );
  NAND2X0 U2432 ( .IN1(\ab[20][28] ), .IN2(\CARRYB[19][28] ), .QN(n1388) );
  NAND2X1 U2433 ( .IN1(\ab[20][28] ), .IN2(\SUMB[19][29] ), .QN(n1389) );
  NAND2X0 U2434 ( .IN1(\CARRYB[19][28] ), .IN2(\SUMB[19][29] ), .QN(n1390) );
  NAND3X1 U2435 ( .IN1(n1388), .IN2(n1389), .IN3(n1390), .QN(\CARRYB[20][28] )
         );
  XOR2X1 U2436 ( .IN1(\ab[21][28] ), .IN2(\SUMB[20][29] ), .Q(n1391) );
  XOR2X2 U2437 ( .IN1(n1391), .IN2(\CARRYB[20][28] ), .Q(\SUMB[21][28] ) );
  NAND2X0 U2438 ( .IN1(\ab[21][28] ), .IN2(\SUMB[20][29] ), .QN(n1392) );
  NAND2X0 U2439 ( .IN1(\ab[21][28] ), .IN2(\CARRYB[20][28] ), .QN(n1393) );
  NAND2X0 U2440 ( .IN1(\SUMB[20][29] ), .IN2(\CARRYB[20][28] ), .QN(n1394) );
  NAND3X1 U2441 ( .IN1(n1392), .IN2(n1393), .IN3(n1394), .QN(\CARRYB[21][28] )
         );
  XOR3X1 U2442 ( .IN1(\CARRYB[8][28] ), .IN2(\ab[9][28] ), .IN3(\SUMB[8][29] ), 
        .Q(\SUMB[9][28] ) );
  NAND2X0 U2443 ( .IN1(\CARRYB[8][28] ), .IN2(\SUMB[8][29] ), .QN(n1395) );
  NAND2X1 U2444 ( .IN1(\CARRYB[8][28] ), .IN2(\ab[9][28] ), .QN(n1396) );
  NAND2X0 U2445 ( .IN1(\SUMB[8][29] ), .IN2(\ab[9][28] ), .QN(n1397) );
  XOR3X1 U2446 ( .IN1(\CARRYB[6][28] ), .IN2(\ab[7][28] ), .IN3(\SUMB[6][29] ), 
        .Q(\SUMB[7][28] ) );
  NAND2X0 U2447 ( .IN1(\CARRYB[6][28] ), .IN2(\SUMB[6][29] ), .QN(n1398) );
  NAND2X1 U2448 ( .IN1(\CARRYB[6][28] ), .IN2(\ab[7][28] ), .QN(n1399) );
  NAND2X0 U2449 ( .IN1(\SUMB[6][29] ), .IN2(\ab[7][28] ), .QN(n1400) );
  NAND3X0 U2450 ( .IN1(n1398), .IN2(n1399), .IN3(n1400), .QN(\CARRYB[7][28] )
         );
  XOR2X1 U2451 ( .IN1(n933), .IN2(\ab[0][29] ), .Q(\SUMB[1][28] ) );
  DELLN1X2 U2452 ( .INP(n2211), .Z(n2100) );
  NBUFFX4 U2453 ( .INP(n2211), .Z(n2098) );
  XOR3X1 U2454 ( .IN1(\ab[16][27] ), .IN2(\CARRYB[15][27] ), .IN3(
        \SUMB[15][28] ), .Q(\SUMB[16][27] ) );
  NAND2X0 U2455 ( .IN1(\ab[16][27] ), .IN2(\CARRYB[15][27] ), .QN(n1401) );
  NAND2X1 U2456 ( .IN1(\ab[16][27] ), .IN2(\SUMB[15][28] ), .QN(n1402) );
  NAND2X0 U2457 ( .IN1(\CARRYB[15][27] ), .IN2(\SUMB[15][28] ), .QN(n1403) );
  NAND3X1 U2458 ( .IN1(n1401), .IN2(n1402), .IN3(n1403), .QN(\CARRYB[16][27] )
         );
  XOR2X1 U2459 ( .IN1(\ab[17][27] ), .IN2(\SUMB[16][28] ), .Q(n1404) );
  NAND2X0 U2460 ( .IN1(\ab[17][27] ), .IN2(\SUMB[16][28] ), .QN(n1405) );
  NAND2X0 U2461 ( .IN1(\ab[17][27] ), .IN2(\CARRYB[16][27] ), .QN(n1406) );
  NAND2X0 U2462 ( .IN1(\SUMB[16][28] ), .IN2(\CARRYB[16][27] ), .QN(n1407) );
  XOR3X1 U2463 ( .IN1(\CARRYB[8][27] ), .IN2(\ab[9][27] ), .IN3(\SUMB[8][28] ), 
        .Q(\SUMB[9][27] ) );
  NAND2X0 U2464 ( .IN1(\CARRYB[8][27] ), .IN2(\SUMB[8][28] ), .QN(n1408) );
  NAND2X0 U2465 ( .IN1(\SUMB[8][28] ), .IN2(\ab[9][27] ), .QN(n1410) );
  XOR3X1 U2466 ( .IN1(\ab[10][27] ), .IN2(\CARRYB[9][27] ), .IN3(\SUMB[9][28] ), .Q(\SUMB[10][27] ) );
  NAND2X1 U2467 ( .IN1(\ab[10][27] ), .IN2(\CARRYB[9][27] ), .QN(n1411) );
  NAND2X0 U2468 ( .IN1(\ab[10][27] ), .IN2(\SUMB[9][28] ), .QN(n1412) );
  NAND2X0 U2469 ( .IN1(\CARRYB[9][27] ), .IN2(\SUMB[9][28] ), .QN(n1413) );
  XOR2X1 U2470 ( .IN1(\ab[11][27] ), .IN2(\SUMB[10][28] ), .Q(n1414) );
  NAND2X0 U2471 ( .IN1(\ab[11][27] ), .IN2(\SUMB[10][28] ), .QN(n1415) );
  NAND2X0 U2472 ( .IN1(\ab[11][27] ), .IN2(\CARRYB[10][27] ), .QN(n1416) );
  NAND2X0 U2473 ( .IN1(\SUMB[10][28] ), .IN2(\CARRYB[10][27] ), .QN(n1417) );
  XOR3X1 U2474 ( .IN1(\ab[28][27] ), .IN2(\CARRYB[27][27] ), .IN3(
        \SUMB[27][28] ), .Q(\SUMB[28][27] ) );
  NAND2X0 U2475 ( .IN1(\ab[28][27] ), .IN2(\CARRYB[27][27] ), .QN(n1418) );
  NAND2X1 U2476 ( .IN1(\ab[28][27] ), .IN2(\SUMB[27][28] ), .QN(n1419) );
  NAND2X0 U2477 ( .IN1(\CARRYB[27][27] ), .IN2(\SUMB[27][28] ), .QN(n1420) );
  XOR2X1 U2478 ( .IN1(\ab[29][27] ), .IN2(\SUMB[28][28] ), .Q(n1421) );
  NAND2X0 U2479 ( .IN1(\ab[29][27] ), .IN2(\SUMB[28][28] ), .QN(n1422) );
  NAND2X0 U2480 ( .IN1(\ab[29][27] ), .IN2(\CARRYB[28][27] ), .QN(n1423) );
  NAND2X0 U2481 ( .IN1(\SUMB[28][28] ), .IN2(\CARRYB[28][27] ), .QN(n1424) );
  DELLN1X2 U2482 ( .INP(n2212), .Z(n2102) );
  DELLN1X2 U2483 ( .INP(n2212), .Z(n2103) );
  DELLN1X2 U2484 ( .INP(n2212), .Z(n2101) );
  XOR3X1 U2485 ( .IN1(\ab[24][26] ), .IN2(\CARRYB[23][26] ), .IN3(
        \SUMB[23][27] ), .Q(\SUMB[24][26] ) );
  NAND2X0 U2486 ( .IN1(\ab[24][26] ), .IN2(\CARRYB[23][26] ), .QN(n1426) );
  NAND2X1 U2487 ( .IN1(\ab[24][26] ), .IN2(\SUMB[23][27] ), .QN(n1427) );
  NAND2X0 U2488 ( .IN1(\CARRYB[23][26] ), .IN2(\SUMB[23][27] ), .QN(n1428) );
  NAND3X0 U2489 ( .IN1(n1426), .IN2(n1427), .IN3(n1428), .QN(\CARRYB[24][26] )
         );
  NAND2X0 U2490 ( .IN1(\ab[25][26] ), .IN2(\SUMB[24][27] ), .QN(n1429) );
  NAND2X0 U2491 ( .IN1(\ab[25][26] ), .IN2(\CARRYB[24][26] ), .QN(n1430) );
  NAND2X0 U2492 ( .IN1(\SUMB[24][27] ), .IN2(\CARRYB[24][26] ), .QN(n1431) );
  XOR3X1 U2493 ( .IN1(\ab[17][1] ), .IN2(\CARRYB[16][1] ), .IN3(\SUMB[16][2] ), 
        .Q(\SUMB[17][1] ) );
  NAND2X0 U2494 ( .IN1(\ab[17][1] ), .IN2(\CARRYB[16][1] ), .QN(n1432) );
  NAND2X0 U2495 ( .IN1(\CARRYB[16][1] ), .IN2(\SUMB[16][2] ), .QN(n1434) );
  NAND3X1 U2496 ( .IN1(n1433), .IN2(n1432), .IN3(n1434), .QN(\CARRYB[17][1] )
         );
  XOR2X1 U2497 ( .IN1(\ab[18][1] ), .IN2(\SUMB[17][2] ), .Q(n1435) );
  NAND2X0 U2498 ( .IN1(\ab[18][1] ), .IN2(\SUMB[17][2] ), .QN(n1436) );
  NAND2X0 U2499 ( .IN1(\ab[18][1] ), .IN2(\CARRYB[17][1] ), .QN(n1437) );
  NAND2X0 U2500 ( .IN1(\SUMB[17][2] ), .IN2(n19), .QN(n1438) );
  NAND3X1 U2501 ( .IN1(n1436), .IN2(n1437), .IN3(n1438), .QN(\CARRYB[18][1] )
         );
  DELLN1X2 U2502 ( .INP(n2213), .Z(n2106) );
  DELLN1X2 U2503 ( .INP(n2236), .Z(n2168) );
  XOR3X1 U2504 ( .IN1(\ab[30][25] ), .IN2(\CARRYB[29][25] ), .IN3(
        \SUMB[29][26] ), .Q(\SUMB[30][25] ) );
  NAND2X0 U2505 ( .IN1(\ab[30][25] ), .IN2(\CARRYB[29][25] ), .QN(n1439) );
  NAND2X1 U2506 ( .IN1(\ab[30][25] ), .IN2(\SUMB[29][26] ), .QN(n1440) );
  NAND2X0 U2507 ( .IN1(\CARRYB[29][25] ), .IN2(\SUMB[29][26] ), .QN(n1441) );
  XOR2X1 U2508 ( .IN1(\ab[31][25] ), .IN2(\SUMB[30][26] ), .Q(n1442) );
  NAND2X0 U2509 ( .IN1(\ab[31][25] ), .IN2(\SUMB[30][26] ), .QN(n1443) );
  NAND2X0 U2510 ( .IN1(\ab[31][25] ), .IN2(\CARRYB[30][25] ), .QN(n1444) );
  NAND2X0 U2511 ( .IN1(\SUMB[30][26] ), .IN2(\CARRYB[30][25] ), .QN(n1445) );
  XOR3X1 U2512 ( .IN1(\ab[8][25] ), .IN2(\CARRYB[7][25] ), .IN3(\SUMB[7][26] ), 
        .Q(\SUMB[8][25] ) );
  NAND2X0 U2513 ( .IN1(\ab[8][25] ), .IN2(\CARRYB[7][25] ), .QN(n1446) );
  NAND2X0 U2514 ( .IN1(\CARRYB[7][25] ), .IN2(\SUMB[7][26] ), .QN(n1448) );
  XOR2X1 U2515 ( .IN1(\ab[9][25] ), .IN2(\SUMB[8][26] ), .Q(n1449) );
  NAND2X0 U2516 ( .IN1(\ab[9][25] ), .IN2(\SUMB[8][26] ), .QN(n1450) );
  NAND2X0 U2517 ( .IN1(\ab[9][25] ), .IN2(\CARRYB[8][25] ), .QN(n1451) );
  NAND2X0 U2518 ( .IN1(\SUMB[8][26] ), .IN2(\CARRYB[8][25] ), .QN(n1452) );
  NAND3X1 U2519 ( .IN1(n1450), .IN2(n1451), .IN3(n1452), .QN(\CARRYB[9][25] )
         );
  XOR3X1 U2520 ( .IN1(\ab[2][25] ), .IN2(n10), .IN3(\SUMB[1][26] ), .Q(
        \SUMB[2][25] ) );
  NAND2X0 U2521 ( .IN1(\ab[2][25] ), .IN2(n10), .QN(n1453) );
  NAND2X1 U2522 ( .IN1(\ab[2][25] ), .IN2(\SUMB[1][26] ), .QN(n1454) );
  NAND2X0 U2523 ( .IN1(n10), .IN2(\SUMB[1][26] ), .QN(n1455) );
  NAND3X1 U2524 ( .IN1(n1453), .IN2(n1454), .IN3(n1455), .QN(\CARRYB[2][25] )
         );
  XOR2X1 U2525 ( .IN1(\ab[3][25] ), .IN2(\SUMB[2][26] ), .Q(n1456) );
  NAND2X0 U2526 ( .IN1(\ab[3][25] ), .IN2(\SUMB[2][26] ), .QN(n1457) );
  NAND2X0 U2527 ( .IN1(\ab[3][25] ), .IN2(\CARRYB[2][25] ), .QN(n1458) );
  NAND2X0 U2528 ( .IN1(\SUMB[2][26] ), .IN2(\CARRYB[2][25] ), .QN(n1459) );
  XOR3X1 U2529 ( .IN1(\ab[25][25] ), .IN2(\CARRYB[24][25] ), .IN3(
        \SUMB[24][26] ), .Q(\SUMB[25][25] ) );
  NAND2X0 U2530 ( .IN1(\ab[25][25] ), .IN2(\CARRYB[24][25] ), .QN(n1460) );
  NAND2X1 U2531 ( .IN1(\ab[25][25] ), .IN2(\SUMB[24][26] ), .QN(n1461) );
  NAND2X0 U2532 ( .IN1(\CARRYB[24][25] ), .IN2(\SUMB[24][26] ), .QN(n1462) );
  XOR2X1 U2533 ( .IN1(\ab[26][25] ), .IN2(\SUMB[25][26] ), .Q(n1463) );
  XOR2X2 U2534 ( .IN1(n1463), .IN2(\CARRYB[25][25] ), .Q(\SUMB[26][25] ) );
  NAND2X0 U2535 ( .IN1(\ab[26][25] ), .IN2(n836), .QN(n1464) );
  NAND2X1 U2536 ( .IN1(\ab[26][25] ), .IN2(\CARRYB[25][25] ), .QN(n1465) );
  NAND2X0 U2537 ( .IN1(\CARRYB[25][25] ), .IN2(n836), .QN(n1466) );
  XOR3X1 U2538 ( .IN1(\CARRYB[23][25] ), .IN2(\ab[24][25] ), .IN3(
        \SUMB[23][26] ), .Q(\SUMB[24][25] ) );
  NAND2X0 U2539 ( .IN1(\CARRYB[23][25] ), .IN2(\SUMB[23][26] ), .QN(n1467) );
  NAND2X0 U2540 ( .IN1(\CARRYB[23][25] ), .IN2(\ab[24][25] ), .QN(n1468) );
  NAND2X0 U2541 ( .IN1(\SUMB[23][26] ), .IN2(\ab[24][25] ), .QN(n1469) );
  XOR2X2 U2542 ( .IN1(\ab[1][25] ), .IN2(\ab[0][26] ), .Q(\SUMB[1][25] ) );
  XOR2X1 U2543 ( .IN1(\ab[26][14] ), .IN2(\CARRYB[25][14] ), .Q(n1470) );
  NAND2X0 U2544 ( .IN1(\ab[25][15] ), .IN2(\SUMB[24][16] ), .QN(n1472) );
  NAND2X0 U2545 ( .IN1(\CARRYB[24][15] ), .IN2(\SUMB[24][16] ), .QN(n1473) );
  NAND2X0 U2546 ( .IN1(\ab[26][14] ), .IN2(\CARRYB[25][14] ), .QN(n1474) );
  NAND2X0 U2547 ( .IN1(\ab[26][14] ), .IN2(\SUMB[25][15] ), .QN(n1475) );
  NAND2X0 U2548 ( .IN1(\CARRYB[25][14] ), .IN2(\SUMB[25][15] ), .QN(n1476) );
  NAND2X0 U2549 ( .IN1(\ab[21][16] ), .IN2(\CARRYB[20][16] ), .QN(n1477) );
  NAND2X1 U2550 ( .IN1(\ab[21][16] ), .IN2(\SUMB[20][17] ), .QN(n1478) );
  NAND2X0 U2551 ( .IN1(\CARRYB[20][16] ), .IN2(\SUMB[20][17] ), .QN(n1479) );
  XOR2X1 U2552 ( .IN1(\ab[22][16] ), .IN2(\SUMB[21][17] ), .Q(n1480) );
  NAND2X0 U2553 ( .IN1(\ab[22][16] ), .IN2(\SUMB[21][17] ), .QN(n1481) );
  NAND2X0 U2554 ( .IN1(\ab[22][16] ), .IN2(\CARRYB[21][16] ), .QN(n1482) );
  NAND2X0 U2555 ( .IN1(\SUMB[21][17] ), .IN2(\CARRYB[21][16] ), .QN(n1483) );
  XOR3X1 U2556 ( .IN1(\ab[30][24] ), .IN2(\CARRYB[29][24] ), .IN3(
        \SUMB[29][25] ), .Q(\SUMB[30][24] ) );
  NAND2X0 U2557 ( .IN1(\ab[30][24] ), .IN2(\CARRYB[29][24] ), .QN(n1484) );
  NAND2X1 U2558 ( .IN1(\ab[30][24] ), .IN2(\SUMB[29][25] ), .QN(n1485) );
  NAND2X0 U2559 ( .IN1(\CARRYB[29][24] ), .IN2(\SUMB[29][25] ), .QN(n1486) );
  XOR2X1 U2560 ( .IN1(\ab[31][24] ), .IN2(\SUMB[30][25] ), .Q(n1487) );
  NAND2X0 U2561 ( .IN1(\ab[31][24] ), .IN2(\SUMB[30][25] ), .QN(n1488) );
  NAND2X0 U2562 ( .IN1(\ab[31][24] ), .IN2(\CARRYB[30][24] ), .QN(n1489) );
  NAND2X0 U2563 ( .IN1(\SUMB[30][25] ), .IN2(\CARRYB[30][24] ), .QN(n1490) );
  XOR3X1 U2564 ( .IN1(\ab[8][24] ), .IN2(\CARRYB[7][24] ), .IN3(\SUMB[7][25] ), 
        .Q(\SUMB[8][24] ) );
  NAND2X0 U2565 ( .IN1(\ab[8][24] ), .IN2(\CARRYB[7][24] ), .QN(n1491) );
  NAND2X1 U2566 ( .IN1(\ab[8][24] ), .IN2(\SUMB[7][25] ), .QN(n1492) );
  NAND2X0 U2567 ( .IN1(\CARRYB[7][24] ), .IN2(\SUMB[7][25] ), .QN(n1493) );
  NAND3X1 U2568 ( .IN1(n1491), .IN2(n1492), .IN3(n1493), .QN(\CARRYB[8][24] )
         );
  XOR2X1 U2569 ( .IN1(\ab[9][24] ), .IN2(\SUMB[8][25] ), .Q(n1494) );
  NAND2X0 U2570 ( .IN1(\ab[9][24] ), .IN2(\SUMB[8][25] ), .QN(n1495) );
  NAND2X0 U2571 ( .IN1(\ab[9][24] ), .IN2(\CARRYB[8][24] ), .QN(n1496) );
  NAND2X0 U2572 ( .IN1(\SUMB[8][25] ), .IN2(\CARRYB[8][24] ), .QN(n1497) );
  XOR3X1 U2573 ( .IN1(\ab[2][24] ), .IN2(n11), .IN3(\SUMB[1][25] ), .Q(
        \SUMB[2][24] ) );
  NAND2X0 U2574 ( .IN1(\ab[2][24] ), .IN2(n11), .QN(n1498) );
  NAND2X1 U2575 ( .IN1(\ab[2][24] ), .IN2(\SUMB[1][25] ), .QN(n1499) );
  NAND2X0 U2576 ( .IN1(n11), .IN2(\SUMB[1][25] ), .QN(n1500) );
  NAND3X1 U2577 ( .IN1(n1498), .IN2(n1499), .IN3(n1500), .QN(\CARRYB[2][24] )
         );
  XOR2X1 U2578 ( .IN1(\ab[3][24] ), .IN2(\SUMB[2][25] ), .Q(n1501) );
  XOR2X2 U2579 ( .IN1(n1501), .IN2(\CARRYB[2][24] ), .Q(\SUMB[3][24] ) );
  NAND2X0 U2580 ( .IN1(\ab[3][24] ), .IN2(\SUMB[2][25] ), .QN(n1502) );
  NAND2X0 U2581 ( .IN1(\ab[3][24] ), .IN2(\CARRYB[2][24] ), .QN(n1503) );
  NAND2X0 U2582 ( .IN1(\SUMB[2][25] ), .IN2(\CARRYB[2][24] ), .QN(n1504) );
  XOR3X1 U2583 ( .IN1(\ab[25][24] ), .IN2(\CARRYB[24][24] ), .IN3(
        \SUMB[24][25] ), .Q(\SUMB[25][24] ) );
  NAND2X0 U2584 ( .IN1(\ab[25][24] ), .IN2(\CARRYB[24][24] ), .QN(n1505) );
  NAND2X0 U2585 ( .IN1(\CARRYB[24][24] ), .IN2(\SUMB[24][25] ), .QN(n1507) );
  XOR2X1 U2586 ( .IN1(\ab[26][24] ), .IN2(\SUMB[25][25] ), .Q(n1508) );
  NAND2X0 U2587 ( .IN1(\ab[26][24] ), .IN2(\SUMB[25][25] ), .QN(n1509) );
  NAND2X0 U2588 ( .IN1(\ab[26][24] ), .IN2(\CARRYB[25][24] ), .QN(n1510) );
  NAND2X0 U2589 ( .IN1(\SUMB[25][25] ), .IN2(\CARRYB[25][24] ), .QN(n1511) );
  NAND2X0 U2590 ( .IN1(\CARRYB[23][24] ), .IN2(\SUMB[23][25] ), .QN(n1512) );
  NAND2X0 U2591 ( .IN1(\CARRYB[23][24] ), .IN2(\ab[24][24] ), .QN(n1513) );
  NAND2X0 U2592 ( .IN1(\SUMB[23][25] ), .IN2(\ab[24][24] ), .QN(n1514) );
  XOR2X2 U2593 ( .IN1(\ab[1][24] ), .IN2(\ab[0][25] ), .Q(\SUMB[1][24] ) );
  XOR3X1 U2594 ( .IN1(\ab[24][23] ), .IN2(\CARRYB[23][23] ), .IN3(
        \SUMB[23][24] ), .Q(\SUMB[24][23] ) );
  NAND2X0 U2595 ( .IN1(\ab[24][23] ), .IN2(\CARRYB[23][23] ), .QN(n1515) );
  NAND2X1 U2596 ( .IN1(\ab[24][23] ), .IN2(\SUMB[23][24] ), .QN(n1516) );
  NAND2X0 U2597 ( .IN1(\CARRYB[23][23] ), .IN2(\SUMB[23][24] ), .QN(n1517) );
  XOR2X1 U2598 ( .IN1(\ab[25][23] ), .IN2(\SUMB[24][24] ), .Q(n1518) );
  NAND2X0 U2599 ( .IN1(\ab[25][23] ), .IN2(\SUMB[24][24] ), .QN(n1519) );
  NAND2X0 U2600 ( .IN1(\ab[25][23] ), .IN2(\CARRYB[24][23] ), .QN(n1520) );
  NAND2X0 U2601 ( .IN1(\SUMB[24][24] ), .IN2(\CARRYB[24][23] ), .QN(n1521) );
  NAND3X1 U2602 ( .IN1(n1519), .IN2(n1520), .IN3(n1521), .QN(\CARRYB[25][23] )
         );
  XOR3X1 U2603 ( .IN1(\CARRYB[4][23] ), .IN2(\ab[5][23] ), .IN3(\SUMB[4][24] ), 
        .Q(\SUMB[5][23] ) );
  NAND2X0 U2604 ( .IN1(\CARRYB[4][23] ), .IN2(\SUMB[4][24] ), .QN(n1522) );
  NAND2X0 U2605 ( .IN1(\SUMB[4][24] ), .IN2(\ab[5][23] ), .QN(n1524) );
  NAND2X0 U2606 ( .IN1(\CARRYB[12][16] ), .IN2(\SUMB[12][17] ), .QN(n1525) );
  NAND2X0 U2607 ( .IN1(\SUMB[12][17] ), .IN2(\ab[13][16] ), .QN(n1527) );
  NAND2X1 U2608 ( .IN1(\ab[26][15] ), .IN2(\CARRYB[25][15] ), .QN(n1528) );
  NAND2X0 U2609 ( .IN1(\ab[26][15] ), .IN2(\SUMB[25][16] ), .QN(n1529) );
  NAND2X0 U2610 ( .IN1(\CARRYB[25][15] ), .IN2(\SUMB[25][16] ), .QN(n1530) );
  XOR2X1 U2611 ( .IN1(\ab[27][15] ), .IN2(\SUMB[26][16] ), .Q(n1531) );
  XOR2X2 U2612 ( .IN1(n1531), .IN2(\CARRYB[26][15] ), .Q(\SUMB[27][15] ) );
  NAND2X0 U2613 ( .IN1(\ab[27][15] ), .IN2(\SUMB[26][16] ), .QN(n1532) );
  NAND2X0 U2614 ( .IN1(\ab[27][15] ), .IN2(\CARRYB[26][15] ), .QN(n1533) );
  NAND2X0 U2615 ( .IN1(\SUMB[26][16] ), .IN2(\CARRYB[26][15] ), .QN(n1534) );
  NAND2X0 U2616 ( .IN1(\ab[24][22] ), .IN2(\CARRYB[23][22] ), .QN(n1535) );
  NAND2X0 U2617 ( .IN1(\CARRYB[23][22] ), .IN2(\SUMB[23][23] ), .QN(n1537) );
  NAND3X1 U2618 ( .IN1(n1535), .IN2(n1536), .IN3(n1537), .QN(\CARRYB[24][22] )
         );
  XOR2X1 U2619 ( .IN1(\ab[25][22] ), .IN2(\SUMB[24][23] ), .Q(n1538) );
  NAND2X0 U2620 ( .IN1(\ab[25][22] ), .IN2(\SUMB[24][23] ), .QN(n1539) );
  NAND2X0 U2621 ( .IN1(\ab[25][22] ), .IN2(\CARRYB[24][22] ), .QN(n1540) );
  NAND2X0 U2622 ( .IN1(\SUMB[24][23] ), .IN2(\CARRYB[24][22] ), .QN(n1541) );
  XOR3X1 U2623 ( .IN1(\ab[5][22] ), .IN2(\CARRYB[4][22] ), .IN3(\SUMB[4][23] ), 
        .Q(\SUMB[5][22] ) );
  NAND2X0 U2624 ( .IN1(\ab[5][22] ), .IN2(\CARRYB[4][22] ), .QN(n1542) );
  NAND2X1 U2625 ( .IN1(\ab[5][22] ), .IN2(\SUMB[4][23] ), .QN(n1543) );
  NAND2X0 U2626 ( .IN1(\CARRYB[4][22] ), .IN2(\SUMB[4][23] ), .QN(n1544) );
  XOR2X1 U2627 ( .IN1(\ab[6][22] ), .IN2(\SUMB[5][23] ), .Q(n1545) );
  XOR2X2 U2628 ( .IN1(n1545), .IN2(\CARRYB[5][22] ), .Q(\SUMB[6][22] ) );
  NAND2X0 U2629 ( .IN1(\ab[6][22] ), .IN2(\SUMB[5][23] ), .QN(n1546) );
  NAND2X0 U2630 ( .IN1(\ab[6][22] ), .IN2(\CARRYB[5][22] ), .QN(n1547) );
  NAND2X0 U2631 ( .IN1(\SUMB[5][23] ), .IN2(\CARRYB[5][22] ), .QN(n1548) );
  NAND3X1 U2632 ( .IN1(n1546), .IN2(n1547), .IN3(n1548), .QN(\CARRYB[6][22] )
         );
  DELLN1X2 U2633 ( .INP(n2217), .Z(n2116) );
  DELLN1X2 U2634 ( .INP(n2217), .Z(n2118) );
  XOR3X1 U2635 ( .IN1(\ab[10][14] ), .IN2(\CARRYB[9][14] ), .IN3(\SUMB[9][15] ), .Q(\SUMB[10][14] ) );
  NAND2X0 U2636 ( .IN1(\ab[10][14] ), .IN2(\CARRYB[9][14] ), .QN(n1549) );
  NAND2X1 U2637 ( .IN1(\ab[10][14] ), .IN2(\SUMB[9][15] ), .QN(n1550) );
  NAND2X0 U2638 ( .IN1(\CARRYB[9][14] ), .IN2(\SUMB[9][15] ), .QN(n1551) );
  NAND3X1 U2639 ( .IN1(n1549), .IN2(n1550), .IN3(n1551), .QN(\CARRYB[10][14] )
         );
  XOR2X1 U2640 ( .IN1(\ab[11][14] ), .IN2(n49), .Q(n1552) );
  XOR2X2 U2641 ( .IN1(n1552), .IN2(\CARRYB[10][14] ), .Q(\SUMB[11][14] ) );
  NAND2X0 U2642 ( .IN1(\ab[11][14] ), .IN2(\SUMB[10][15] ), .QN(n1553) );
  NAND2X0 U2643 ( .IN1(\ab[11][14] ), .IN2(\CARRYB[10][14] ), .QN(n1554) );
  NAND2X0 U2644 ( .IN1(\SUMB[10][15] ), .IN2(\CARRYB[10][14] ), .QN(n1555) );
  XOR3X1 U2645 ( .IN1(\ab[15][11] ), .IN2(\CARRYB[14][11] ), .IN3(
        \SUMB[14][12] ), .Q(\SUMB[15][11] ) );
  NAND2X1 U2646 ( .IN1(\ab[15][11] ), .IN2(\CARRYB[14][11] ), .QN(n1556) );
  NAND2X0 U2647 ( .IN1(\ab[15][11] ), .IN2(\SUMB[14][12] ), .QN(n1557) );
  NAND2X0 U2648 ( .IN1(\CARRYB[14][11] ), .IN2(\SUMB[14][12] ), .QN(n1558) );
  XOR2X1 U2649 ( .IN1(\ab[16][11] ), .IN2(\SUMB[15][12] ), .Q(n1559) );
  XOR2X2 U2650 ( .IN1(n1559), .IN2(\CARRYB[15][11] ), .Q(\SUMB[16][11] ) );
  NAND2X0 U2651 ( .IN1(\ab[16][11] ), .IN2(\SUMB[15][12] ), .QN(n1560) );
  NAND2X0 U2652 ( .IN1(\ab[16][11] ), .IN2(\CARRYB[15][11] ), .QN(n1561) );
  NAND2X0 U2653 ( .IN1(\SUMB[15][12] ), .IN2(\CARRYB[15][11] ), .QN(n1562) );
  XOR3X1 U2654 ( .IN1(\ab[26][30] ), .IN2(\CARRYB[25][30] ), .IN3(\ab[25][31] ), .Q(\SUMB[26][30] ) );
  NAND2X0 U2655 ( .IN1(\ab[26][30] ), .IN2(\CARRYB[25][30] ), .QN(n1563) );
  NAND2X1 U2656 ( .IN1(\ab[26][30] ), .IN2(\ab[25][31] ), .QN(n1564) );
  NAND2X0 U2657 ( .IN1(\CARRYB[25][30] ), .IN2(\ab[25][31] ), .QN(n1565) );
  XOR2X1 U2658 ( .IN1(\ab[27][30] ), .IN2(\ab[26][31] ), .Q(n1566) );
  XOR2X1 U2659 ( .IN1(n1566), .IN2(\CARRYB[26][30] ), .Q(\SUMB[27][30] ) );
  NAND2X1 U2660 ( .IN1(\ab[27][30] ), .IN2(\ab[26][31] ), .QN(n1567) );
  NAND2X0 U2661 ( .IN1(\ab[27][30] ), .IN2(\CARRYB[26][30] ), .QN(n1568) );
  NAND2X0 U2662 ( .IN1(\ab[26][31] ), .IN2(\CARRYB[26][30] ), .QN(n1569) );
  XOR2X1 U2663 ( .IN1(\ab[25][30] ), .IN2(\ab[24][31] ), .Q(n1570) );
  XOR2X1 U2664 ( .IN1(n1570), .IN2(\CARRYB[24][30] ), .Q(\SUMB[25][30] ) );
  NAND2X0 U2665 ( .IN1(\CARRYB[24][30] ), .IN2(\ab[24][31] ), .QN(n1571) );
  NAND2X0 U2666 ( .IN1(\CARRYB[24][30] ), .IN2(\ab[25][30] ), .QN(n1572) );
  NAND2X1 U2667 ( .IN1(\ab[24][31] ), .IN2(\ab[25][30] ), .QN(n1573) );
  XOR3X1 U2668 ( .IN1(\ab[16][30] ), .IN2(\CARRYB[15][30] ), .IN3(\ab[15][31] ), .Q(\SUMB[16][30] ) );
  NAND2X0 U2669 ( .IN1(\ab[16][30] ), .IN2(\CARRYB[15][30] ), .QN(n1574) );
  NAND2X1 U2670 ( .IN1(\ab[16][30] ), .IN2(\ab[15][31] ), .QN(n1575) );
  NAND2X0 U2671 ( .IN1(\CARRYB[15][30] ), .IN2(\ab[15][31] ), .QN(n1576) );
  XOR2X1 U2672 ( .IN1(\ab[17][30] ), .IN2(\ab[16][31] ), .Q(n1577) );
  XOR2X1 U2673 ( .IN1(n1577), .IN2(\CARRYB[16][30] ), .Q(\SUMB[17][30] ) );
  NAND2X1 U2674 ( .IN1(\ab[17][30] ), .IN2(\ab[16][31] ), .QN(n1578) );
  NAND2X0 U2675 ( .IN1(\ab[17][30] ), .IN2(\CARRYB[16][30] ), .QN(n1579) );
  NAND2X0 U2676 ( .IN1(\ab[16][31] ), .IN2(\CARRYB[16][30] ), .QN(n1580) );
  DELLN1X2 U2677 ( .INP(n2208), .Z(n2094) );
  XOR3X1 U2678 ( .IN1(\ab[24][20] ), .IN2(\CARRYB[23][20] ), .IN3(
        \SUMB[23][21] ), .Q(\SUMB[24][20] ) );
  NAND2X0 U2679 ( .IN1(\ab[24][20] ), .IN2(\CARRYB[23][20] ), .QN(n1582) );
  NAND2X1 U2680 ( .IN1(\ab[24][20] ), .IN2(\SUMB[23][21] ), .QN(n1583) );
  NAND2X0 U2681 ( .IN1(\CARRYB[23][20] ), .IN2(\SUMB[23][21] ), .QN(n1584) );
  NAND3X1 U2682 ( .IN1(n1582), .IN2(n1583), .IN3(n1584), .QN(\CARRYB[24][20] )
         );
  XOR2X1 U2683 ( .IN1(\ab[25][20] ), .IN2(\SUMB[24][21] ), .Q(n1585) );
  XOR2X2 U2684 ( .IN1(n1585), .IN2(\CARRYB[24][20] ), .Q(\SUMB[25][20] ) );
  NAND2X0 U2685 ( .IN1(\ab[25][20] ), .IN2(\SUMB[24][21] ), .QN(n1586) );
  NAND2X0 U2686 ( .IN1(\ab[25][20] ), .IN2(\CARRYB[24][20] ), .QN(n1587) );
  NAND2X0 U2687 ( .IN1(\CARRYB[24][20] ), .IN2(\SUMB[24][21] ), .QN(n1588) );
  NAND3X1 U2688 ( .IN1(n1586), .IN2(n1587), .IN3(n1588), .QN(\CARRYB[25][20] )
         );
  XOR3X1 U2689 ( .IN1(\ab[5][20] ), .IN2(\CARRYB[4][20] ), .IN3(\SUMB[4][21] ), 
        .Q(\SUMB[5][20] ) );
  NAND2X0 U2690 ( .IN1(\ab[5][20] ), .IN2(\CARRYB[4][20] ), .QN(n1589) );
  NAND2X1 U2691 ( .IN1(\ab[5][20] ), .IN2(\SUMB[4][21] ), .QN(n1590) );
  NAND2X0 U2692 ( .IN1(\CARRYB[4][20] ), .IN2(\SUMB[4][21] ), .QN(n1591) );
  NAND3X1 U2693 ( .IN1(n1589), .IN2(n1590), .IN3(n1591), .QN(\CARRYB[5][20] )
         );
  XOR2X1 U2694 ( .IN1(\ab[6][20] ), .IN2(\SUMB[5][21] ), .Q(n1592) );
  XOR2X2 U2695 ( .IN1(n1592), .IN2(\CARRYB[5][20] ), .Q(\SUMB[6][20] ) );
  NAND2X0 U2696 ( .IN1(\ab[6][20] ), .IN2(\SUMB[5][21] ), .QN(n1593) );
  NAND2X0 U2697 ( .IN1(\ab[6][20] ), .IN2(\CARRYB[5][20] ), .QN(n1594) );
  NAND2X0 U2698 ( .IN1(\SUMB[5][21] ), .IN2(\CARRYB[5][20] ), .QN(n1595) );
  NAND3X1 U2699 ( .IN1(n1593), .IN2(n1594), .IN3(n1595), .QN(\CARRYB[6][20] )
         );
  XOR3X1 U2700 ( .IN1(\CARRYB[2][19] ), .IN2(\ab[3][19] ), .IN3(\SUMB[2][20] ), 
        .Q(\SUMB[3][19] ) );
  NAND2X0 U2701 ( .IN1(\CARRYB[2][19] ), .IN2(\SUMB[2][20] ), .QN(n1596) );
  NAND2X0 U2702 ( .IN1(\CARRYB[2][19] ), .IN2(\ab[3][19] ), .QN(n1597) );
  NAND2X0 U2703 ( .IN1(\SUMB[2][20] ), .IN2(\ab[3][19] ), .QN(n1598) );
  NAND3X0 U2704 ( .IN1(n1596), .IN2(n1597), .IN3(n1598), .QN(\CARRYB[3][19] )
         );
  XOR3X1 U2705 ( .IN1(\ab[4][19] ), .IN2(\CARRYB[3][19] ), .IN3(\SUMB[3][20] ), 
        .Q(\SUMB[4][19] ) );
  NAND2X1 U2706 ( .IN1(\ab[4][19] ), .IN2(\CARRYB[3][19] ), .QN(n1599) );
  NAND2X0 U2707 ( .IN1(\ab[4][19] ), .IN2(\SUMB[3][20] ), .QN(n1600) );
  NAND2X0 U2708 ( .IN1(\CARRYB[3][19] ), .IN2(\SUMB[3][20] ), .QN(n1601) );
  XOR2X1 U2709 ( .IN1(\ab[5][19] ), .IN2(\SUMB[4][20] ), .Q(n1602) );
  NAND2X0 U2710 ( .IN1(\ab[5][19] ), .IN2(\SUMB[4][20] ), .QN(n1603) );
  NAND2X0 U2711 ( .IN1(\ab[5][19] ), .IN2(\CARRYB[4][19] ), .QN(n1604) );
  NAND2X0 U2712 ( .IN1(\SUMB[4][20] ), .IN2(\CARRYB[4][19] ), .QN(n1605) );
  NAND2X0 U2713 ( .IN1(\ab[15][19] ), .IN2(\CARRYB[14][19] ), .QN(n1606) );
  NAND2X1 U2714 ( .IN1(\ab[15][19] ), .IN2(\SUMB[14][20] ), .QN(n1607) );
  NAND2X0 U2715 ( .IN1(\CARRYB[14][19] ), .IN2(\SUMB[14][20] ), .QN(n1608) );
  NAND3X1 U2716 ( .IN1(n1606), .IN2(n1607), .IN3(n1608), .QN(\CARRYB[15][19] )
         );
  XOR2X1 U2717 ( .IN1(\ab[16][19] ), .IN2(\SUMB[15][20] ), .Q(n1609) );
  XOR2X2 U2718 ( .IN1(n1609), .IN2(\CARRYB[15][19] ), .Q(\SUMB[16][19] ) );
  NAND2X0 U2719 ( .IN1(\ab[16][19] ), .IN2(\SUMB[15][20] ), .QN(n1610) );
  NAND2X0 U2720 ( .IN1(\ab[16][19] ), .IN2(\CARRYB[15][19] ), .QN(n1611) );
  NAND2X0 U2721 ( .IN1(\SUMB[15][20] ), .IN2(\CARRYB[15][19] ), .QN(n1612) );
  XOR3X1 U2722 ( .IN1(\ab[13][12] ), .IN2(\CARRYB[12][12] ), .IN3(
        \SUMB[12][13] ), .Q(\SUMB[13][12] ) );
  NAND2X0 U2723 ( .IN1(\ab[13][12] ), .IN2(\CARRYB[12][12] ), .QN(n1613) );
  NAND2X1 U2724 ( .IN1(\ab[13][12] ), .IN2(\SUMB[12][13] ), .QN(n1614) );
  NAND2X0 U2725 ( .IN1(\CARRYB[12][12] ), .IN2(\SUMB[12][13] ), .QN(n1615) );
  NAND3X1 U2726 ( .IN1(n1613), .IN2(n1614), .IN3(n1615), .QN(\CARRYB[13][12] )
         );
  XOR2X1 U2727 ( .IN1(\ab[14][12] ), .IN2(\SUMB[13][13] ), .Q(n1616) );
  NAND2X0 U2728 ( .IN1(\ab[14][12] ), .IN2(\SUMB[13][13] ), .QN(n1617) );
  NAND2X0 U2729 ( .IN1(\ab[14][12] ), .IN2(\CARRYB[13][12] ), .QN(n1618) );
  NAND2X0 U2730 ( .IN1(\SUMB[13][13] ), .IN2(\CARRYB[13][12] ), .QN(n1619) );
  XOR3X1 U2731 ( .IN1(\ab[4][13] ), .IN2(\CARRYB[3][13] ), .IN3(\SUMB[3][14] ), 
        .Q(\SUMB[4][13] ) );
  NAND2X0 U2732 ( .IN1(\ab[4][13] ), .IN2(\CARRYB[3][13] ), .QN(n1620) );
  NAND2X1 U2733 ( .IN1(\ab[4][13] ), .IN2(\SUMB[3][14] ), .QN(n1621) );
  NAND2X0 U2734 ( .IN1(\CARRYB[3][13] ), .IN2(\SUMB[3][14] ), .QN(n1622) );
  XOR2X1 U2735 ( .IN1(\ab[5][13] ), .IN2(\SUMB[4][14] ), .Q(n1623) );
  NAND2X0 U2736 ( .IN1(\ab[5][13] ), .IN2(\SUMB[4][14] ), .QN(n1624) );
  NAND2X0 U2737 ( .IN1(\ab[5][13] ), .IN2(\CARRYB[4][13] ), .QN(n1625) );
  NAND2X0 U2738 ( .IN1(\SUMB[4][14] ), .IN2(\CARRYB[4][13] ), .QN(n1626) );
  XOR3X1 U2739 ( .IN1(n14), .IN2(\ab[2][18] ), .IN3(\SUMB[1][19] ), .Q(
        \SUMB[2][18] ) );
  NAND2X1 U2740 ( .IN1(n14), .IN2(\SUMB[1][19] ), .QN(n1627) );
  NAND2X1 U2741 ( .IN1(n14), .IN2(\ab[2][18] ), .QN(n1628) );
  NAND2X0 U2742 ( .IN1(\SUMB[1][19] ), .IN2(\ab[2][18] ), .QN(n1629) );
  NAND3X0 U2743 ( .IN1(n1627), .IN2(n1628), .IN3(n1629), .QN(\CARRYB[2][18] )
         );
  XOR3X1 U2744 ( .IN1(\ab[3][18] ), .IN2(\CARRYB[2][18] ), .IN3(\SUMB[2][19] ), 
        .Q(\SUMB[3][18] ) );
  NAND2X1 U2745 ( .IN1(\ab[3][18] ), .IN2(\CARRYB[2][18] ), .QN(n1630) );
  NAND2X0 U2746 ( .IN1(\ab[3][18] ), .IN2(\SUMB[2][19] ), .QN(n1631) );
  NAND2X0 U2747 ( .IN1(\CARRYB[2][18] ), .IN2(\SUMB[2][19] ), .QN(n1632) );
  NAND3X1 U2748 ( .IN1(n1630), .IN2(n1631), .IN3(n1632), .QN(\CARRYB[3][18] )
         );
  XOR2X1 U2749 ( .IN1(\ab[4][18] ), .IN2(\SUMB[3][19] ), .Q(n1633) );
  NAND2X0 U2750 ( .IN1(\ab[4][18] ), .IN2(\SUMB[3][19] ), .QN(n1634) );
  NAND2X0 U2751 ( .IN1(\ab[4][18] ), .IN2(\CARRYB[3][18] ), .QN(n1635) );
  NAND2X0 U2752 ( .IN1(\SUMB[3][19] ), .IN2(\CARRYB[3][18] ), .QN(n1636) );
  XOR3X1 U2753 ( .IN1(\ab[20][18] ), .IN2(\CARRYB[19][18] ), .IN3(
        \SUMB[19][19] ), .Q(\SUMB[20][18] ) );
  NAND2X0 U2754 ( .IN1(\ab[20][18] ), .IN2(\CARRYB[19][18] ), .QN(n1637) );
  NAND2X1 U2755 ( .IN1(\ab[20][18] ), .IN2(\SUMB[19][19] ), .QN(n1638) );
  NAND2X0 U2756 ( .IN1(\CARRYB[19][18] ), .IN2(\SUMB[19][19] ), .QN(n1639) );
  XOR2X1 U2757 ( .IN1(\ab[21][18] ), .IN2(\SUMB[20][19] ), .Q(n1640) );
  XOR2X2 U2758 ( .IN1(n1640), .IN2(\CARRYB[20][18] ), .Q(\SUMB[21][18] ) );
  NAND2X0 U2759 ( .IN1(\ab[21][18] ), .IN2(\SUMB[20][19] ), .QN(n1641) );
  NAND2X0 U2760 ( .IN1(\ab[21][18] ), .IN2(\CARRYB[20][18] ), .QN(n1642) );
  NAND2X0 U2761 ( .IN1(\SUMB[20][19] ), .IN2(\CARRYB[20][18] ), .QN(n1643) );
  XOR3X1 U2762 ( .IN1(\ab[12][11] ), .IN2(\CARRYB[11][11] ), .IN3(
        \SUMB[11][12] ), .Q(\SUMB[12][11] ) );
  XOR2X1 U2763 ( .IN1(\ab[13][10] ), .IN2(\CARRYB[12][10] ), .Q(n1644) );
  NAND2X0 U2764 ( .IN1(\ab[12][11] ), .IN2(\CARRYB[11][11] ), .QN(n1645) );
  NAND2X0 U2765 ( .IN1(\ab[12][11] ), .IN2(\SUMB[11][12] ), .QN(n1646) );
  NAND2X0 U2766 ( .IN1(\CARRYB[11][11] ), .IN2(\SUMB[11][12] ), .QN(n1647) );
  NAND2X0 U2767 ( .IN1(\ab[13][10] ), .IN2(\CARRYB[12][10] ), .QN(n1648) );
  NAND2X0 U2768 ( .IN1(\ab[13][10] ), .IN2(\SUMB[12][11] ), .QN(n1649) );
  NAND2X0 U2769 ( .IN1(\SUMB[12][11] ), .IN2(\CARRYB[12][10] ), .QN(n1650) );
  NAND2X0 U2770 ( .IN1(\CARRYB[10][11] ), .IN2(\SUMB[10][12] ), .QN(n1651) );
  NAND2X0 U2771 ( .IN1(\CARRYB[10][11] ), .IN2(\ab[11][11] ), .QN(n1652) );
  XOR3X1 U2772 ( .IN1(\ab[29][17] ), .IN2(\CARRYB[28][17] ), .IN3(
        \SUMB[28][18] ), .Q(\SUMB[29][17] ) );
  NAND2X0 U2773 ( .IN1(\ab[29][17] ), .IN2(\CARRYB[28][17] ), .QN(n1654) );
  NAND2X1 U2774 ( .IN1(\ab[29][17] ), .IN2(\SUMB[28][18] ), .QN(n1655) );
  NAND2X0 U2775 ( .IN1(\CARRYB[28][17] ), .IN2(\SUMB[28][18] ), .QN(n1656) );
  NAND3X1 U2776 ( .IN1(n1654), .IN2(n1655), .IN3(n1656), .QN(\CARRYB[29][17] )
         );
  XOR2X1 U2777 ( .IN1(\ab[30][17] ), .IN2(\SUMB[29][18] ), .Q(n1657) );
  NAND2X0 U2778 ( .IN1(\ab[30][17] ), .IN2(\SUMB[29][18] ), .QN(n1658) );
  NAND2X0 U2779 ( .IN1(\ab[30][17] ), .IN2(\CARRYB[29][17] ), .QN(n1659) );
  NAND2X0 U2780 ( .IN1(\SUMB[29][18] ), .IN2(\CARRYB[29][17] ), .QN(n1660) );
  XOR3X1 U2781 ( .IN1(\ab[20][17] ), .IN2(\CARRYB[19][17] ), .IN3(
        \SUMB[19][18] ), .Q(\SUMB[20][17] ) );
  NAND2X0 U2782 ( .IN1(\ab[20][17] ), .IN2(\CARRYB[19][17] ), .QN(n1661) );
  NAND2X0 U2783 ( .IN1(\CARRYB[19][17] ), .IN2(\SUMB[19][18] ), .QN(n1663) );
  NAND3X1 U2784 ( .IN1(n1661), .IN2(n1662), .IN3(n1663), .QN(\CARRYB[20][17] )
         );
  XOR2X1 U2785 ( .IN1(\ab[21][17] ), .IN2(\SUMB[20][18] ), .Q(n1664) );
  NAND2X0 U2786 ( .IN1(\ab[21][17] ), .IN2(\SUMB[20][18] ), .QN(n1665) );
  NAND2X0 U2787 ( .IN1(\ab[21][17] ), .IN2(\CARRYB[20][17] ), .QN(n1666) );
  NAND2X0 U2788 ( .IN1(\SUMB[20][18] ), .IN2(\CARRYB[20][17] ), .QN(n1667) );
  XOR3X1 U2789 ( .IN1(\ab[26][16] ), .IN2(\CARRYB[25][16] ), .IN3(
        \SUMB[25][17] ), .Q(\SUMB[26][16] ) );
  NAND2X0 U2790 ( .IN1(\ab[26][16] ), .IN2(\CARRYB[25][16] ), .QN(n1668) );
  NAND2X1 U2791 ( .IN1(\ab[26][16] ), .IN2(\SUMB[25][17] ), .QN(n1669) );
  NAND2X0 U2792 ( .IN1(\CARRYB[25][16] ), .IN2(\SUMB[25][17] ), .QN(n1670) );
  NAND3X1 U2793 ( .IN1(n1668), .IN2(n1669), .IN3(n1670), .QN(\CARRYB[26][16] )
         );
  XOR2X1 U2794 ( .IN1(\ab[27][16] ), .IN2(\SUMB[26][17] ), .Q(n1671) );
  NAND2X0 U2795 ( .IN1(\ab[27][16] ), .IN2(\SUMB[26][17] ), .QN(n1672) );
  NAND2X0 U2796 ( .IN1(\ab[27][16] ), .IN2(\CARRYB[26][16] ), .QN(n1673) );
  NAND2X0 U2797 ( .IN1(\SUMB[26][17] ), .IN2(\CARRYB[26][16] ), .QN(n1674) );
  XOR3X1 U2798 ( .IN1(\ab[13][11] ), .IN2(\CARRYB[12][11] ), .IN3(
        \SUMB[12][12] ), .Q(\SUMB[13][11] ) );
  NAND2X0 U2799 ( .IN1(\ab[13][11] ), .IN2(\CARRYB[12][11] ), .QN(n1675) );
  NAND2X1 U2800 ( .IN1(\ab[13][11] ), .IN2(\SUMB[12][12] ), .QN(n1676) );
  NAND2X0 U2801 ( .IN1(\CARRYB[12][11] ), .IN2(\SUMB[12][12] ), .QN(n1677) );
  XOR2X1 U2802 ( .IN1(\ab[14][11] ), .IN2(\SUMB[13][12] ), .Q(n1678) );
  NAND2X0 U2803 ( .IN1(\ab[14][11] ), .IN2(\SUMB[13][12] ), .QN(n1679) );
  NAND2X0 U2804 ( .IN1(\ab[14][11] ), .IN2(\CARRYB[13][11] ), .QN(n1680) );
  NAND2X0 U2805 ( .IN1(\SUMB[13][12] ), .IN2(\CARRYB[13][11] ), .QN(n1681) );
  XOR3X1 U2806 ( .IN1(\ab[18][14] ), .IN2(\CARRYB[17][14] ), .IN3(
        \SUMB[17][15] ), .Q(\SUMB[18][14] ) );
  NAND2X0 U2807 ( .IN1(\ab[18][14] ), .IN2(\CARRYB[17][14] ), .QN(n1682) );
  NAND2X1 U2808 ( .IN1(\ab[18][14] ), .IN2(\SUMB[17][15] ), .QN(n1683) );
  NAND2X0 U2809 ( .IN1(\CARRYB[17][14] ), .IN2(\SUMB[17][15] ), .QN(n1684) );
  XOR2X1 U2810 ( .IN1(\ab[19][14] ), .IN2(\SUMB[18][15] ), .Q(n1685) );
  NAND2X0 U2811 ( .IN1(\ab[19][14] ), .IN2(\SUMB[18][15] ), .QN(n1686) );
  NAND2X0 U2812 ( .IN1(\ab[19][14] ), .IN2(\CARRYB[18][14] ), .QN(n1687) );
  NAND2X0 U2813 ( .IN1(\SUMB[18][15] ), .IN2(\CARRYB[18][14] ), .QN(n1688) );
  XOR3X1 U2814 ( .IN1(\ab[27][6] ), .IN2(\CARRYB[26][6] ), .IN3(\SUMB[26][7] ), 
        .Q(\SUMB[27][6] ) );
  NAND2X0 U2815 ( .IN1(\ab[27][6] ), .IN2(\CARRYB[26][6] ), .QN(n1690) );
  NAND2X1 U2816 ( .IN1(\ab[27][6] ), .IN2(\SUMB[26][7] ), .QN(n1691) );
  NAND2X0 U2817 ( .IN1(\CARRYB[26][6] ), .IN2(\SUMB[26][7] ), .QN(n1692) );
  XOR2X1 U2818 ( .IN1(\ab[28][6] ), .IN2(\SUMB[27][7] ), .Q(n1693) );
  XOR2X2 U2819 ( .IN1(n1693), .IN2(\CARRYB[27][6] ), .Q(\SUMB[28][6] ) );
  NAND2X0 U2820 ( .IN1(\ab[28][6] ), .IN2(\SUMB[27][7] ), .QN(n1694) );
  NAND2X0 U2821 ( .IN1(\ab[28][6] ), .IN2(\CARRYB[27][6] ), .QN(n1695) );
  NAND2X0 U2822 ( .IN1(\SUMB[27][7] ), .IN2(\CARRYB[27][6] ), .QN(n1696) );
  XOR3X1 U2823 ( .IN1(\ab[29][6] ), .IN2(\CARRYB[28][6] ), .IN3(\SUMB[28][7] ), 
        .Q(\SUMB[29][6] ) );
  NAND2X1 U2824 ( .IN1(\ab[29][6] ), .IN2(\CARRYB[28][6] ), .QN(n1697) );
  NAND2X0 U2825 ( .IN1(\ab[29][6] ), .IN2(\SUMB[28][7] ), .QN(n1698) );
  NAND2X0 U2826 ( .IN1(\CARRYB[28][6] ), .IN2(\SUMB[28][7] ), .QN(n1699) );
  NAND2X0 U2827 ( .IN1(\ab[30][6] ), .IN2(\SUMB[29][7] ), .QN(n1700) );
  NAND2X0 U2828 ( .IN1(\ab[30][6] ), .IN2(\CARRYB[29][6] ), .QN(n1701) );
  NAND2X0 U2829 ( .IN1(\SUMB[29][7] ), .IN2(\CARRYB[29][6] ), .QN(n1702) );
  XOR3X1 U2830 ( .IN1(\ab[17][6] ), .IN2(\CARRYB[16][6] ), .IN3(\SUMB[16][7] ), 
        .Q(\SUMB[17][6] ) );
  NAND2X0 U2831 ( .IN1(\ab[17][6] ), .IN2(\CARRYB[16][6] ), .QN(n1703) );
  NAND2X1 U2832 ( .IN1(\ab[17][6] ), .IN2(\SUMB[16][7] ), .QN(n1704) );
  NAND2X0 U2833 ( .IN1(\CARRYB[16][6] ), .IN2(\SUMB[16][7] ), .QN(n1705) );
  NAND3X1 U2834 ( .IN1(n1703), .IN2(n1704), .IN3(n1705), .QN(\CARRYB[17][6] )
         );
  XOR2X1 U2835 ( .IN1(\ab[18][6] ), .IN2(\SUMB[17][7] ), .Q(n1706) );
  NAND2X0 U2836 ( .IN1(\ab[18][6] ), .IN2(\SUMB[17][7] ), .QN(n1707) );
  NAND2X0 U2837 ( .IN1(\ab[18][6] ), .IN2(\CARRYB[17][6] ), .QN(n1708) );
  NAND2X0 U2838 ( .IN1(\SUMB[17][7] ), .IN2(\CARRYB[17][6] ), .QN(n1709) );
  NAND3X1 U2839 ( .IN1(n1707), .IN2(n1708), .IN3(n1709), .QN(\CARRYB[18][6] )
         );
  XOR3X1 U2840 ( .IN1(\ab[2][6] ), .IN2(n12), .IN3(\SUMB[1][7] ), .Q(
        \SUMB[2][6] ) );
  NAND2X0 U2841 ( .IN1(\ab[2][6] ), .IN2(n12), .QN(n1710) );
  NAND2X0 U2842 ( .IN1(\ab[2][6] ), .IN2(\SUMB[1][7] ), .QN(n1711) );
  NAND2X0 U2843 ( .IN1(n12), .IN2(\SUMB[1][7] ), .QN(n1712) );
  NAND3X1 U2844 ( .IN1(n1710), .IN2(n1711), .IN3(n1712), .QN(\CARRYB[2][6] )
         );
  XOR2X1 U2845 ( .IN1(\ab[3][6] ), .IN2(\SUMB[2][7] ), .Q(n1713) );
  NAND2X0 U2846 ( .IN1(\ab[3][6] ), .IN2(\SUMB[2][7] ), .QN(n1714) );
  NAND2X0 U2847 ( .IN1(\ab[3][6] ), .IN2(\CARRYB[2][6] ), .QN(n1715) );
  NAND2X0 U2848 ( .IN1(\SUMB[2][7] ), .IN2(\CARRYB[2][6] ), .QN(n1716) );
  XOR3X1 U2849 ( .IN1(\ab[12][13] ), .IN2(\CARRYB[11][13] ), .IN3(
        \SUMB[11][14] ), .Q(\SUMB[12][13] ) );
  NAND2X0 U2850 ( .IN1(\ab[12][13] ), .IN2(\CARRYB[11][13] ), .QN(n1717) );
  NAND2X1 U2851 ( .IN1(\ab[12][13] ), .IN2(\SUMB[11][14] ), .QN(n1718) );
  NAND2X0 U2852 ( .IN1(\CARRYB[11][13] ), .IN2(\SUMB[11][14] ), .QN(n1719) );
  NAND3X1 U2853 ( .IN1(n1717), .IN2(n1718), .IN3(n1719), .QN(\CARRYB[12][13] )
         );
  XOR2X1 U2854 ( .IN1(\ab[13][13] ), .IN2(\SUMB[12][14] ), .Q(n1720) );
  XOR2X2 U2855 ( .IN1(n1720), .IN2(\CARRYB[12][13] ), .Q(\SUMB[13][13] ) );
  NAND2X0 U2856 ( .IN1(\ab[13][13] ), .IN2(\SUMB[12][14] ), .QN(n1721) );
  NAND2X0 U2857 ( .IN1(\ab[13][13] ), .IN2(\CARRYB[12][13] ), .QN(n1722) );
  NAND2X0 U2858 ( .IN1(\SUMB[12][14] ), .IN2(\CARRYB[12][13] ), .QN(n1723) );
  XOR3X1 U2859 ( .IN1(\ab[27][13] ), .IN2(\CARRYB[26][13] ), .IN3(
        \SUMB[26][14] ), .Q(\SUMB[27][13] ) );
  NAND2X0 U2860 ( .IN1(\ab[27][13] ), .IN2(\CARRYB[26][13] ), .QN(n1724) );
  NAND2X1 U2861 ( .IN1(\ab[27][13] ), .IN2(\SUMB[26][14] ), .QN(n1725) );
  NAND2X0 U2862 ( .IN1(\CARRYB[26][13] ), .IN2(\SUMB[26][14] ), .QN(n1726) );
  NAND3X1 U2863 ( .IN1(n1724), .IN2(n1725), .IN3(n1726), .QN(\CARRYB[27][13] )
         );
  XOR2X1 U2864 ( .IN1(\ab[28][13] ), .IN2(\SUMB[27][14] ), .Q(n1727) );
  NAND2X0 U2865 ( .IN1(\ab[28][13] ), .IN2(\SUMB[27][14] ), .QN(n1728) );
  NAND2X0 U2866 ( .IN1(\ab[28][13] ), .IN2(\CARRYB[27][13] ), .QN(n1729) );
  NAND2X0 U2867 ( .IN1(\SUMB[27][14] ), .IN2(\CARRYB[27][13] ), .QN(n1730) );
  XOR3X1 U2868 ( .IN1(\CARRYB[24][13] ), .IN2(\ab[25][13] ), .IN3(
        \SUMB[24][14] ), .Q(\SUMB[25][13] ) );
  NAND2X0 U2869 ( .IN1(\CARRYB[24][13] ), .IN2(\SUMB[24][14] ), .QN(n1731) );
  NAND2X0 U2870 ( .IN1(\CARRYB[24][13] ), .IN2(\ab[25][13] ), .QN(n1732) );
  NAND2X0 U2871 ( .IN1(\SUMB[24][14] ), .IN2(\ab[25][13] ), .QN(n1733) );
  XOR3X1 U2872 ( .IN1(\ab[7][13] ), .IN2(\CARRYB[6][13] ), .IN3(\SUMB[6][14] ), 
        .Q(\SUMB[7][13] ) );
  NAND2X0 U2873 ( .IN1(\ab[7][13] ), .IN2(\CARRYB[6][13] ), .QN(n1734) );
  NAND2X0 U2874 ( .IN1(\CARRYB[6][13] ), .IN2(\SUMB[6][14] ), .QN(n1736) );
  NAND3X1 U2875 ( .IN1(n1734), .IN2(n1735), .IN3(n1736), .QN(\CARRYB[7][13] )
         );
  XOR2X1 U2876 ( .IN1(\ab[8][13] ), .IN2(\SUMB[7][14] ), .Q(n1737) );
  XOR2X2 U2877 ( .IN1(n1737), .IN2(\CARRYB[7][13] ), .Q(\SUMB[8][13] ) );
  NAND2X0 U2878 ( .IN1(\ab[8][13] ), .IN2(\SUMB[7][14] ), .QN(n1738) );
  NAND2X0 U2879 ( .IN1(\ab[8][13] ), .IN2(\CARRYB[7][13] ), .QN(n1739) );
  NAND2X0 U2880 ( .IN1(\SUMB[7][14] ), .IN2(\CARRYB[7][13] ), .QN(n1740) );
  XOR2X1 U2881 ( .IN1(\ab[31][7] ), .IN2(\SUMB[30][8] ), .Q(n1741) );
  XOR2X1 U2882 ( .IN1(n1741), .IN2(\CARRYB[30][7] ), .Q(\SUMB[31][7] ) );
  NAND2X0 U2883 ( .IN1(\CARRYB[30][7] ), .IN2(\SUMB[30][8] ), .QN(n1742) );
  NAND2X0 U2884 ( .IN1(\CARRYB[30][7] ), .IN2(\ab[31][7] ), .QN(n1743) );
  NAND2X1 U2885 ( .IN1(\SUMB[30][8] ), .IN2(\ab[31][7] ), .QN(n1744) );
  XOR2X1 U2886 ( .IN1(\ab[30][7] ), .IN2(\SUMB[29][8] ), .Q(n1745) );
  NAND2X0 U2887 ( .IN1(\CARRYB[29][7] ), .IN2(\SUMB[29][8] ), .QN(n1746) );
  NAND2X0 U2888 ( .IN1(\CARRYB[29][7] ), .IN2(\ab[30][7] ), .QN(n1747) );
  NAND2X1 U2889 ( .IN1(\SUMB[29][8] ), .IN2(\ab[30][7] ), .QN(n1748) );
  XOR3X1 U2890 ( .IN1(\ab[20][7] ), .IN2(\CARRYB[19][7] ), .IN3(\SUMB[19][8] ), 
        .Q(\SUMB[20][7] ) );
  NAND2X0 U2891 ( .IN1(\ab[20][7] ), .IN2(\CARRYB[19][7] ), .QN(n1749) );
  NAND2X1 U2892 ( .IN1(\ab[20][7] ), .IN2(\SUMB[19][8] ), .QN(n1750) );
  NAND2X0 U2893 ( .IN1(\CARRYB[19][7] ), .IN2(\SUMB[19][8] ), .QN(n1751) );
  XOR2X1 U2894 ( .IN1(\ab[21][7] ), .IN2(\SUMB[20][8] ), .Q(n1752) );
  NAND2X0 U2895 ( .IN1(\ab[21][7] ), .IN2(\SUMB[20][8] ), .QN(n1753) );
  NAND2X0 U2896 ( .IN1(\ab[21][7] ), .IN2(\CARRYB[20][7] ), .QN(n1754) );
  NAND2X0 U2897 ( .IN1(\SUMB[20][8] ), .IN2(\CARRYB[20][7] ), .QN(n1755) );
  XOR3X1 U2898 ( .IN1(\ab[11][7] ), .IN2(\CARRYB[10][7] ), .IN3(\SUMB[10][8] ), 
        .Q(\SUMB[11][7] ) );
  NAND2X0 U2899 ( .IN1(\ab[11][7] ), .IN2(\CARRYB[10][7] ), .QN(n1756) );
  NAND2X1 U2900 ( .IN1(\ab[11][7] ), .IN2(\SUMB[10][8] ), .QN(n1757) );
  NAND2X0 U2901 ( .IN1(\CARRYB[10][7] ), .IN2(\SUMB[10][8] ), .QN(n1758) );
  NAND3X1 U2902 ( .IN1(n1756), .IN2(n1757), .IN3(n1758), .QN(\CARRYB[11][7] )
         );
  XOR2X1 U2903 ( .IN1(\ab[12][7] ), .IN2(\SUMB[11][8] ), .Q(n1759) );
  NAND2X0 U2904 ( .IN1(\ab[12][7] ), .IN2(\SUMB[11][8] ), .QN(n1760) );
  NAND2X0 U2905 ( .IN1(\ab[12][7] ), .IN2(\CARRYB[11][7] ), .QN(n1761) );
  NAND2X0 U2906 ( .IN1(\SUMB[11][8] ), .IN2(\CARRYB[11][7] ), .QN(n1762) );
  NAND3X1 U2907 ( .IN1(n1760), .IN2(n1761), .IN3(n1762), .QN(\CARRYB[12][7] )
         );
  XOR3X1 U2908 ( .IN1(\ab[19][9] ), .IN2(\CARRYB[18][9] ), .IN3(\SUMB[18][10] ), .Q(\SUMB[19][9] ) );
  NAND2X0 U2909 ( .IN1(\ab[19][9] ), .IN2(\CARRYB[18][9] ), .QN(n1764) );
  NAND2X1 U2910 ( .IN1(\ab[19][9] ), .IN2(\SUMB[18][10] ), .QN(n1765) );
  NAND2X0 U2911 ( .IN1(\CARRYB[18][9] ), .IN2(\SUMB[18][10] ), .QN(n1766) );
  XOR2X1 U2912 ( .IN1(\ab[20][9] ), .IN2(\SUMB[19][10] ), .Q(n1767) );
  XOR2X2 U2913 ( .IN1(n1767), .IN2(\CARRYB[19][9] ), .Q(\SUMB[20][9] ) );
  NAND2X0 U2914 ( .IN1(\ab[20][9] ), .IN2(\SUMB[19][10] ), .QN(n1768) );
  NAND2X0 U2915 ( .IN1(\ab[20][9] ), .IN2(\CARRYB[19][9] ), .QN(n1769) );
  NAND2X0 U2916 ( .IN1(\SUMB[19][10] ), .IN2(\CARRYB[19][9] ), .QN(n1770) );
  NAND3X1 U2917 ( .IN1(n1768), .IN2(n1769), .IN3(n1770), .QN(\CARRYB[20][9] )
         );
  XOR2X1 U2918 ( .IN1(\ab[18][9] ), .IN2(\SUMB[17][10] ), .Q(n1771) );
  NAND2X0 U2919 ( .IN1(\CARRYB[17][9] ), .IN2(\SUMB[17][10] ), .QN(n1772) );
  NAND2X0 U2920 ( .IN1(\CARRYB[17][9] ), .IN2(\ab[18][9] ), .QN(n1773) );
  NAND2X0 U2921 ( .IN1(\SUMB[17][10] ), .IN2(\ab[18][9] ), .QN(n1774) );
  XOR3X1 U2922 ( .IN1(\ab[6][9] ), .IN2(\CARRYB[5][9] ), .IN3(\SUMB[5][10] ), 
        .Q(\SUMB[6][9] ) );
  NAND2X0 U2923 ( .IN1(\ab[6][9] ), .IN2(\SUMB[5][10] ), .QN(n1776) );
  NAND2X0 U2924 ( .IN1(\CARRYB[5][9] ), .IN2(\SUMB[5][10] ), .QN(n1777) );
  NAND3X1 U2925 ( .IN1(n1775), .IN2(n1776), .IN3(n1777), .QN(\CARRYB[6][9] )
         );
  XOR2X1 U2926 ( .IN1(\ab[7][9] ), .IN2(\SUMB[6][10] ), .Q(n1778) );
  NAND2X0 U2927 ( .IN1(\ab[7][9] ), .IN2(\SUMB[6][10] ), .QN(n1779) );
  NAND2X0 U2928 ( .IN1(\ab[7][9] ), .IN2(\CARRYB[6][9] ), .QN(n1780) );
  NAND2X0 U2929 ( .IN1(\SUMB[6][10] ), .IN2(\CARRYB[6][9] ), .QN(n1781) );
  NAND3X1 U2930 ( .IN1(n1779), .IN2(n1780), .IN3(n1781), .QN(\CARRYB[7][9] )
         );
  XOR3X1 U2931 ( .IN1(\ab[28][3] ), .IN2(\CARRYB[27][3] ), .IN3(\SUMB[27][4] ), 
        .Q(\SUMB[28][3] ) );
  NAND2X0 U2932 ( .IN1(\ab[28][3] ), .IN2(\CARRYB[27][3] ), .QN(n1783) );
  NAND2X1 U2933 ( .IN1(\ab[28][3] ), .IN2(\SUMB[27][4] ), .QN(n1784) );
  NAND2X0 U2934 ( .IN1(\CARRYB[27][3] ), .IN2(\SUMB[27][4] ), .QN(n1785) );
  XOR2X1 U2935 ( .IN1(\ab[29][3] ), .IN2(\SUMB[28][4] ), .Q(n1786) );
  NAND2X0 U2936 ( .IN1(\ab[29][3] ), .IN2(\SUMB[28][4] ), .QN(n1787) );
  NAND2X0 U2937 ( .IN1(\ab[29][3] ), .IN2(\CARRYB[28][3] ), .QN(n1788) );
  NAND2X0 U2938 ( .IN1(\SUMB[28][4] ), .IN2(\CARRYB[28][3] ), .QN(n1789) );
  XOR2X1 U2939 ( .IN1(\ab[27][3] ), .IN2(\SUMB[26][4] ), .Q(n1790) );
  XOR2X1 U2940 ( .IN1(n1790), .IN2(\CARRYB[26][3] ), .Q(\SUMB[27][3] ) );
  NAND2X0 U2941 ( .IN1(\CARRYB[26][3] ), .IN2(\SUMB[26][4] ), .QN(n1791) );
  NAND2X0 U2942 ( .IN1(\CARRYB[26][3] ), .IN2(\ab[27][3] ), .QN(n1792) );
  NAND2X1 U2943 ( .IN1(\SUMB[26][4] ), .IN2(\ab[27][3] ), .QN(n1793) );
  NAND2X0 U2944 ( .IN1(\ab[15][3] ), .IN2(\CARRYB[14][3] ), .QN(n1794) );
  NAND2X1 U2945 ( .IN1(\ab[15][3] ), .IN2(\SUMB[14][4] ), .QN(n1795) );
  NAND2X0 U2946 ( .IN1(\CARRYB[14][3] ), .IN2(\SUMB[14][4] ), .QN(n1796) );
  XOR2X1 U2947 ( .IN1(\ab[16][3] ), .IN2(\SUMB[15][4] ), .Q(n1797) );
  NAND2X0 U2948 ( .IN1(\ab[16][3] ), .IN2(\SUMB[15][4] ), .QN(n1798) );
  NAND2X0 U2949 ( .IN1(\ab[16][3] ), .IN2(\CARRYB[15][3] ), .QN(n1799) );
  NAND2X0 U2950 ( .IN1(\SUMB[15][4] ), .IN2(\CARRYB[15][3] ), .QN(n1800) );
  XOR3X1 U2951 ( .IN1(\ab[17][3] ), .IN2(\CARRYB[16][3] ), .IN3(\SUMB[16][4] ), 
        .Q(\SUMB[17][3] ) );
  NAND2X1 U2952 ( .IN1(\ab[17][3] ), .IN2(\CARRYB[16][3] ), .QN(n1801) );
  NAND2X0 U2953 ( .IN1(\ab[17][3] ), .IN2(\SUMB[16][4] ), .QN(n1802) );
  NAND2X0 U2954 ( .IN1(\CARRYB[16][3] ), .IN2(\SUMB[16][4] ), .QN(n1803) );
  XOR2X1 U2955 ( .IN1(\ab[18][3] ), .IN2(\SUMB[17][4] ), .Q(n1804) );
  XOR2X2 U2956 ( .IN1(n1804), .IN2(\CARRYB[17][3] ), .Q(\SUMB[18][3] ) );
  NAND2X0 U2957 ( .IN1(\ab[18][3] ), .IN2(\SUMB[17][4] ), .QN(n1805) );
  NAND2X0 U2958 ( .IN1(\ab[18][3] ), .IN2(\CARRYB[17][3] ), .QN(n1806) );
  NAND2X0 U2959 ( .IN1(\SUMB[17][4] ), .IN2(\CARRYB[17][3] ), .QN(n1807) );
  NAND3X1 U2960 ( .IN1(n1805), .IN2(n1806), .IN3(n1807), .QN(\CARRYB[18][3] )
         );
  XOR2X1 U2961 ( .IN1(n1812), .IN2(\CARRYB[25][4] ), .Q(\SUMB[26][4] ) );
  XOR3X1 U2962 ( .IN1(\ab[25][4] ), .IN2(\CARRYB[24][4] ), .IN3(\SUMB[24][5] ), 
        .Q(\SUMB[25][4] ) );
  NAND2X0 U2963 ( .IN1(\ab[25][4] ), .IN2(\CARRYB[24][4] ), .QN(n1809) );
  NAND2X1 U2964 ( .IN1(\ab[25][4] ), .IN2(\SUMB[24][5] ), .QN(n1810) );
  NAND2X0 U2965 ( .IN1(\CARRYB[24][4] ), .IN2(\SUMB[24][5] ), .QN(n1811) );
  XOR2X1 U2966 ( .IN1(\ab[26][4] ), .IN2(\SUMB[25][5] ), .Q(n1812) );
  NAND2X0 U2967 ( .IN1(\ab[26][4] ), .IN2(\SUMB[25][5] ), .QN(n1813) );
  NAND2X0 U2968 ( .IN1(\ab[26][4] ), .IN2(\CARRYB[25][4] ), .QN(n1814) );
  NAND2X0 U2969 ( .IN1(\SUMB[25][5] ), .IN2(\CARRYB[25][4] ), .QN(n1815) );
  XOR3X1 U2970 ( .IN1(\ab[20][4] ), .IN2(\CARRYB[19][4] ), .IN3(\SUMB[19][5] ), 
        .Q(\SUMB[20][4] ) );
  NAND2X0 U2971 ( .IN1(\ab[20][4] ), .IN2(\CARRYB[19][4] ), .QN(n1816) );
  NAND2X1 U2972 ( .IN1(\ab[20][4] ), .IN2(\SUMB[19][5] ), .QN(n1817) );
  NAND2X0 U2973 ( .IN1(\SUMB[19][5] ), .IN2(\CARRYB[19][4] ), .QN(n1818) );
  NAND3X1 U2974 ( .IN1(n1816), .IN2(n1817), .IN3(n1818), .QN(\CARRYB[20][4] )
         );
  NAND2X0 U2975 ( .IN1(\ab[21][4] ), .IN2(\SUMB[20][5] ), .QN(n1819) );
  NAND2X0 U2976 ( .IN1(\ab[21][4] ), .IN2(\CARRYB[20][4] ), .QN(n1820) );
  NAND2X0 U2977 ( .IN1(\SUMB[20][5] ), .IN2(\CARRYB[20][4] ), .QN(n1821) );
  NAND3X1 U2978 ( .IN1(n1819), .IN2(n1820), .IN3(n1821), .QN(\CARRYB[21][4] )
         );
  XOR2X1 U2979 ( .IN1(\ab[19][4] ), .IN2(\SUMB[18][5] ), .Q(n1822) );
  XOR2X1 U2980 ( .IN1(n1822), .IN2(\CARRYB[18][4] ), .Q(\SUMB[19][4] ) );
  NAND2X0 U2981 ( .IN1(\CARRYB[18][4] ), .IN2(\SUMB[18][5] ), .QN(n1823) );
  NAND2X0 U2982 ( .IN1(\CARRYB[18][4] ), .IN2(\ab[19][4] ), .QN(n1824) );
  NAND2X1 U2983 ( .IN1(\SUMB[18][5] ), .IN2(\ab[19][4] ), .QN(n1825) );
  NAND3X1 U2984 ( .IN1(n1823), .IN2(n1824), .IN3(n1825), .QN(\CARRYB[19][4] )
         );
  XOR3X1 U2985 ( .IN1(\ab[11][4] ), .IN2(\CARRYB[10][4] ), .IN3(\SUMB[10][5] ), 
        .Q(\SUMB[11][4] ) );
  NAND2X0 U2986 ( .IN1(\ab[11][4] ), .IN2(\CARRYB[10][4] ), .QN(n1826) );
  NAND2X1 U2987 ( .IN1(\ab[11][4] ), .IN2(\SUMB[10][5] ), .QN(n1827) );
  NAND2X0 U2988 ( .IN1(\CARRYB[10][4] ), .IN2(\SUMB[10][5] ), .QN(n1828) );
  XOR2X1 U2989 ( .IN1(\ab[12][4] ), .IN2(\SUMB[11][5] ), .Q(n1829) );
  NAND2X0 U2990 ( .IN1(\ab[12][4] ), .IN2(\SUMB[11][5] ), .QN(n1830) );
  NAND2X0 U2991 ( .IN1(\ab[12][4] ), .IN2(\CARRYB[11][4] ), .QN(n1831) );
  NAND2X0 U2992 ( .IN1(\SUMB[11][5] ), .IN2(\CARRYB[11][4] ), .QN(n1832) );
  NAND3X1 U2993 ( .IN1(n1830), .IN2(n1831), .IN3(n1832), .QN(\CARRYB[12][4] )
         );
  XOR3X1 U2994 ( .IN1(\CARRYB[30][8] ), .IN2(\ab[31][8] ), .IN3(\SUMB[30][9] ), 
        .Q(\SUMB[31][8] ) );
  NAND2X0 U2995 ( .IN1(\CARRYB[30][8] ), .IN2(\SUMB[30][9] ), .QN(n1833) );
  NAND2X0 U2996 ( .IN1(\CARRYB[30][8] ), .IN2(\ab[31][8] ), .QN(n1834) );
  XOR3X1 U2997 ( .IN1(\CARRYB[29][8] ), .IN2(\ab[30][8] ), .IN3(\SUMB[29][9] ), 
        .Q(\SUMB[30][8] ) );
  NAND2X0 U2998 ( .IN1(\CARRYB[29][8] ), .IN2(\SUMB[29][9] ), .QN(n1836) );
  NAND2X0 U2999 ( .IN1(\CARRYB[29][8] ), .IN2(\ab[30][8] ), .QN(n1837) );
  NAND2X0 U3000 ( .IN1(\SUMB[29][9] ), .IN2(\ab[30][8] ), .QN(n1838) );
  XOR3X1 U3001 ( .IN1(\ab[22][8] ), .IN2(\CARRYB[21][8] ), .IN3(\SUMB[21][9] ), 
        .Q(\SUMB[22][8] ) );
  NAND2X0 U3002 ( .IN1(\ab[22][8] ), .IN2(\CARRYB[21][8] ), .QN(n1839) );
  NAND2X1 U3003 ( .IN1(\ab[22][8] ), .IN2(\SUMB[21][9] ), .QN(n1840) );
  NAND2X0 U3004 ( .IN1(\CARRYB[21][8] ), .IN2(\SUMB[21][9] ), .QN(n1841) );
  NAND3X1 U3005 ( .IN1(n1839), .IN2(n1840), .IN3(n1841), .QN(\CARRYB[22][8] )
         );
  XOR2X1 U3006 ( .IN1(\ab[23][8] ), .IN2(\SUMB[22][9] ), .Q(n1842) );
  NAND2X0 U3007 ( .IN1(\ab[23][8] ), .IN2(\SUMB[22][9] ), .QN(n1843) );
  NAND2X0 U3008 ( .IN1(\ab[23][8] ), .IN2(\CARRYB[22][8] ), .QN(n1844) );
  NAND2X0 U3009 ( .IN1(\SUMB[22][9] ), .IN2(\CARRYB[22][8] ), .QN(n1845) );
  XOR3X1 U3010 ( .IN1(\ab[12][8] ), .IN2(\CARRYB[11][8] ), .IN3(\SUMB[11][9] ), 
        .Q(\SUMB[12][8] ) );
  NAND2X0 U3011 ( .IN1(\ab[12][8] ), .IN2(\CARRYB[11][8] ), .QN(n1846) );
  NAND2X0 U3012 ( .IN1(\CARRYB[11][8] ), .IN2(\SUMB[11][9] ), .QN(n1848) );
  NAND3X1 U3013 ( .IN1(n1846), .IN2(n1847), .IN3(n1848), .QN(\CARRYB[12][8] )
         );
  XOR2X1 U3014 ( .IN1(\ab[13][8] ), .IN2(\SUMB[12][9] ), .Q(n1849) );
  XOR2X2 U3015 ( .IN1(n1849), .IN2(\CARRYB[12][8] ), .Q(\SUMB[13][8] ) );
  NAND2X0 U3016 ( .IN1(\ab[13][8] ), .IN2(\SUMB[12][9] ), .QN(n1850) );
  NAND2X0 U3017 ( .IN1(\ab[13][8] ), .IN2(\CARRYB[12][8] ), .QN(n1851) );
  NAND2X0 U3018 ( .IN1(\SUMB[12][9] ), .IN2(\CARRYB[12][8] ), .QN(n1852) );
  NAND3X1 U3019 ( .IN1(n1850), .IN2(n1851), .IN3(n1852), .QN(\CARRYB[13][8] )
         );
  NAND2X0 U3020 ( .IN1(\ab[14][1] ), .IN2(\CARRYB[13][1] ), .QN(n1853) );
  NAND2X0 U3021 ( .IN1(\ab[14][1] ), .IN2(\SUMB[13][2] ), .QN(n1854) );
  NAND2X0 U3022 ( .IN1(\CARRYB[13][1] ), .IN2(\SUMB[13][2] ), .QN(n1855) );
  NAND3X1 U3023 ( .IN1(n1853), .IN2(n1854), .IN3(n1855), .QN(\CARRYB[14][1] )
         );
  XOR2X1 U3024 ( .IN1(n1856), .IN2(\CARRYB[14][1] ), .Q(\SUMB[15][1] ) );
  NAND2X0 U3025 ( .IN1(\ab[15][1] ), .IN2(\SUMB[14][2] ), .QN(n1857) );
  NAND2X0 U3026 ( .IN1(\ab[15][1] ), .IN2(\CARRYB[14][1] ), .QN(n1858) );
  NAND2X0 U3027 ( .IN1(\SUMB[14][2] ), .IN2(\CARRYB[14][1] ), .QN(n1859) );
  NAND3X1 U3028 ( .IN1(n1857), .IN2(n1858), .IN3(n1859), .QN(\CARRYB[15][1] )
         );
  XOR3X1 U3029 ( .IN1(\CARRYB[11][1] ), .IN2(\ab[12][1] ), .IN3(\SUMB[11][2] ), 
        .Q(\SUMB[12][1] ) );
  NAND2X0 U3030 ( .IN1(\CARRYB[11][1] ), .IN2(\SUMB[11][2] ), .QN(n1860) );
  NAND2X0 U3031 ( .IN1(\CARRYB[11][1] ), .IN2(\ab[12][1] ), .QN(n1861) );
  NAND2X1 U3032 ( .IN1(\SUMB[11][2] ), .IN2(\ab[12][1] ), .QN(n1862) );
  NAND3X0 U3033 ( .IN1(n1860), .IN2(n1861), .IN3(n1862), .QN(\CARRYB[12][1] )
         );
  XOR3X1 U3034 ( .IN1(\CARRYB[9][1] ), .IN2(\ab[10][1] ), .IN3(\SUMB[9][2] ), 
        .Q(\SUMB[10][1] ) );
  NAND2X0 U3035 ( .IN1(\CARRYB[9][1] ), .IN2(\SUMB[9][2] ), .QN(n1863) );
  NAND2X0 U3036 ( .IN1(\CARRYB[9][1] ), .IN2(\ab[10][1] ), .QN(n1864) );
  NAND2X1 U3037 ( .IN1(\SUMB[9][2] ), .IN2(\ab[10][1] ), .QN(n1865) );
  NAND3X0 U3038 ( .IN1(n1863), .IN2(n1864), .IN3(n1865), .QN(\CARRYB[10][1] )
         );
  XOR2X1 U3039 ( .IN1(\ab[11][1] ), .IN2(\CARRYB[10][1] ), .Q(n1866) );
  XOR2X1 U3040 ( .IN1(n1866), .IN2(\SUMB[10][2] ), .Q(\SUMB[11][1] ) );
  NAND2X0 U3041 ( .IN1(\SUMB[10][2] ), .IN2(\CARRYB[10][1] ), .QN(n1867) );
  NAND2X0 U3042 ( .IN1(\SUMB[10][2] ), .IN2(\ab[11][1] ), .QN(n1868) );
  NAND2X1 U3043 ( .IN1(\CARRYB[10][1] ), .IN2(\ab[11][1] ), .QN(n1869) );
  XOR3X1 U3044 ( .IN1(\CARRYB[8][10] ), .IN2(\ab[9][10] ), .IN3(\SUMB[8][11] ), 
        .Q(\SUMB[9][10] ) );
  NAND2X0 U3045 ( .IN1(\ab[9][10] ), .IN2(\CARRYB[8][10] ), .QN(n1870) );
  NAND2X1 U3046 ( .IN1(\ab[9][10] ), .IN2(\SUMB[8][11] ), .QN(n1871) );
  NAND2X0 U3047 ( .IN1(\SUMB[8][11] ), .IN2(\CARRYB[8][10] ), .QN(n1872) );
  NAND3X1 U3048 ( .IN1(n1872), .IN2(n1871), .IN3(n1870), .QN(\CARRYB[9][10] )
         );
  XOR2X1 U3049 ( .IN1(\ab[10][10] ), .IN2(\SUMB[9][11] ), .Q(n1873) );
  XOR2X2 U3050 ( .IN1(n1873), .IN2(\CARRYB[9][10] ), .Q(\SUMB[10][10] ) );
  NAND2X0 U3051 ( .IN1(\ab[10][10] ), .IN2(\SUMB[9][11] ), .QN(n1874) );
  NAND2X0 U3052 ( .IN1(\ab[10][10] ), .IN2(\CARRYB[9][10] ), .QN(n1875) );
  NAND2X0 U3053 ( .IN1(\SUMB[9][11] ), .IN2(\CARRYB[9][10] ), .QN(n1876) );
  NAND3X1 U3054 ( .IN1(n1875), .IN2(n1874), .IN3(n1876), .QN(\CARRYB[10][10] )
         );
  XOR3X1 U3055 ( .IN1(\CARRYB[6][10] ), .IN2(\ab[7][10] ), .IN3(\SUMB[6][11] ), 
        .Q(\SUMB[7][10] ) );
  NAND2X0 U3056 ( .IN1(\CARRYB[6][10] ), .IN2(\SUMB[6][11] ), .QN(n1877) );
  NAND2X0 U3057 ( .IN1(\CARRYB[6][10] ), .IN2(\ab[7][10] ), .QN(n1878) );
  NAND2X1 U3058 ( .IN1(\SUMB[6][11] ), .IN2(\ab[7][10] ), .QN(n1879) );
  NAND3X0 U3059 ( .IN1(n1877), .IN2(n1878), .IN3(n1879), .QN(\CARRYB[7][10] )
         );
  XOR3X1 U3060 ( .IN1(\CARRYB[27][12] ), .IN2(\ab[28][12] ), .IN3(
        \SUMB[27][13] ), .Q(\SUMB[28][12] ) );
  NAND2X1 U3061 ( .IN1(\CARRYB[27][12] ), .IN2(\SUMB[27][13] ), .QN(n1880) );
  NAND2X1 U3062 ( .IN1(\CARRYB[27][12] ), .IN2(\ab[28][12] ), .QN(n1881) );
  NAND2X1 U3063 ( .IN1(\SUMB[27][13] ), .IN2(\ab[28][12] ), .QN(n1882) );
  NAND3X0 U3064 ( .IN1(n1880), .IN2(n1881), .IN3(n1882), .QN(\CARRYB[28][12] )
         );
  XOR3X1 U3065 ( .IN1(\ab[29][12] ), .IN2(\CARRYB[28][12] ), .IN3(
        \SUMB[28][13] ), .Q(\SUMB[29][12] ) );
  NAND2X1 U3066 ( .IN1(\ab[29][12] ), .IN2(\CARRYB[28][12] ), .QN(n1883) );
  NAND2X0 U3067 ( .IN1(\ab[29][12] ), .IN2(\SUMB[28][13] ), .QN(n1884) );
  NAND2X0 U3068 ( .IN1(\CARRYB[28][12] ), .IN2(\SUMB[28][13] ), .QN(n1885) );
  XOR2X1 U3069 ( .IN1(\ab[30][12] ), .IN2(\SUMB[29][13] ), .Q(n1886) );
  NAND2X0 U3070 ( .IN1(\ab[30][12] ), .IN2(\SUMB[29][13] ), .QN(n1887) );
  NAND2X0 U3071 ( .IN1(\ab[30][12] ), .IN2(\CARRYB[29][12] ), .QN(n1888) );
  NAND2X0 U3072 ( .IN1(\SUMB[29][13] ), .IN2(\CARRYB[29][12] ), .QN(n1889) );
  XOR3X1 U3073 ( .IN1(\CARRYB[16][12] ), .IN2(\ab[17][12] ), .IN3(
        \SUMB[16][13] ), .Q(\SUMB[17][12] ) );
  NAND2X1 U3074 ( .IN1(\CARRYB[16][12] ), .IN2(\ab[17][12] ), .QN(n1891) );
  XOR3X1 U3075 ( .IN1(\ab[18][12] ), .IN2(\CARRYB[17][12] ), .IN3(
        \SUMB[17][13] ), .Q(\SUMB[18][12] ) );
  NAND2X1 U3076 ( .IN1(\ab[18][12] ), .IN2(\CARRYB[17][12] ), .QN(n1893) );
  NAND2X0 U3077 ( .IN1(\ab[18][12] ), .IN2(\SUMB[17][13] ), .QN(n1894) );
  NAND2X0 U3078 ( .IN1(\CARRYB[17][12] ), .IN2(\SUMB[17][13] ), .QN(n1895) );
  NAND3X1 U3079 ( .IN1(n1893), .IN2(n1894), .IN3(n1895), .QN(\CARRYB[18][12] )
         );
  NAND2X0 U3080 ( .IN1(\ab[19][12] ), .IN2(\SUMB[18][13] ), .QN(n1896) );
  NAND2X0 U3081 ( .IN1(\ab[19][12] ), .IN2(\CARRYB[18][12] ), .QN(n1897) );
  NAND2X0 U3082 ( .IN1(\SUMB[18][13] ), .IN2(\CARRYB[18][12] ), .QN(n1898) );
  XOR2X2 U3083 ( .IN1(n1899), .IN2(\ab[2][12] ), .Q(\SUMB[2][12] ) );
  NAND2X1 U3084 ( .IN1(\ab[2][12] ), .IN2(n9), .QN(n1900) );
  NAND2X0 U3085 ( .IN1(\ab[2][12] ), .IN2(\SUMB[1][13] ), .QN(n1901) );
  DELLN1X2 U3086 ( .INP(n2227), .Z(n1903) );
  DELLN1X2 U3087 ( .INP(n2227), .Z(n1904) );
  XOR2X2 U3088 ( .IN1(\ab[1][13] ), .IN2(\ab[0][14] ), .Q(\SUMB[1][13] ) );
  XOR3X1 U3089 ( .IN1(\ab[28][5] ), .IN2(\CARRYB[27][5] ), .IN3(\SUMB[27][6] ), 
        .Q(\SUMB[28][5] ) );
  NAND2X0 U3090 ( .IN1(\ab[28][5] ), .IN2(\CARRYB[27][5] ), .QN(n1905) );
  NAND2X1 U3091 ( .IN1(\ab[28][5] ), .IN2(\SUMB[27][6] ), .QN(n1906) );
  NAND2X0 U3092 ( .IN1(\CARRYB[27][5] ), .IN2(\SUMB[27][6] ), .QN(n1907) );
  XOR2X1 U3093 ( .IN1(\ab[29][5] ), .IN2(\SUMB[28][6] ), .Q(n1908) );
  NAND2X0 U3094 ( .IN1(\ab[29][5] ), .IN2(\SUMB[28][6] ), .QN(n1909) );
  NAND2X0 U3095 ( .IN1(\ab[29][5] ), .IN2(\CARRYB[28][5] ), .QN(n1910) );
  NAND2X0 U3096 ( .IN1(\SUMB[28][6] ), .IN2(\CARRYB[28][5] ), .QN(n1911) );
  XOR3X1 U3097 ( .IN1(\ab[18][5] ), .IN2(\CARRYB[17][5] ), .IN3(\SUMB[17][6] ), 
        .Q(\SUMB[18][5] ) );
  NAND2X0 U3098 ( .IN1(\ab[18][5] ), .IN2(\CARRYB[17][5] ), .QN(n1912) );
  NAND2X0 U3099 ( .IN1(\CARRYB[17][5] ), .IN2(\SUMB[17][6] ), .QN(n1914) );
  NAND3X1 U3100 ( .IN1(n1912), .IN2(n1913), .IN3(n1914), .QN(\CARRYB[18][5] )
         );
  XOR2X1 U3101 ( .IN1(\ab[19][5] ), .IN2(\SUMB[18][6] ), .Q(n1915) );
  XOR2X2 U3102 ( .IN1(n1915), .IN2(\CARRYB[18][5] ), .Q(\SUMB[19][5] ) );
  NAND2X0 U3103 ( .IN1(\ab[19][5] ), .IN2(\SUMB[18][6] ), .QN(n1916) );
  NAND2X0 U3104 ( .IN1(\ab[19][5] ), .IN2(\CARRYB[18][5] ), .QN(n1917) );
  NAND2X0 U3105 ( .IN1(\SUMB[18][6] ), .IN2(\CARRYB[18][5] ), .QN(n1918) );
  XOR3X1 U3106 ( .IN1(\ab[8][5] ), .IN2(\CARRYB[7][5] ), .IN3(\SUMB[7][6] ), 
        .Q(\SUMB[8][5] ) );
  NAND2X0 U3107 ( .IN1(\ab[8][5] ), .IN2(\CARRYB[7][5] ), .QN(n1919) );
  NAND2X1 U3108 ( .IN1(\ab[8][5] ), .IN2(\SUMB[7][6] ), .QN(n1920) );
  NAND2X0 U3109 ( .IN1(\CARRYB[7][5] ), .IN2(\SUMB[7][6] ), .QN(n1921) );
  NAND3X1 U3110 ( .IN1(n1919), .IN2(n1920), .IN3(n1921), .QN(\CARRYB[8][5] )
         );
  XOR2X1 U3111 ( .IN1(\ab[9][5] ), .IN2(\SUMB[8][6] ), .Q(n1922) );
  NAND2X0 U3112 ( .IN1(\ab[9][5] ), .IN2(\SUMB[8][6] ), .QN(n1923) );
  NAND2X0 U3113 ( .IN1(\ab[9][5] ), .IN2(\CARRYB[8][5] ), .QN(n1924) );
  NAND2X0 U3114 ( .IN1(\CARRYB[8][5] ), .IN2(\SUMB[8][6] ), .QN(n1925) );
  NAND3X1 U3115 ( .IN1(n1923), .IN2(n1924), .IN3(n1925), .QN(\CARRYB[9][5] )
         );
  NAND2X0 U3116 ( .IN1(\CARRYB[22][2] ), .IN2(\SUMB[22][3] ), .QN(n1926) );
  NAND2X0 U3117 ( .IN1(\CARRYB[22][2] ), .IN2(\ab[23][2] ), .QN(n1927) );
  NAND2X1 U3118 ( .IN1(\SUMB[22][3] ), .IN2(\ab[23][2] ), .QN(n1928) );
  NAND3X0 U3119 ( .IN1(n1926), .IN2(n1927), .IN3(n1928), .QN(\CARRYB[23][2] )
         );
  XOR3X1 U3120 ( .IN1(\ab[24][2] ), .IN2(\CARRYB[23][2] ), .IN3(\SUMB[23][3] ), 
        .Q(\SUMB[24][2] ) );
  NAND2X1 U3121 ( .IN1(\ab[24][2] ), .IN2(\CARRYB[23][2] ), .QN(n1929) );
  NAND2X0 U3122 ( .IN1(\ab[24][2] ), .IN2(\SUMB[23][3] ), .QN(n1930) );
  NAND2X0 U3123 ( .IN1(\CARRYB[23][2] ), .IN2(\SUMB[23][3] ), .QN(n1931) );
  XOR2X1 U3124 ( .IN1(\ab[25][2] ), .IN2(\SUMB[24][3] ), .Q(n1932) );
  NAND2X0 U3125 ( .IN1(\ab[25][2] ), .IN2(\SUMB[24][3] ), .QN(n1933) );
  NAND2X0 U3126 ( .IN1(\ab[25][2] ), .IN2(\CARRYB[24][2] ), .QN(n1934) );
  NAND2X0 U3127 ( .IN1(\SUMB[24][3] ), .IN2(\CARRYB[24][2] ), .QN(n1935) );
  XOR3X1 U3128 ( .IN1(\CARRYB[13][2] ), .IN2(\ab[14][2] ), .IN3(\SUMB[13][3] ), 
        .Q(\SUMB[14][2] ) );
  NAND2X0 U3129 ( .IN1(\CARRYB[13][2] ), .IN2(\SUMB[13][3] ), .QN(n1936) );
  NAND2X0 U3130 ( .IN1(\CARRYB[13][2] ), .IN2(\ab[14][2] ), .QN(n1937) );
  NAND2X1 U3131 ( .IN1(\SUMB[13][3] ), .IN2(\ab[14][2] ), .QN(n1938) );
  NAND3X0 U3132 ( .IN1(n1936), .IN2(n1937), .IN3(n1938), .QN(\CARRYB[14][2] )
         );
  XOR3X1 U3133 ( .IN1(\ab[15][2] ), .IN2(\CARRYB[14][2] ), .IN3(\SUMB[14][3] ), 
        .Q(\SUMB[15][2] ) );
  NAND2X1 U3134 ( .IN1(\ab[15][2] ), .IN2(\CARRYB[14][2] ), .QN(n1939) );
  NAND2X0 U3135 ( .IN1(\ab[15][2] ), .IN2(\SUMB[14][3] ), .QN(n1940) );
  NAND2X0 U3136 ( .IN1(\CARRYB[14][2] ), .IN2(\SUMB[14][3] ), .QN(n1941) );
  NAND3X1 U3137 ( .IN1(n1939), .IN2(n1940), .IN3(n1941), .QN(\CARRYB[15][2] )
         );
  NAND2X0 U3138 ( .IN1(\ab[16][2] ), .IN2(\SUMB[15][3] ), .QN(n1942) );
  NAND2X0 U3139 ( .IN1(\ab[16][2] ), .IN2(\CARRYB[15][2] ), .QN(n1943) );
  NAND2X0 U3140 ( .IN1(\SUMB[15][3] ), .IN2(\CARRYB[15][2] ), .QN(n1944) );
  DELLN1X2 U3141 ( .INP(n2237), .Z(n1945) );
  DELLN1X2 U3142 ( .INP(n2237), .Z(n1946) );
  XOR2X1 U3143 ( .IN1(ZA), .IN2(n148), .Q(n1947) );
  XOR2X1 U3144 ( .IN1(n1947), .IN2(\SUMB[31][0] ), .Q(\A1[29] ) );
  NAND2X0 U3145 ( .IN1(\ab[31][0] ), .IN2(\CARRYB[30][0] ), .QN(n1948) );
  NAND2X0 U3146 ( .IN1(\ab[31][0] ), .IN2(\SUMB[30][1] ), .QN(n1949) );
  NAND2X0 U3147 ( .IN1(\CARRYB[30][0] ), .IN2(\SUMB[30][1] ), .QN(n1950) );
  NAND3X1 U3148 ( .IN1(n1948), .IN2(n1949), .IN3(n1950), .QN(\CARRYB[31][0] )
         );
  NAND2X0 U3149 ( .IN1(ZA), .IN2(n148), .QN(n1951) );
  NAND2X0 U3150 ( .IN1(ZA), .IN2(\SUMB[31][0] ), .QN(n1952) );
  NAND2X0 U3151 ( .IN1(n148), .IN2(\SUMB[31][0] ), .QN(n1953) );
  NAND3X1 U3152 ( .IN1(n1951), .IN2(n1952), .IN3(n1953), .QN(\A2[30] ) );
  XOR3X1 U3153 ( .IN1(\ab[21][0] ), .IN2(\CARRYB[20][0] ), .IN3(\SUMB[20][1] ), 
        .Q(\A1[19] ) );
  NAND2X1 U3154 ( .IN1(\ab[21][0] ), .IN2(\SUMB[20][1] ), .QN(n1955) );
  XOR2X1 U3155 ( .IN1(\ab[22][0] ), .IN2(\SUMB[21][1] ), .Q(n1957) );
  XOR2X1 U3156 ( .IN1(n1957), .IN2(n197), .Q(\A1[20] ) );
  NAND2X0 U3157 ( .IN1(\ab[22][0] ), .IN2(\SUMB[21][1] ), .QN(n1958) );
  NAND2X0 U3158 ( .IN1(\ab[22][0] ), .IN2(\CARRYB[21][0] ), .QN(n1959) );
  NAND2X0 U3159 ( .IN1(\SUMB[21][1] ), .IN2(n197), .QN(n1960) );
  NAND3X1 U3160 ( .IN1(n1958), .IN2(n1959), .IN3(n1960), .QN(\CARRYB[22][0] )
         );
  XOR3X1 U3161 ( .IN1(\ab[9][0] ), .IN2(\CARRYB[8][0] ), .IN3(\SUMB[8][1] ), 
        .Q(\A1[7] ) );
  NAND2X1 U3162 ( .IN1(\ab[9][0] ), .IN2(\SUMB[8][1] ), .QN(n1962) );
  NAND3X1 U3163 ( .IN1(n1961), .IN2(n1962), .IN3(n1963), .QN(\CARRYB[9][0] )
         );
  XOR2X1 U3164 ( .IN1(\ab[10][0] ), .IN2(\SUMB[9][1] ), .Q(n1964) );
  XOR2X1 U3165 ( .IN1(n1964), .IN2(\CARRYB[9][0] ), .Q(\A1[8] ) );
  NAND2X0 U3166 ( .IN1(\ab[10][0] ), .IN2(\SUMB[9][1] ), .QN(n1965) );
  NAND2X0 U3167 ( .IN1(\ab[10][0] ), .IN2(\CARRYB[9][0] ), .QN(n1966) );
  NAND2X0 U3168 ( .IN1(\SUMB[9][1] ), .IN2(\CARRYB[9][0] ), .QN(n1967) );
  NAND2X0 U3169 ( .IN1(\CARRYB[29][0] ), .IN2(\SUMB[29][1] ), .QN(n1968) );
  NAND2X0 U3170 ( .IN1(\SUMB[29][1] ), .IN2(\ab[30][0] ), .QN(n1970) );
  NAND3X1 U3171 ( .IN1(n1968), .IN2(n1969), .IN3(n1970), .QN(\CARRYB[30][0] )
         );
  DELLN1X2 U3172 ( .INP(n2221), .Z(n2129) );
  DELLN1X2 U3173 ( .INP(n2225), .Z(n2141) );
  NBUFFX2 U3174 ( .INP(n2229), .Z(n2151) );
  DELLN1X2 U3175 ( .INP(n2205), .Z(n2089) );
  NBUFFX2 U3176 ( .INP(n2234), .Z(n2163) );
  DELLN1X2 U3177 ( .INP(n2225), .Z(n2140) );
  DELLN1X2 U3178 ( .INP(n2224), .Z(n2138) );
  DELLN1X2 U3179 ( .INP(n2223), .Z(n2135) );
  DELLN1X2 U3180 ( .INP(n2222), .Z(n2132) );
  NBUFFX2 U3181 ( .INP(n2237), .Z(n2169) );
  NBUFFX4 U3182 ( .INP(n2215), .Z(n2111) );
  NBUFFX4 U3183 ( .INP(n2214), .Z(n2108) );
  DELLN1X2 U3184 ( .INP(n2204), .Z(n2086) );
  DELLN1X2 U3185 ( .INP(n2203), .Z(n2083) );
  DELLN1X2 U3186 ( .INP(n2202), .Z(n2080) );
  DELLN1X2 U3187 ( .INP(n2201), .Z(n2077) );
  DELLN1X2 U3188 ( .INP(n2200), .Z(n2074) );
  DELLN1X2 U3189 ( .INP(n2199), .Z(n2071) );
  DELLN1X2 U3190 ( .INP(n2198), .Z(n2068) );
  INVX0 U3191 ( .INP(A[0]), .ZN(n1971) );
  NBUFFX4 U3192 ( .INP(n2233), .Z(n2161) );
  AND2X1 U3193 ( .IN1(\CARRYB[31][11] ), .IN2(\SUMB[31][12] ), .Q(n1972) );
  AND2X1 U3194 ( .IN1(\CARRYB[31][6] ), .IN2(\SUMB[31][7] ), .Q(n1973) );
  AND2X1 U3195 ( .IN1(\CARRYB[31][3] ), .IN2(\SUMB[31][4] ), .Q(n1974) );
  AND2X1 U3196 ( .IN1(\CARRYB[31][7] ), .IN2(\SUMB[31][8] ), .Q(n1975) );
  AND2X1 U3197 ( .IN1(\CARRYB[31][5] ), .IN2(\SUMB[31][6] ), .Q(n1978) );
  AND2X1 U3198 ( .IN1(\CARRYB[31][13] ), .IN2(\SUMB[31][14] ), .Q(n1979) );
  AND2X1 U3199 ( .IN1(\CARRYB[31][14] ), .IN2(\SUMB[31][15] ), .Q(n1980) );
  AND2X1 U3200 ( .IN1(\CARRYB[31][4] ), .IN2(\SUMB[31][5] ), .Q(n1982) );
  AND2X1 U3201 ( .IN1(\CARRYB[31][12] ), .IN2(\SUMB[31][13] ), .Q(n1983) );
  AND2X1 U3202 ( .IN1(\CARRYB[31][0] ), .IN2(\SUMB[31][1] ), .Q(n1984) );
  AND2X1 U3203 ( .IN1(\CARRYB[31][10] ), .IN2(\SUMB[31][11] ), .Q(n1985) );
  AND2X1 U3204 ( .IN1(\CARRYB[31][2] ), .IN2(\SUMB[31][3] ), .Q(n1986) );
  NBUFFX2 U3205 ( .INP(n2221), .Z(n2130) );
  AND2X1 U3206 ( .IN1(\CARRYB[31][29] ), .IN2(\SUMB[31][30] ), .Q(n1987) );
  AND2X1 U3207 ( .IN1(\CARRYB[31][15] ), .IN2(\SUMB[31][16] ), .Q(n1988) );
  AND2X1 U3208 ( .IN1(\CARRYB[31][16] ), .IN2(\SUMB[31][17] ), .Q(n1989) );
  AND2X1 U3209 ( .IN1(\CARRYB[31][17] ), .IN2(\SUMB[31][18] ), .Q(n1990) );
  AND2X1 U3210 ( .IN1(\CARRYB[31][18] ), .IN2(\SUMB[31][19] ), .Q(n1991) );
  AND2X1 U3211 ( .IN1(\CARRYB[31][19] ), .IN2(\SUMB[31][20] ), .Q(n1992) );
  NBUFFX2 U3212 ( .INP(n2220), .Z(n2127) );
  NBUFFX2 U3213 ( .INP(n2215), .Z(n2112) );
  AND2X1 U3214 ( .IN1(\CARRYB[31][28] ), .IN2(\SUMB[31][29] ), .Q(n1994) );
  AND2X1 U3215 ( .IN1(\CARRYB[31][21] ), .IN2(\SUMB[31][22] ), .Q(n1995) );
  AND2X1 U3216 ( .IN1(\CARRYB[31][22] ), .IN2(\SUMB[31][23] ), .Q(n1996) );
  AND2X1 U3217 ( .IN1(\CARRYB[31][23] ), .IN2(\SUMB[31][24] ), .Q(n1997) );
  AND2X1 U3218 ( .IN1(\CARRYB[31][24] ), .IN2(\SUMB[31][25] ), .Q(n1998) );
  AND2X1 U3219 ( .IN1(\CARRYB[31][27] ), .IN2(\SUMB[31][28] ), .Q(n1999) );
  AND2X1 U3220 ( .IN1(\CARRYB[31][25] ), .IN2(\SUMB[31][26] ), .Q(n2000) );
  AND2X1 U3221 ( .IN1(\CARRYB[31][26] ), .IN2(\SUMB[31][27] ), .Q(n2001) );
  NBUFFX2 U3222 ( .INP(n2221), .Z(n2128) );
  NBUFFX2 U3223 ( .INP(n2220), .Z(n2125) );
  NBUFFX2 U3224 ( .INP(n2214), .Z(n2109) );
  NBUFFX2 U3225 ( .INP(n2215), .Z(n2110) );
  NBUFFX2 U3226 ( .INP(n2214), .Z(n2107) );
  NBUFFX2 U3227 ( .INP(n2204), .Z(n2087) );
  NBUFFX2 U3228 ( .INP(n2204), .Z(n2088) );
  NBUFFX2 U3229 ( .INP(n2203), .Z(n2084) );
  NBUFFX2 U3230 ( .INP(n2203), .Z(n2085) );
  NBUFFX2 U3231 ( .INP(n2202), .Z(n2081) );
  NBUFFX2 U3232 ( .INP(n2202), .Z(n2082) );
  NBUFFX2 U3233 ( .INP(n2201), .Z(n2078) );
  NBUFFX2 U3234 ( .INP(n2201), .Z(n2079) );
  NBUFFX2 U3235 ( .INP(n2200), .Z(n2075) );
  NBUFFX2 U3236 ( .INP(n2200), .Z(n2076) );
  NBUFFX2 U3237 ( .INP(n2199), .Z(n2072) );
  NBUFFX2 U3238 ( .INP(n2199), .Z(n2073) );
  NBUFFX2 U3239 ( .INP(n2198), .Z(n2069) );
  NBUFFX2 U3240 ( .INP(n2197), .Z(n2066) );
  NBUFFX2 U3241 ( .INP(n2198), .Z(n2070) );
  NBUFFX2 U3242 ( .INP(n2239), .Z(n2174) );
  NBUFFX2 U3243 ( .INP(n2197), .Z(n2065) );
  NBUFFX2 U3244 ( .INP(n2197), .Z(n2067) );
  NBUFFX2 U3245 ( .INP(n2196), .Z(n2062) );
  NBUFFX2 U3246 ( .INP(n2196), .Z(n2063) );
  NBUFFX2 U3247 ( .INP(n2196), .Z(n2064) );
  NBUFFX2 U3248 ( .INP(n2195), .Z(n2059) );
  NBUFFX2 U3249 ( .INP(n2195), .Z(n2060) );
  NBUFFX2 U3250 ( .INP(n2195), .Z(n2061) );
  NBUFFX2 U3251 ( .INP(n2194), .Z(n2056) );
  NBUFFX2 U3252 ( .INP(n2194), .Z(n2057) );
  NBUFFX2 U3253 ( .INP(n2194), .Z(n2058) );
  NBUFFX2 U3254 ( .INP(n2239), .Z(n2173) );
  NBUFFX2 U3255 ( .INP(n2229), .Z(n2150) );
  NBUFFX2 U3256 ( .INP(n2193), .Z(n2054) );
  NBUFFX2 U3257 ( .INP(n2193), .Z(n2053) );
  NBUFFX2 U3258 ( .INP(n2193), .Z(n2055) );
  NBUFFX2 U3259 ( .INP(n2192), .Z(n2050) );
  NBUFFX2 U3260 ( .INP(n2192), .Z(n2051) );
  NBUFFX2 U3261 ( .INP(n2192), .Z(n2052) );
  NBUFFX2 U3262 ( .INP(n2191), .Z(n2047) );
  NBUFFX2 U3263 ( .INP(n2191), .Z(n2048) );
  NBUFFX2 U3264 ( .INP(n2191), .Z(n2049) );
  NBUFFX2 U3265 ( .INP(n2190), .Z(n2044) );
  NBUFFX2 U3266 ( .INP(n2190), .Z(n2045) );
  NBUFFX2 U3267 ( .INP(n2190), .Z(n2046) );
  NBUFFX2 U3268 ( .INP(n2189), .Z(n2041) );
  NBUFFX2 U3269 ( .INP(n2189), .Z(n2042) );
  NBUFFX2 U3270 ( .INP(n2189), .Z(n2043) );
  NBUFFX2 U3271 ( .INP(n2188), .Z(n2038) );
  NBUFFX2 U3272 ( .INP(n2188), .Z(n2039) );
  NBUFFX2 U3273 ( .INP(n2188), .Z(n2040) );
  NBUFFX2 U3274 ( .INP(n2187), .Z(n2035) );
  NBUFFX2 U3275 ( .INP(n2187), .Z(n2036) );
  NBUFFX2 U3276 ( .INP(n2187), .Z(n2037) );
  NBUFFX2 U3277 ( .INP(n2186), .Z(n2032) );
  NBUFFX2 U3278 ( .INP(n2186), .Z(n2033) );
  NBUFFX2 U3279 ( .INP(n2186), .Z(n2034) );
  NBUFFX2 U3280 ( .INP(n2185), .Z(n2029) );
  NBUFFX2 U3281 ( .INP(n2185), .Z(n2030) );
  NBUFFX2 U3282 ( .INP(n2185), .Z(n2031) );
  NBUFFX2 U3283 ( .INP(n2184), .Z(n2027) );
  NBUFFX2 U3284 ( .INP(n2184), .Z(n2026) );
  NBUFFX2 U3285 ( .INP(n2184), .Z(n2028) );
  NBUFFX2 U3286 ( .INP(n2183), .Z(n2023) );
  NBUFFX2 U3287 ( .INP(n2183), .Z(n2024) );
  NBUFFX2 U3288 ( .INP(n2183), .Z(n2025) );
  NBUFFX2 U3289 ( .INP(n2182), .Z(n2020) );
  NBUFFX2 U3290 ( .INP(n2182), .Z(n2021) );
  NBUFFX2 U3291 ( .INP(n2182), .Z(n2022) );
  NBUFFX2 U3292 ( .INP(n2181), .Z(n2017) );
  NBUFFX2 U3293 ( .INP(n2181), .Z(n2018) );
  NBUFFX2 U3294 ( .INP(n2181), .Z(n2019) );
  NBUFFX2 U3295 ( .INP(n2180), .Z(n2014) );
  NBUFFX2 U3296 ( .INP(n2180), .Z(n2015) );
  NBUFFX2 U3297 ( .INP(n2180), .Z(n2016) );
  NBUFFX2 U3298 ( .INP(n2179), .Z(n2011) );
  NBUFFX2 U3299 ( .INP(n2179), .Z(n2012) );
  NBUFFX2 U3300 ( .INP(n2179), .Z(n2013) );
  NBUFFX2 U3301 ( .INP(n2178), .Z(n2008) );
  NBUFFX2 U3302 ( .INP(n2178), .Z(n2009) );
  NBUFFX2 U3303 ( .INP(n2178), .Z(n2010) );
  NBUFFX2 U3304 ( .INP(n2177), .Z(n2005) );
  NBUFFX2 U3305 ( .INP(n2177), .Z(n2006) );
  NBUFFX2 U3306 ( .INP(n2177), .Z(n2007) );
  INVX0 U3307 ( .INP(B[14]), .ZN(n2225) );
  INVX0 U3308 ( .INP(B[15]), .ZN(n2224) );
  INVX0 U3309 ( .INP(B[4]), .ZN(n2235) );
  INVX0 U3310 ( .INP(B[8]), .ZN(n2231) );
  INVX0 U3311 ( .INP(ZB), .ZN(n2208) );
  INVX0 U3312 ( .INP(B[16]), .ZN(n2223) );
  INVX0 U3313 ( .INP(B[17]), .ZN(n2222) );
  INVX0 U3314 ( .INP(B[18]), .ZN(n2221) );
  INVX0 U3315 ( .INP(B[19]), .ZN(n2220) );
  INVX0 U3316 ( .INP(B[20]), .ZN(n2219) );
  INVX0 U3317 ( .INP(B[21]), .ZN(n2218) );
  INVX0 U3318 ( .INP(A[2]), .ZN(n2205) );
  INVX0 U3319 ( .INP(B[22]), .ZN(n2217) );
  INVX0 U3320 ( .INP(B[23]), .ZN(n2216) );
  INVX0 U3321 ( .INP(B[24]), .ZN(n2215) );
  INVX0 U3322 ( .INP(B[25]), .ZN(n2214) );
  INVX0 U3323 ( .INP(B[26]), .ZN(n2213) );
  INVX0 U3324 ( .INP(B[27]), .ZN(n2212) );
  INVX0 U3325 ( .INP(B[28]), .ZN(n2211) );
  INVX0 U3326 ( .INP(B[29]), .ZN(n2210) );
  INVX0 U3327 ( .INP(B[30]), .ZN(n2209) );
  INVX0 U3328 ( .INP(A[3]), .ZN(n2204) );
  INVX0 U3329 ( .INP(A[4]), .ZN(n2203) );
  INVX0 U3330 ( .INP(A[5]), .ZN(n2202) );
  INVX0 U3331 ( .INP(A[6]), .ZN(n2201) );
  INVX0 U3332 ( .INP(A[7]), .ZN(n2200) );
  INVX0 U3333 ( .INP(A[8]), .ZN(n2199) );
  INVX0 U3334 ( .INP(A[9]), .ZN(n2198) );
  INVX0 U3335 ( .INP(A[10]), .ZN(n2197) );
  INVX0 U3336 ( .INP(A[11]), .ZN(n2196) );
  INVX0 U3337 ( .INP(A[12]), .ZN(n2195) );
  INVX0 U3338 ( .INP(A[13]), .ZN(n2194) );
  INVX0 U3339 ( .INP(A[14]), .ZN(n2193) );
  INVX0 U3340 ( .INP(A[15]), .ZN(n2192) );
  INVX0 U3341 ( .INP(A[16]), .ZN(n2191) );
  INVX0 U3342 ( .INP(A[17]), .ZN(n2190) );
  INVX0 U3343 ( .INP(A[18]), .ZN(n2189) );
  INVX0 U3344 ( .INP(A[19]), .ZN(n2188) );
  INVX0 U3345 ( .INP(A[20]), .ZN(n2187) );
  INVX0 U3346 ( .INP(A[21]), .ZN(n2186) );
  INVX0 U3347 ( .INP(A[22]), .ZN(n2185) );
  INVX0 U3348 ( .INP(A[23]), .ZN(n2184) );
  INVX0 U3349 ( .INP(A[24]), .ZN(n2183) );
  INVX0 U3350 ( .INP(A[25]), .ZN(n2182) );
  INVX0 U3351 ( .INP(A[26]), .ZN(n2181) );
  INVX0 U3352 ( .INP(A[27]), .ZN(n2180) );
  INVX0 U3353 ( .INP(A[28]), .ZN(n2179) );
  NBUFFX4 U3354 ( .INP(n2176), .Z(n2004) );
  INVX0 U3355 ( .INP(ZA), .ZN(n2176) );
  INVX0 U3356 ( .INP(A[29]), .ZN(n2178) );
  INVX0 U3357 ( .INP(A[30]), .ZN(n2177) );
  XOR2X1 U3358 ( .IN1(\CARRYB[31][0] ), .IN2(\SUMB[31][1] ), .Q(\A1[30] ) );
  XOR2X1 U3359 ( .IN1(\CARRYB[31][4] ), .IN2(\SUMB[31][5] ), .Q(\A1[34] ) );
  XOR2X1 U3360 ( .IN1(\CARRYB[31][5] ), .IN2(\SUMB[31][6] ), .Q(\A1[35] ) );
  XOR2X1 U3361 ( .IN1(\CARRYB[31][12] ), .IN2(\SUMB[31][13] ), .Q(\A1[42] ) );
  XOR2X1 U3362 ( .IN1(\CARRYB[31][13] ), .IN2(\SUMB[31][14] ), .Q(\A1[43] ) );
  XOR2X1 U3363 ( .IN1(\CARRYB[31][14] ), .IN2(\SUMB[31][15] ), .Q(\A1[44] ) );
  XOR2X1 U3364 ( .IN1(\CARRYB[31][15] ), .IN2(\SUMB[31][16] ), .Q(\A1[45] ) );
  XOR2X1 U3365 ( .IN1(\CARRYB[31][16] ), .IN2(\SUMB[31][17] ), .Q(\A1[46] ) );
  XOR2X1 U3366 ( .IN1(\CARRYB[31][17] ), .IN2(\SUMB[31][18] ), .Q(\A1[47] ) );
  XOR2X1 U3367 ( .IN1(\CARRYB[31][18] ), .IN2(\SUMB[31][19] ), .Q(\A1[48] ) );
  XOR2X1 U3368 ( .IN1(\CARRYB[31][19] ), .IN2(\SUMB[31][20] ), .Q(\A1[49] ) );
  XOR2X1 U3369 ( .IN1(\CARRYB[31][20] ), .IN2(\SUMB[31][21] ), .Q(\A1[50] ) );
  XOR2X1 U3370 ( .IN1(\CARRYB[31][21] ), .IN2(\SUMB[31][22] ), .Q(\A1[51] ) );
  XOR2X1 U3371 ( .IN1(\CARRYB[31][22] ), .IN2(\SUMB[31][23] ), .Q(\A1[52] ) );
  XOR2X1 U3372 ( .IN1(\CARRYB[31][23] ), .IN2(\SUMB[31][24] ), .Q(\A1[53] ) );
  XOR2X1 U3373 ( .IN1(\CARRYB[31][24] ), .IN2(\SUMB[31][25] ), .Q(\A1[54] ) );
  XOR2X1 U3374 ( .IN1(\CARRYB[31][25] ), .IN2(\SUMB[31][26] ), .Q(\A1[55] ) );
  XOR2X1 U3375 ( .IN1(\CARRYB[31][26] ), .IN2(\SUMB[31][27] ), .Q(\A1[56] ) );
  XOR2X1 U3376 ( .IN1(\CARRYB[31][27] ), .IN2(\SUMB[31][28] ), .Q(\A1[57] ) );
  XOR2X1 U3377 ( .IN1(\CARRYB[31][28] ), .IN2(\SUMB[31][29] ), .Q(\A1[58] ) );
  XOR2X1 U3378 ( .IN1(\CARRYB[31][29] ), .IN2(\SUMB[31][30] ), .Q(\A1[59] ) );
  XOR2X1 U3379 ( .IN1(\CARRYB[31][30] ), .IN2(\SUMB[31][31] ), .Q(\A1[60] ) );
  XOR2X1 U3380 ( .IN1(\ab[1][0] ), .IN2(\ab[0][1] ), .Q(PRODUCT[1]) );
  XOR2X1 U3381 ( .IN1(\ab[1][1] ), .IN2(\ab[0][2] ), .Q(\SUMB[1][1] ) );
  XOR2X1 U3382 ( .IN1(\ab[1][2] ), .IN2(\ab[0][3] ), .Q(\SUMB[1][2] ) );
  XOR2X1 U3383 ( .IN1(\ab[1][5] ), .IN2(\ab[0][6] ), .Q(\SUMB[1][5] ) );
  XOR2X1 U3384 ( .IN1(\ab[1][6] ), .IN2(\ab[0][7] ), .Q(\SUMB[1][6] ) );
  XOR2X1 U3385 ( .IN1(\ab[1][7] ), .IN2(\ab[0][8] ), .Q(\SUMB[1][7] ) );
  XOR2X1 U3386 ( .IN1(\ab[1][10] ), .IN2(\ab[0][11] ), .Q(\SUMB[1][10] ) );
  XOR2X1 U3387 ( .IN1(\ab[1][15] ), .IN2(\ab[0][16] ), .Q(\SUMB[1][15] ) );
  XOR2X1 U3388 ( .IN1(\ab[1][18] ), .IN2(\ab[0][19] ), .Q(\SUMB[1][18] ) );
  INVX0 U3389 ( .INP(B[9]), .ZN(n2230) );
  DELLN1X2 U3390 ( .INP(n2206), .Z(n2002) );
  DELLN1X2 U3391 ( .INP(n2206), .Z(n2003) );
  INVX0 U3392 ( .INP(B[13]), .ZN(n2226) );
  INVX0 U3393 ( .INP(A[0]), .ZN(n2207) );
  INVX0 U3394 ( .INP(B[12]), .ZN(n2227) );
  INVX0 U3395 ( .INP(B[10]), .ZN(n2229) );
  INVX0 U3396 ( .INP(B[6]), .ZN(n2233) );
  INVX0 U3397 ( .INP(B[5]), .ZN(n2234) );
  INVX0 U3398 ( .INP(B[11]), .ZN(n2228) );
  INVX0 U3399 ( .INP(B[7]), .ZN(n2232) );
  INVX0 U3400 ( .INP(B[0]), .ZN(n2239) );
  INVX0 U3401 ( .INP(B[3]), .ZN(n2236) );
  INVX0 U3402 ( .INP(B[1]), .ZN(n2238) );
  INVX0 U3403 ( .INP(A[1]), .ZN(n2206) );
  INVX0 U3404 ( .INP(B[2]), .ZN(n2237) );
  DELLN1X2 U3405 ( .INP(n1971), .Z(n2093) );
  DELLN1X2 U3406 ( .INP(n2226), .Z(n2143) );
  DELLN1X2 U3407 ( .INP(n2226), .Z(n2144) );
  DELLN1X2 U3408 ( .INP(n2226), .Z(n2145) );
  DELLN1X2 U3409 ( .INP(n2227), .Z(n2146) );
  DELLN1X2 U3410 ( .INP(n2229), .Z(n2149) );
  DELLN1X2 U3411 ( .INP(n2230), .Z(n2153) );
  DELLN1X2 U3412 ( .INP(n2232), .Z(n2158) );
  DELLN1X2 U3413 ( .INP(n2233), .Z(n2160) );
  DELLN1X2 U3414 ( .INP(n2234), .Z(n2162) );
  DELLN1X2 U3415 ( .INP(n2238), .Z(n2170) );
  DELLN1X2 U3416 ( .INP(n2239), .Z(n2172) );
  NOR2X0 U3417 ( .IN1(n2070), .IN2(n2152), .QN(\ab[9][9] ) );
  NOR2X0 U3418 ( .IN1(n2070), .IN2(n2155), .QN(\ab[9][8] ) );
  NOR2X0 U3419 ( .IN1(n2070), .IN2(n2158), .QN(\ab[9][7] ) );
  NOR2X0 U3420 ( .IN1(n2070), .IN2(n2160), .QN(\ab[9][6] ) );
  NOR2X0 U3421 ( .IN1(n2070), .IN2(n2162), .QN(\ab[9][5] ) );
  NOR2X0 U3422 ( .IN1(n2070), .IN2(n2164), .QN(\ab[9][4] ) );
  NOR2X0 U3423 ( .IN1(n2070), .IN2(n2168), .QN(\ab[9][3] ) );
  NOR2X0 U3424 ( .IN1(A[9]), .IN2(n2094), .QN(\ab[9][31] ) );
  NOR2X0 U3425 ( .IN1(n2069), .IN2(n2096), .QN(\ab[9][30] ) );
  NOR2X0 U3426 ( .IN1(n2069), .IN2(n2169), .QN(\ab[9][2] ) );
  NOR2X0 U3427 ( .IN1(n2069), .IN2(n580), .QN(\ab[9][29] ) );
  NOR2X0 U3428 ( .IN1(n2069), .IN2(n2099), .QN(\ab[9][28] ) );
  NOR2X0 U3429 ( .IN1(n2069), .IN2(n2101), .QN(\ab[9][27] ) );
  NOR2X0 U3430 ( .IN1(n2069), .IN2(n2106), .QN(\ab[9][26] ) );
  NOR2X0 U3431 ( .IN1(n2069), .IN2(n2107), .QN(\ab[9][25] ) );
  NOR2X0 U3432 ( .IN1(n2069), .IN2(n2110), .QN(\ab[9][24] ) );
  NOR2X0 U3433 ( .IN1(n2069), .IN2(n2114), .QN(\ab[9][23] ) );
  NOR2X0 U3434 ( .IN1(n2069), .IN2(n2117), .QN(\ab[9][22] ) );
  NOR2X0 U3435 ( .IN1(n2069), .IN2(n2119), .QN(\ab[9][21] ) );
  NOR2X0 U3436 ( .IN1(n2069), .IN2(n2123), .QN(\ab[9][20] ) );
  NOR2X0 U3437 ( .IN1(n2068), .IN2(n2170), .QN(\ab[9][1] ) );
  NOR2X0 U3438 ( .IN1(n2068), .IN2(n2125), .QN(\ab[9][19] ) );
  NOR2X0 U3439 ( .IN1(n2068), .IN2(n2128), .QN(\ab[9][18] ) );
  NOR2X0 U3440 ( .IN1(n2068), .IN2(n2131), .QN(\ab[9][17] ) );
  NOR2X0 U3441 ( .IN1(n2068), .IN2(n2134), .QN(\ab[9][16] ) );
  NOR2X0 U3442 ( .IN1(n2068), .IN2(n2137), .QN(\ab[9][15] ) );
  NOR2X0 U3443 ( .IN1(n2068), .IN2(n2140), .QN(\ab[9][14] ) );
  NOR2X0 U3444 ( .IN1(n2068), .IN2(n2143), .QN(\ab[9][13] ) );
  NOR2X0 U3445 ( .IN1(n2068), .IN2(n2146), .QN(\ab[9][12] ) );
  NOR2X0 U3446 ( .IN1(n2068), .IN2(n2148), .QN(\ab[9][11] ) );
  NOR2X0 U3447 ( .IN1(n2068), .IN2(n2149), .QN(\ab[9][10] ) );
  NOR2X0 U3448 ( .IN1(n2068), .IN2(n2172), .QN(\ab[9][0] ) );
  NOR2X0 U3449 ( .IN1(n2153), .IN2(n2073), .QN(\ab[8][9] ) );
  NOR2X0 U3450 ( .IN1(n2157), .IN2(n2073), .QN(\ab[8][8] ) );
  NOR2X0 U3451 ( .IN1(n2158), .IN2(n2073), .QN(\ab[8][7] ) );
  NOR2X0 U3452 ( .IN1(n2160), .IN2(n2073), .QN(\ab[8][6] ) );
  NOR2X0 U3453 ( .IN1(n2162), .IN2(n2073), .QN(\ab[8][5] ) );
  NOR2X0 U3454 ( .IN1(n2166), .IN2(n2073), .QN(\ab[8][4] ) );
  NOR2X0 U3455 ( .IN1(n2168), .IN2(n2073), .QN(\ab[8][3] ) );
  NOR2X0 U3456 ( .IN1(A[8]), .IN2(n2094), .QN(\ab[8][31] ) );
  NOR2X0 U3457 ( .IN1(n2095), .IN2(n2072), .QN(\ab[8][30] ) );
  NOR2X0 U3458 ( .IN1(n2169), .IN2(n2072), .QN(\ab[8][2] ) );
  NOR2X0 U3459 ( .IN1(n578), .IN2(n2072), .QN(\ab[8][29] ) );
  NOR2X0 U3460 ( .IN1(n2100), .IN2(n2072), .QN(\ab[8][28] ) );
  NOR2X0 U3461 ( .IN1(n2102), .IN2(n2072), .QN(\ab[8][27] ) );
  NOR2X0 U3462 ( .IN1(n2104), .IN2(n2072), .QN(\ab[8][26] ) );
  NOR2X0 U3463 ( .IN1(n2107), .IN2(n2072), .QN(\ab[8][25] ) );
  NOR2X0 U3464 ( .IN1(n2110), .IN2(n2072), .QN(\ab[8][24] ) );
  NOR2X0 U3465 ( .IN1(n2115), .IN2(n2072), .QN(\ab[8][23] ) );
  NOR2X0 U3466 ( .IN1(n2118), .IN2(n2072), .QN(\ab[8][22] ) );
  NOR2X0 U3467 ( .IN1(n2119), .IN2(n2072), .QN(\ab[8][21] ) );
  NOR2X0 U3468 ( .IN1(n2124), .IN2(n2072), .QN(\ab[8][20] ) );
  NOR2X0 U3469 ( .IN1(n2171), .IN2(n2071), .QN(\ab[8][1] ) );
  NOR2X0 U3470 ( .IN1(n2125), .IN2(n2071), .QN(\ab[8][19] ) );
  NOR2X0 U3471 ( .IN1(n2128), .IN2(n2071), .QN(\ab[8][18] ) );
  NOR2X0 U3472 ( .IN1(n2131), .IN2(n2071), .QN(\ab[8][17] ) );
  NOR2X0 U3473 ( .IN1(n2137), .IN2(n2071), .QN(\ab[8][15] ) );
  NOR2X0 U3474 ( .IN1(n2142), .IN2(n2071), .QN(\ab[8][14] ) );
  NOR2X0 U3475 ( .IN1(n2143), .IN2(n2071), .QN(\ab[8][13] ) );
  NOR2X0 U3476 ( .IN1(n1903), .IN2(n2071), .QN(\ab[8][12] ) );
  NOR2X0 U3477 ( .IN1(n2148), .IN2(n2071), .QN(\ab[8][11] ) );
  NOR2X0 U3478 ( .IN1(n2149), .IN2(n2071), .QN(\ab[8][10] ) );
  NOR2X0 U3479 ( .IN1(n2172), .IN2(n2071), .QN(\ab[8][0] ) );
  NOR2X0 U3480 ( .IN1(n2152), .IN2(n2076), .QN(\ab[7][9] ) );
  NOR2X0 U3481 ( .IN1(n2155), .IN2(n2076), .QN(\ab[7][8] ) );
  NOR2X0 U3482 ( .IN1(n2159), .IN2(n2076), .QN(\ab[7][7] ) );
  NOR2X0 U3483 ( .IN1(n2161), .IN2(n2076), .QN(\ab[7][6] ) );
  NOR2X0 U3484 ( .IN1(n2162), .IN2(n2076), .QN(\ab[7][5] ) );
  NOR2X0 U3485 ( .IN1(n2164), .IN2(n2076), .QN(\ab[7][4] ) );
  NOR2X0 U3486 ( .IN1(n2168), .IN2(n2076), .QN(\ab[7][3] ) );
  NOR2X0 U3487 ( .IN1(A[7]), .IN2(n2094), .QN(\ab[7][31] ) );
  NOR2X0 U3488 ( .IN1(n2096), .IN2(n2075), .QN(\ab[7][30] ) );
  NOR2X0 U3489 ( .IN1(n1945), .IN2(n2075), .QN(\ab[7][2] ) );
  NOR2X0 U3490 ( .IN1(n579), .IN2(n2075), .QN(\ab[7][29] ) );
  NOR2X0 U3491 ( .IN1(n2098), .IN2(n2075), .QN(\ab[7][28] ) );
  NOR2X0 U3492 ( .IN1(n2101), .IN2(n2075), .QN(\ab[7][27] ) );
  NOR2X0 U3493 ( .IN1(n2106), .IN2(n2075), .QN(\ab[7][26] ) );
  NOR2X0 U3494 ( .IN1(n2107), .IN2(n2075), .QN(\ab[7][25] ) );
  NOR2X0 U3495 ( .IN1(n2110), .IN2(n2075), .QN(\ab[7][24] ) );
  NOR2X0 U3496 ( .IN1(n2113), .IN2(n2075), .QN(\ab[7][23] ) );
  NOR2X0 U3497 ( .IN1(n2116), .IN2(n2075), .QN(\ab[7][22] ) );
  NOR2X0 U3498 ( .IN1(n2119), .IN2(n2075), .QN(\ab[7][21] ) );
  NOR2X0 U3499 ( .IN1(n2122), .IN2(n2075), .QN(\ab[7][20] ) );
  NOR2X0 U3500 ( .IN1(n2170), .IN2(n2074), .QN(\ab[7][1] ) );
  NOR2X0 U3501 ( .IN1(n2125), .IN2(n2074), .QN(\ab[7][19] ) );
  NOR2X0 U3502 ( .IN1(n2128), .IN2(n2074), .QN(\ab[7][18] ) );
  NOR2X0 U3503 ( .IN1(n2131), .IN2(n2074), .QN(\ab[7][17] ) );
  NOR2X0 U3504 ( .IN1(n2134), .IN2(n2074), .QN(\ab[7][16] ) );
  NOR2X0 U3505 ( .IN1(n2137), .IN2(n2074), .QN(\ab[7][15] ) );
  NOR2X0 U3506 ( .IN1(n2140), .IN2(n2074), .QN(\ab[7][14] ) );
  NOR2X0 U3507 ( .IN1(n2143), .IN2(n2074), .QN(\ab[7][13] ) );
  NOR2X0 U3508 ( .IN1(n1904), .IN2(n2074), .QN(\ab[7][12] ) );
  NOR2X0 U3509 ( .IN1(n2148), .IN2(n2074), .QN(\ab[7][11] ) );
  NOR2X0 U3510 ( .IN1(n2149), .IN2(n2074), .QN(\ab[7][10] ) );
  NOR2X0 U3511 ( .IN1(n2172), .IN2(n2074), .QN(\ab[7][0] ) );
  NOR2X0 U3512 ( .IN1(n2153), .IN2(n2079), .QN(\ab[6][9] ) );
  NOR2X0 U3513 ( .IN1(n2157), .IN2(n2079), .QN(\ab[6][8] ) );
  NOR2X0 U3514 ( .IN1(n2158), .IN2(n2079), .QN(\ab[6][7] ) );
  NOR2X0 U3515 ( .IN1(n2160), .IN2(n2079), .QN(\ab[6][6] ) );
  NOR2X0 U3516 ( .IN1(n2162), .IN2(n2079), .QN(\ab[6][5] ) );
  NOR2X0 U3517 ( .IN1(n2166), .IN2(n2079), .QN(\ab[6][4] ) );
  NOR2X0 U3518 ( .IN1(n2168), .IN2(n2079), .QN(\ab[6][3] ) );
  NOR2X0 U3519 ( .IN1(A[6]), .IN2(n2208), .QN(\ab[6][31] ) );
  NOR2X0 U3520 ( .IN1(n2095), .IN2(n2078), .QN(\ab[6][30] ) );
  NOR2X0 U3521 ( .IN1(n1946), .IN2(n2078), .QN(\ab[6][2] ) );
  NOR2X0 U3522 ( .IN1(n2097), .IN2(n2078), .QN(\ab[6][29] ) );
  NOR2X0 U3523 ( .IN1(n2099), .IN2(n2078), .QN(\ab[6][28] ) );
  NOR2X0 U3524 ( .IN1(n2102), .IN2(n2078), .QN(\ab[6][27] ) );
  NOR2X0 U3525 ( .IN1(n2104), .IN2(n2078), .QN(\ab[6][26] ) );
  NOR2X0 U3526 ( .IN1(n2107), .IN2(n2078), .QN(\ab[6][25] ) );
  NOR2X0 U3527 ( .IN1(n2110), .IN2(n2078), .QN(\ab[6][24] ) );
  NOR2X0 U3528 ( .IN1(n2114), .IN2(n2078), .QN(\ab[6][23] ) );
  NOR2X0 U3529 ( .IN1(n2117), .IN2(n2078), .QN(\ab[6][22] ) );
  NOR2X0 U3530 ( .IN1(n2119), .IN2(n2078), .QN(\ab[6][21] ) );
  NOR2X0 U3531 ( .IN1(n2123), .IN2(n2078), .QN(\ab[6][20] ) );
  NOR2X0 U3532 ( .IN1(n2171), .IN2(n2077), .QN(\ab[6][1] ) );
  NOR2X0 U3533 ( .IN1(n2125), .IN2(n2077), .QN(\ab[6][19] ) );
  NOR2X0 U3534 ( .IN1(n2128), .IN2(n2077), .QN(\ab[6][18] ) );
  NOR2X0 U3535 ( .IN1(n2131), .IN2(n2077), .QN(\ab[6][17] ) );
  NOR2X0 U3536 ( .IN1(n2134), .IN2(n2077), .QN(\ab[6][16] ) );
  NOR2X0 U3537 ( .IN1(n2137), .IN2(n2077), .QN(\ab[6][15] ) );
  NOR2X0 U3538 ( .IN1(n2142), .IN2(n2077), .QN(\ab[6][14] ) );
  NOR2X0 U3539 ( .IN1(n2143), .IN2(n2077), .QN(\ab[6][13] ) );
  NOR2X0 U3540 ( .IN1(n1903), .IN2(n2077), .QN(\ab[6][12] ) );
  NOR2X0 U3541 ( .IN1(n2148), .IN2(n2077), .QN(\ab[6][11] ) );
  NOR2X0 U3542 ( .IN1(n2149), .IN2(n2077), .QN(\ab[6][10] ) );
  NOR2X0 U3543 ( .IN1(n2172), .IN2(n2077), .QN(\ab[6][0] ) );
  NOR2X0 U3544 ( .IN1(n2152), .IN2(n2082), .QN(\ab[5][9] ) );
  NOR2X0 U3545 ( .IN1(n2155), .IN2(n2082), .QN(\ab[5][8] ) );
  NOR2X0 U3546 ( .IN1(n2158), .IN2(n2082), .QN(\ab[5][7] ) );
  NOR2X0 U3547 ( .IN1(n2160), .IN2(n2082), .QN(\ab[5][6] ) );
  NOR2X0 U3548 ( .IN1(n2162), .IN2(n2082), .QN(\ab[5][5] ) );
  NOR2X0 U3549 ( .IN1(n2164), .IN2(n2082), .QN(\ab[5][4] ) );
  NOR2X0 U3550 ( .IN1(n2168), .IN2(n2082), .QN(\ab[5][3] ) );
  NOR2X0 U3551 ( .IN1(A[5]), .IN2(n2208), .QN(\ab[5][31] ) );
  NOR2X0 U3552 ( .IN1(n2096), .IN2(n2081), .QN(\ab[5][30] ) );
  NOR2X0 U3553 ( .IN1(n2169), .IN2(n2081), .QN(\ab[5][2] ) );
  NOR2X0 U3554 ( .IN1(n578), .IN2(n2081), .QN(\ab[5][29] ) );
  NOR2X0 U3555 ( .IN1(n2100), .IN2(n2081), .QN(\ab[5][28] ) );
  NOR2X0 U3556 ( .IN1(n2101), .IN2(n2081), .QN(\ab[5][27] ) );
  NOR2X0 U3557 ( .IN1(n2106), .IN2(n2081), .QN(\ab[5][26] ) );
  NOR2X0 U3558 ( .IN1(n2107), .IN2(n2081), .QN(\ab[5][25] ) );
  NOR2X0 U3559 ( .IN1(n2110), .IN2(n2081), .QN(\ab[5][24] ) );
  NOR2X0 U3560 ( .IN1(n2115), .IN2(n2081), .QN(\ab[5][23] ) );
  NOR2X0 U3561 ( .IN1(n2118), .IN2(n2081), .QN(\ab[5][22] ) );
  NOR2X0 U3562 ( .IN1(n2119), .IN2(n2081), .QN(\ab[5][21] ) );
  NOR2X0 U3563 ( .IN1(n2124), .IN2(n2081), .QN(\ab[5][20] ) );
  NOR2X0 U3564 ( .IN1(n2170), .IN2(n2080), .QN(\ab[5][1] ) );
  NOR2X0 U3565 ( .IN1(n2125), .IN2(n2080), .QN(\ab[5][19] ) );
  NOR2X0 U3566 ( .IN1(n2128), .IN2(n2080), .QN(\ab[5][18] ) );
  NOR2X0 U3567 ( .IN1(n2131), .IN2(n2080), .QN(\ab[5][17] ) );
  NOR2X0 U3568 ( .IN1(n2134), .IN2(n2080), .QN(\ab[5][16] ) );
  NOR2X0 U3569 ( .IN1(n2137), .IN2(n2080), .QN(\ab[5][15] ) );
  NOR2X0 U3570 ( .IN1(n2140), .IN2(n2080), .QN(\ab[5][14] ) );
  NOR2X0 U3571 ( .IN1(n2143), .IN2(n2080), .QN(\ab[5][13] ) );
  NOR2X0 U3572 ( .IN1(n1904), .IN2(n2080), .QN(\ab[5][12] ) );
  NOR2X0 U3573 ( .IN1(n2148), .IN2(n2080), .QN(\ab[5][11] ) );
  NOR2X0 U3574 ( .IN1(n2149), .IN2(n2080), .QN(\ab[5][10] ) );
  NOR2X0 U3575 ( .IN1(n2172), .IN2(n2080), .QN(\ab[5][0] ) );
  NOR2X0 U3576 ( .IN1(n2152), .IN2(n2085), .QN(\ab[4][9] ) );
  NOR2X0 U3577 ( .IN1(n2157), .IN2(n2085), .QN(\ab[4][8] ) );
  NOR2X0 U3578 ( .IN1(n2159), .IN2(n2085), .QN(\ab[4][7] ) );
  NOR2X0 U3579 ( .IN1(n2161), .IN2(n2085), .QN(\ab[4][6] ) );
  NOR2X0 U3580 ( .IN1(n2162), .IN2(n2085), .QN(\ab[4][5] ) );
  NOR2X0 U3581 ( .IN1(n2166), .IN2(n2085), .QN(\ab[4][4] ) );
  NOR2X0 U3582 ( .IN1(n2168), .IN2(n2085), .QN(\ab[4][3] ) );
  NOR2X0 U3583 ( .IN1(A[4]), .IN2(n2208), .QN(\ab[4][31] ) );
  NOR2X0 U3584 ( .IN1(n2095), .IN2(n2084), .QN(\ab[4][30] ) );
  NOR2X0 U3585 ( .IN1(n1945), .IN2(n2084), .QN(\ab[4][2] ) );
  NOR2X0 U3586 ( .IN1(n579), .IN2(n2084), .QN(\ab[4][29] ) );
  NOR2X0 U3587 ( .IN1(n2098), .IN2(n2084), .QN(\ab[4][28] ) );
  NOR2X0 U3588 ( .IN1(n2102), .IN2(n2084), .QN(\ab[4][27] ) );
  NOR2X0 U3589 ( .IN1(n2104), .IN2(n2084), .QN(\ab[4][26] ) );
  NOR2X0 U3590 ( .IN1(n2107), .IN2(n2084), .QN(\ab[4][25] ) );
  NOR2X0 U3591 ( .IN1(n2110), .IN2(n2084), .QN(\ab[4][24] ) );
  NOR2X0 U3592 ( .IN1(n2113), .IN2(n2084), .QN(\ab[4][23] ) );
  NOR2X0 U3593 ( .IN1(n2116), .IN2(n2084), .QN(\ab[4][22] ) );
  NOR2X0 U3594 ( .IN1(n2119), .IN2(n2084), .QN(\ab[4][21] ) );
  NOR2X0 U3595 ( .IN1(n2122), .IN2(n2084), .QN(\ab[4][20] ) );
  NOR2X0 U3596 ( .IN1(n2171), .IN2(n2083), .QN(\ab[4][1] ) );
  NOR2X0 U3597 ( .IN1(n2125), .IN2(n2083), .QN(\ab[4][19] ) );
  NOR2X0 U3598 ( .IN1(n2128), .IN2(n2083), .QN(\ab[4][18] ) );
  NOR2X0 U3599 ( .IN1(n2131), .IN2(n2083), .QN(\ab[4][17] ) );
  NOR2X0 U3600 ( .IN1(n2134), .IN2(n2083), .QN(\ab[4][16] ) );
  NOR2X0 U3601 ( .IN1(n2137), .IN2(n2083), .QN(\ab[4][15] ) );
  NOR2X0 U3602 ( .IN1(n2142), .IN2(n2083), .QN(\ab[4][14] ) );
  NOR2X0 U3603 ( .IN1(n2143), .IN2(n2083), .QN(\ab[4][13] ) );
  NOR2X0 U3604 ( .IN1(n2146), .IN2(n2083), .QN(\ab[4][12] ) );
  NOR2X0 U3605 ( .IN1(n2148), .IN2(n2083), .QN(\ab[4][11] ) );
  NOR2X0 U3606 ( .IN1(n2149), .IN2(n2083), .QN(\ab[4][10] ) );
  NOR2X0 U3607 ( .IN1(n2172), .IN2(n2083), .QN(\ab[4][0] ) );
  NOR2X0 U3608 ( .IN1(n2153), .IN2(n2088), .QN(\ab[3][9] ) );
  NOR2X0 U3609 ( .IN1(n2155), .IN2(n2088), .QN(\ab[3][8] ) );
  NOR2X0 U3610 ( .IN1(n2158), .IN2(n2088), .QN(\ab[3][7] ) );
  NOR2X0 U3611 ( .IN1(n2160), .IN2(n2088), .QN(\ab[3][6] ) );
  NOR2X0 U3612 ( .IN1(n2162), .IN2(n2088), .QN(\ab[3][5] ) );
  NOR2X0 U3613 ( .IN1(n2164), .IN2(n2088), .QN(\ab[3][4] ) );
  NOR2X0 U3614 ( .IN1(n2168), .IN2(n2088), .QN(\ab[3][3] ) );
  NOR2X0 U3615 ( .IN1(A[3]), .IN2(n2208), .QN(\ab[3][31] ) );
  NOR2X0 U3616 ( .IN1(n2096), .IN2(n2087), .QN(\ab[3][30] ) );
  NOR2X0 U3617 ( .IN1(n1946), .IN2(n2087), .QN(\ab[3][2] ) );
  NOR2X0 U3618 ( .IN1(n580), .IN2(n2087), .QN(\ab[3][29] ) );
  NOR2X0 U3619 ( .IN1(n2099), .IN2(n2087), .QN(\ab[3][28] ) );
  NOR2X0 U3620 ( .IN1(n2101), .IN2(n2087), .QN(\ab[3][27] ) );
  NOR2X0 U3621 ( .IN1(n2106), .IN2(n2087), .QN(\ab[3][26] ) );
  NOR2X0 U3622 ( .IN1(n2107), .IN2(n2087), .QN(\ab[3][25] ) );
  NOR2X0 U3623 ( .IN1(n2110), .IN2(n2087), .QN(\ab[3][24] ) );
  NOR2X0 U3624 ( .IN1(n2114), .IN2(n2087), .QN(\ab[3][23] ) );
  NOR2X0 U3625 ( .IN1(n2117), .IN2(n2087), .QN(\ab[3][22] ) );
  NOR2X0 U3626 ( .IN1(n2119), .IN2(n2087), .QN(\ab[3][21] ) );
  NOR2X0 U3627 ( .IN1(n2123), .IN2(n2087), .QN(\ab[3][20] ) );
  NOR2X0 U3628 ( .IN1(n2170), .IN2(n2086), .QN(\ab[3][1] ) );
  NOR2X0 U3629 ( .IN1(n2125), .IN2(n2086), .QN(\ab[3][19] ) );
  NOR2X0 U3630 ( .IN1(n2128), .IN2(n2086), .QN(\ab[3][18] ) );
  NOR2X0 U3631 ( .IN1(n2131), .IN2(n2086), .QN(\ab[3][17] ) );
  NOR2X0 U3632 ( .IN1(n2134), .IN2(n2086), .QN(\ab[3][16] ) );
  NOR2X0 U3633 ( .IN1(n2137), .IN2(n2086), .QN(\ab[3][15] ) );
  NOR2X0 U3634 ( .IN1(n2140), .IN2(n2086), .QN(\ab[3][14] ) );
  NOR2X0 U3635 ( .IN1(n2143), .IN2(n2086), .QN(\ab[3][13] ) );
  NOR2X0 U3636 ( .IN1(n1903), .IN2(n2086), .QN(\ab[3][12] ) );
  NOR2X0 U3637 ( .IN1(n2147), .IN2(n2086), .QN(\ab[3][11] ) );
  NOR2X0 U3638 ( .IN1(n2149), .IN2(n2086), .QN(\ab[3][10] ) );
  NOR2X0 U3639 ( .IN1(n2172), .IN2(n2086), .QN(\ab[3][0] ) );
  NOR2X0 U3640 ( .IN1(B[9]), .IN2(n2004), .QN(\ab[31][9] ) );
  NOR2X0 U3641 ( .IN1(B[8]), .IN2(n2004), .QN(\ab[31][8] ) );
  NOR2X0 U3642 ( .IN1(B[6]), .IN2(n2004), .QN(\ab[31][6] ) );
  NOR2X0 U3643 ( .IN1(B[5]), .IN2(n2004), .QN(\ab[31][5] ) );
  NOR2X0 U3644 ( .IN1(B[4]), .IN2(n2004), .QN(\ab[31][4] ) );
  NOR2X0 U3645 ( .IN1(B[3]), .IN2(n2004), .QN(\ab[31][3] ) );
  NOR2X0 U3646 ( .IN1(n2094), .IN2(n2004), .QN(\ab[31][31] ) );
  NOR2X0 U3647 ( .IN1(n546), .IN2(n2004), .QN(\ab[31][30] ) );
  NOR2X0 U3648 ( .IN1(B[2]), .IN2(n2004), .QN(\ab[31][2] ) );
  NOR2X0 U3649 ( .IN1(B[29]), .IN2(n2004), .QN(\ab[31][29] ) );
  NOR2X0 U3650 ( .IN1(B[28]), .IN2(n2004), .QN(\ab[31][28] ) );
  NOR2X0 U3651 ( .IN1(B[27]), .IN2(n2004), .QN(\ab[31][27] ) );
  NOR2X0 U3652 ( .IN1(B[26]), .IN2(n2004), .QN(\ab[31][26] ) );
  NOR2X0 U3653 ( .IN1(B[25]), .IN2(n2004), .QN(\ab[31][25] ) );
  NOR2X0 U3654 ( .IN1(B[24]), .IN2(n2004), .QN(\ab[31][24] ) );
  NOR2X0 U3655 ( .IN1(B[23]), .IN2(n2004), .QN(\ab[31][23] ) );
  NOR2X0 U3656 ( .IN1(B[22]), .IN2(n2004), .QN(\ab[31][22] ) );
  NOR2X0 U3657 ( .IN1(B[21]), .IN2(n2004), .QN(\ab[31][21] ) );
  NOR2X0 U3658 ( .IN1(B[20]), .IN2(n2004), .QN(\ab[31][20] ) );
  NOR2X0 U3659 ( .IN1(B[1]), .IN2(n2004), .QN(\ab[31][1] ) );
  NOR2X0 U3660 ( .IN1(B[19]), .IN2(n2004), .QN(\ab[31][19] ) );
  NOR2X0 U3661 ( .IN1(B[18]), .IN2(n2004), .QN(\ab[31][18] ) );
  NOR2X0 U3662 ( .IN1(B[17]), .IN2(n2004), .QN(\ab[31][17] ) );
  NOR2X0 U3663 ( .IN1(n20), .IN2(n2004), .QN(\ab[31][16] ) );
  NOR2X0 U3664 ( .IN1(B[15]), .IN2(n2004), .QN(\ab[31][15] ) );
  NOR2X0 U3665 ( .IN1(B[14]), .IN2(n2004), .QN(\ab[31][14] ) );
  NOR2X0 U3666 ( .IN1(n28), .IN2(n2004), .QN(\ab[31][13] ) );
  NOR2X0 U3667 ( .IN1(B[12]), .IN2(n2004), .QN(\ab[31][12] ) );
  NOR2X0 U3668 ( .IN1(B[11]), .IN2(n2004), .QN(\ab[31][11] ) );
  NOR2X0 U3669 ( .IN1(B[0]), .IN2(n2004), .QN(\ab[31][0] ) );
  NOR2X0 U3670 ( .IN1(n2153), .IN2(n2007), .QN(\ab[30][9] ) );
  NOR2X0 U3671 ( .IN1(n2157), .IN2(n2007), .QN(\ab[30][8] ) );
  NOR2X0 U3672 ( .IN1(n2158), .IN2(n2007), .QN(\ab[30][7] ) );
  NOR2X0 U3673 ( .IN1(n2160), .IN2(n2007), .QN(\ab[30][6] ) );
  NOR2X0 U3674 ( .IN1(n2162), .IN2(n2007), .QN(\ab[30][5] ) );
  NOR2X0 U3675 ( .IN1(n2166), .IN2(n2007), .QN(\ab[30][4] ) );
  NOR2X0 U3676 ( .IN1(n2168), .IN2(n2007), .QN(\ab[30][3] ) );
  NOR2X0 U3677 ( .IN1(A[30]), .IN2(n2094), .QN(\ab[30][31] ) );
  NOR2X0 U3678 ( .IN1(n2095), .IN2(n2006), .QN(\ab[30][30] ) );
  NOR2X0 U3679 ( .IN1(n1945), .IN2(n2006), .QN(\ab[30][2] ) );
  NOR2X0 U3680 ( .IN1(n2097), .IN2(n2006), .QN(\ab[30][29] ) );
  NOR2X0 U3681 ( .IN1(n2099), .IN2(n2006), .QN(\ab[30][28] ) );
  NOR2X0 U3682 ( .IN1(n2102), .IN2(n2006), .QN(\ab[30][27] ) );
  NOR2X0 U3683 ( .IN1(n2104), .IN2(n2006), .QN(\ab[30][26] ) );
  NOR2X0 U3684 ( .IN1(n2107), .IN2(n2006), .QN(\ab[30][25] ) );
  NOR2X0 U3685 ( .IN1(n2110), .IN2(n2006), .QN(\ab[30][24] ) );
  NOR2X0 U3686 ( .IN1(n2114), .IN2(n2006), .QN(\ab[30][23] ) );
  NOR2X0 U3687 ( .IN1(n2117), .IN2(n2006), .QN(\ab[30][22] ) );
  NOR2X0 U3688 ( .IN1(n2119), .IN2(n2006), .QN(\ab[30][21] ) );
  NOR2X0 U3689 ( .IN1(n2123), .IN2(n2006), .QN(\ab[30][20] ) );
  NOR2X0 U3690 ( .IN1(n2171), .IN2(n2005), .QN(\ab[30][1] ) );
  NOR2X0 U3691 ( .IN1(n2125), .IN2(n2005), .QN(\ab[30][19] ) );
  NOR2X0 U3692 ( .IN1(n2128), .IN2(n2005), .QN(\ab[30][18] ) );
  NOR2X0 U3693 ( .IN1(n2131), .IN2(n2005), .QN(\ab[30][17] ) );
  NOR2X0 U3694 ( .IN1(n2134), .IN2(n2005), .QN(\ab[30][16] ) );
  NOR2X0 U3695 ( .IN1(n2137), .IN2(n2005), .QN(\ab[30][15] ) );
  NOR2X0 U3696 ( .IN1(n2142), .IN2(n2005), .QN(\ab[30][14] ) );
  NOR2X0 U3697 ( .IN1(n2143), .IN2(n2005), .QN(\ab[30][13] ) );
  NOR2X0 U3698 ( .IN1(n2146), .IN2(n2005), .QN(\ab[30][12] ) );
  NOR2X0 U3699 ( .IN1(n2148), .IN2(n2005), .QN(\ab[30][11] ) );
  NOR2X0 U3700 ( .IN1(n2149), .IN2(n2005), .QN(\ab[30][10] ) );
  NOR2X0 U3701 ( .IN1(n2172), .IN2(n2005), .QN(\ab[30][0] ) );
  NOR2X0 U3702 ( .IN1(n2152), .IN2(n2089), .QN(\ab[2][9] ) );
  NOR2X0 U3703 ( .IN1(n2157), .IN2(n601), .QN(\ab[2][8] ) );
  NOR2X0 U3704 ( .IN1(n2158), .IN2(n600), .QN(\ab[2][7] ) );
  NOR2X0 U3705 ( .IN1(n2160), .IN2(n600), .QN(\ab[2][6] ) );
  NOR2X0 U3706 ( .IN1(n2162), .IN2(n2089), .QN(\ab[2][5] ) );
  NOR2X0 U3707 ( .IN1(n2166), .IN2(n601), .QN(\ab[2][4] ) );
  NOR2X0 U3708 ( .IN1(n2167), .IN2(n600), .QN(\ab[2][3] ) );
  NOR2X0 U3709 ( .IN1(A[2]), .IN2(n2208), .QN(\ab[2][31] ) );
  NOR2X0 U3710 ( .IN1(n2209), .IN2(n2205), .QN(\ab[2][30] ) );
  NOR2X0 U3711 ( .IN1(n2169), .IN2(n601), .QN(\ab[2][2] ) );
  NOR2X0 U3712 ( .IN1(n2210), .IN2(n2205), .QN(\ab[2][29] ) );
  NOR2X0 U3713 ( .IN1(n2098), .IN2(n2089), .QN(\ab[2][28] ) );
  NOR2X0 U3714 ( .IN1(n2102), .IN2(n2089), .QN(\ab[2][27] ) );
  NOR2X0 U3715 ( .IN1(n2105), .IN2(n601), .QN(\ab[2][26] ) );
  NOR2X0 U3716 ( .IN1(n2107), .IN2(n2089), .QN(\ab[2][25] ) );
  NOR2X0 U3717 ( .IN1(n2110), .IN2(n601), .QN(\ab[2][24] ) );
  NOR2X0 U3718 ( .IN1(n2115), .IN2(n2089), .QN(\ab[2][23] ) );
  NOR2X0 U3719 ( .IN1(n2116), .IN2(n600), .QN(\ab[2][22] ) );
  NOR2X0 U3720 ( .IN1(n2119), .IN2(n601), .QN(\ab[2][21] ) );
  NOR2X0 U3721 ( .IN1(n2122), .IN2(n600), .QN(\ab[2][20] ) );
  NOR2X0 U3722 ( .IN1(n2170), .IN2(n600), .QN(\ab[2][1] ) );
  NOR2X0 U3723 ( .IN1(n2125), .IN2(n601), .QN(\ab[2][19] ) );
  NOR2X0 U3724 ( .IN1(n2128), .IN2(n601), .QN(\ab[2][18] ) );
  NOR2X0 U3725 ( .IN1(n2131), .IN2(n2089), .QN(\ab[2][17] ) );
  NOR2X0 U3726 ( .IN1(n2134), .IN2(n600), .QN(\ab[2][16] ) );
  NOR2X0 U3727 ( .IN1(n2137), .IN2(n2089), .QN(\ab[2][15] ) );
  NOR2X0 U3728 ( .IN1(n2142), .IN2(n600), .QN(\ab[2][14] ) );
  NOR2X0 U3729 ( .IN1(n2143), .IN2(n601), .QN(\ab[2][13] ) );
  NOR2X0 U3730 ( .IN1(n2146), .IN2(n600), .QN(\ab[2][12] ) );
  NOR2X0 U3731 ( .IN1(n2147), .IN2(n601), .QN(\ab[2][11] ) );
  NOR2X0 U3732 ( .IN1(n2149), .IN2(n2089), .QN(\ab[2][10] ) );
  NOR2X0 U3733 ( .IN1(n2172), .IN2(n2089), .QN(\ab[2][0] ) );
  NOR2X0 U3734 ( .IN1(n2153), .IN2(n2010), .QN(\ab[29][9] ) );
  NOR2X0 U3735 ( .IN1(n2155), .IN2(n2010), .QN(\ab[29][8] ) );
  NOR2X0 U3736 ( .IN1(n2158), .IN2(n2010), .QN(\ab[29][7] ) );
  NOR2X0 U3737 ( .IN1(n2160), .IN2(n2010), .QN(\ab[29][6] ) );
  NOR2X0 U3738 ( .IN1(n2162), .IN2(n2010), .QN(\ab[29][5] ) );
  NOR2X0 U3739 ( .IN1(n2164), .IN2(n2010), .QN(\ab[29][4] ) );
  NOR2X0 U3740 ( .IN1(n2168), .IN2(n2010), .QN(\ab[29][3] ) );
  NOR2X0 U3741 ( .IN1(A[29]), .IN2(n2094), .QN(\ab[29][31] ) );
  NOR2X0 U3742 ( .IN1(n2096), .IN2(n2009), .QN(\ab[29][30] ) );
  NOR2X0 U3743 ( .IN1(n1946), .IN2(n2009), .QN(\ab[29][2] ) );
  NOR2X0 U3744 ( .IN1(n580), .IN2(n2009), .QN(\ab[29][29] ) );
  NOR2X0 U3745 ( .IN1(n2100), .IN2(n2009), .QN(\ab[29][28] ) );
  NOR2X0 U3746 ( .IN1(n2101), .IN2(n2009), .QN(\ab[29][27] ) );
  NOR2X0 U3747 ( .IN1(n2106), .IN2(n2009), .QN(\ab[29][26] ) );
  NOR2X0 U3748 ( .IN1(n2107), .IN2(n2009), .QN(\ab[29][25] ) );
  NOR2X0 U3749 ( .IN1(n2110), .IN2(n2009), .QN(\ab[29][24] ) );
  NOR2X0 U3750 ( .IN1(n2115), .IN2(n2009), .QN(\ab[29][23] ) );
  NOR2X0 U3751 ( .IN1(n2118), .IN2(n2009), .QN(\ab[29][22] ) );
  NOR2X0 U3752 ( .IN1(n2119), .IN2(n2009), .QN(\ab[29][21] ) );
  NOR2X0 U3753 ( .IN1(n2124), .IN2(n2009), .QN(\ab[29][20] ) );
  NOR2X0 U3754 ( .IN1(n2170), .IN2(n2008), .QN(\ab[29][1] ) );
  NOR2X0 U3755 ( .IN1(n2125), .IN2(n2008), .QN(\ab[29][19] ) );
  NOR2X0 U3756 ( .IN1(n2128), .IN2(n2008), .QN(\ab[29][18] ) );
  NOR2X0 U3757 ( .IN1(n2131), .IN2(n2008), .QN(\ab[29][17] ) );
  NOR2X0 U3758 ( .IN1(n2134), .IN2(n2008), .QN(\ab[29][16] ) );
  NOR2X0 U3759 ( .IN1(n2137), .IN2(n2008), .QN(\ab[29][15] ) );
  NOR2X0 U3760 ( .IN1(n2140), .IN2(n2008), .QN(\ab[29][14] ) );
  NOR2X0 U3761 ( .IN1(n2143), .IN2(n2008), .QN(\ab[29][13] ) );
  NOR2X0 U3762 ( .IN1(n1903), .IN2(n2008), .QN(\ab[29][12] ) );
  NOR2X0 U3763 ( .IN1(n2148), .IN2(n2008), .QN(\ab[29][11] ) );
  NOR2X0 U3764 ( .IN1(n2149), .IN2(n2008), .QN(\ab[29][10] ) );
  NOR2X0 U3765 ( .IN1(n2172), .IN2(n2008), .QN(\ab[29][0] ) );
  NOR2X0 U3766 ( .IN1(n2153), .IN2(n2013), .QN(\ab[28][9] ) );
  NOR2X0 U3767 ( .IN1(n2157), .IN2(n2013), .QN(\ab[28][8] ) );
  NOR2X0 U3768 ( .IN1(n2159), .IN2(n2013), .QN(\ab[28][7] ) );
  NOR2X0 U3769 ( .IN1(n2161), .IN2(n2013), .QN(\ab[28][6] ) );
  NOR2X0 U3770 ( .IN1(n2162), .IN2(n2013), .QN(\ab[28][5] ) );
  NOR2X0 U3771 ( .IN1(n2166), .IN2(n2013), .QN(\ab[28][4] ) );
  NOR2X0 U3772 ( .IN1(n2168), .IN2(n2013), .QN(\ab[28][3] ) );
  NOR2X0 U3773 ( .IN1(A[28]), .IN2(n2094), .QN(\ab[28][31] ) );
  NOR2X0 U3774 ( .IN1(n2095), .IN2(n2012), .QN(\ab[28][30] ) );
  NOR2X0 U3775 ( .IN1(n1945), .IN2(n2012), .QN(\ab[28][2] ) );
  NOR2X0 U3776 ( .IN1(n578), .IN2(n2012), .QN(\ab[28][29] ) );
  NOR2X0 U3777 ( .IN1(n2098), .IN2(n2012), .QN(\ab[28][28] ) );
  NOR2X0 U3778 ( .IN1(n2102), .IN2(n2012), .QN(\ab[28][27] ) );
  NOR2X0 U3779 ( .IN1(n2104), .IN2(n2012), .QN(\ab[28][26] ) );
  NOR2X0 U3780 ( .IN1(n2107), .IN2(n2012), .QN(\ab[28][25] ) );
  NOR2X0 U3781 ( .IN1(n2110), .IN2(n2012), .QN(\ab[28][24] ) );
  NOR2X0 U3782 ( .IN1(n2113), .IN2(n2012), .QN(\ab[28][23] ) );
  NOR2X0 U3783 ( .IN1(n2116), .IN2(n2012), .QN(\ab[28][22] ) );
  NOR2X0 U3784 ( .IN1(n2119), .IN2(n2012), .QN(\ab[28][21] ) );
  NOR2X0 U3785 ( .IN1(n2122), .IN2(n2012), .QN(\ab[28][20] ) );
  NOR2X0 U3786 ( .IN1(n2171), .IN2(n2011), .QN(\ab[28][1] ) );
  NOR2X0 U3787 ( .IN1(n2125), .IN2(n2011), .QN(\ab[28][19] ) );
  NOR2X0 U3788 ( .IN1(n2128), .IN2(n2011), .QN(\ab[28][18] ) );
  NOR2X0 U3789 ( .IN1(n2131), .IN2(n2011), .QN(\ab[28][17] ) );
  NOR2X0 U3790 ( .IN1(n2134), .IN2(n2011), .QN(\ab[28][16] ) );
  NOR2X0 U3791 ( .IN1(n2137), .IN2(n2011), .QN(\ab[28][15] ) );
  NOR2X0 U3792 ( .IN1(n2142), .IN2(n2011), .QN(\ab[28][14] ) );
  NOR2X0 U3793 ( .IN1(n2143), .IN2(n2011), .QN(\ab[28][13] ) );
  NOR2X0 U3794 ( .IN1(n1904), .IN2(n2011), .QN(\ab[28][12] ) );
  NOR2X0 U3795 ( .IN1(n2148), .IN2(n2011), .QN(\ab[28][11] ) );
  NOR2X0 U3796 ( .IN1(n2149), .IN2(n2011), .QN(\ab[28][10] ) );
  NOR2X0 U3797 ( .IN1(n2172), .IN2(n2011), .QN(\ab[28][0] ) );
  NOR2X0 U3798 ( .IN1(n2153), .IN2(n2016), .QN(\ab[27][9] ) );
  NOR2X0 U3799 ( .IN1(n2155), .IN2(n2016), .QN(\ab[27][8] ) );
  NOR2X0 U3800 ( .IN1(n2158), .IN2(n2016), .QN(\ab[27][7] ) );
  NOR2X0 U3801 ( .IN1(n2160), .IN2(n2016), .QN(\ab[27][6] ) );
  NOR2X0 U3802 ( .IN1(n2162), .IN2(n2016), .QN(\ab[27][5] ) );
  NOR2X0 U3803 ( .IN1(n2164), .IN2(n2016), .QN(\ab[27][4] ) );
  NOR2X0 U3804 ( .IN1(n2168), .IN2(n2016), .QN(\ab[27][3] ) );
  NOR2X0 U3805 ( .IN1(A[27]), .IN2(n2094), .QN(\ab[27][31] ) );
  NOR2X0 U3806 ( .IN1(n2096), .IN2(n2015), .QN(\ab[27][30] ) );
  NOR2X0 U3807 ( .IN1(n1946), .IN2(n2015), .QN(\ab[27][2] ) );
  NOR2X0 U3808 ( .IN1(n579), .IN2(n2015), .QN(\ab[27][29] ) );
  NOR2X0 U3809 ( .IN1(n2099), .IN2(n2015), .QN(\ab[27][28] ) );
  NOR2X0 U3810 ( .IN1(n2101), .IN2(n2015), .QN(\ab[27][27] ) );
  NOR2X0 U3811 ( .IN1(n2106), .IN2(n2015), .QN(\ab[27][26] ) );
  NOR2X0 U3812 ( .IN1(n2107), .IN2(n2015), .QN(\ab[27][25] ) );
  NOR2X0 U3813 ( .IN1(n2110), .IN2(n2015), .QN(\ab[27][24] ) );
  NOR2X0 U3814 ( .IN1(n2114), .IN2(n2015), .QN(\ab[27][23] ) );
  NOR2X0 U3815 ( .IN1(n2117), .IN2(n2015), .QN(\ab[27][22] ) );
  NOR2X0 U3816 ( .IN1(n2119), .IN2(n2015), .QN(\ab[27][21] ) );
  NOR2X0 U3817 ( .IN1(n2123), .IN2(n2015), .QN(\ab[27][20] ) );
  NOR2X0 U3818 ( .IN1(n2170), .IN2(n2014), .QN(\ab[27][1] ) );
  NOR2X0 U3819 ( .IN1(n2125), .IN2(n2014), .QN(\ab[27][19] ) );
  NOR2X0 U3820 ( .IN1(n2128), .IN2(n2014), .QN(\ab[27][18] ) );
  NOR2X0 U3821 ( .IN1(n2131), .IN2(n2014), .QN(\ab[27][17] ) );
  NOR2X0 U3822 ( .IN1(n2134), .IN2(n2014), .QN(\ab[27][16] ) );
  NOR2X0 U3823 ( .IN1(n2137), .IN2(n2014), .QN(\ab[27][15] ) );
  NOR2X0 U3824 ( .IN1(n2140), .IN2(n2014), .QN(\ab[27][14] ) );
  NOR2X0 U3825 ( .IN1(n2143), .IN2(n2014), .QN(\ab[27][13] ) );
  NOR2X0 U3826 ( .IN1(n2146), .IN2(n2014), .QN(\ab[27][12] ) );
  NOR2X0 U3827 ( .IN1(n2148), .IN2(n2014), .QN(\ab[27][11] ) );
  NOR2X0 U3828 ( .IN1(n2149), .IN2(n2014), .QN(\ab[27][10] ) );
  NOR2X0 U3829 ( .IN1(n2172), .IN2(n2014), .QN(\ab[27][0] ) );
  NOR2X0 U3830 ( .IN1(n2152), .IN2(n2019), .QN(\ab[26][9] ) );
  NOR2X0 U3831 ( .IN1(n2157), .IN2(n2019), .QN(\ab[26][8] ) );
  NOR2X0 U3832 ( .IN1(n2158), .IN2(n2019), .QN(\ab[26][7] ) );
  NOR2X0 U3833 ( .IN1(n2160), .IN2(n2019), .QN(\ab[26][6] ) );
  NOR2X0 U3834 ( .IN1(n2162), .IN2(n2019), .QN(\ab[26][5] ) );
  NOR2X0 U3835 ( .IN1(n2166), .IN2(n2019), .QN(\ab[26][4] ) );
  NOR2X0 U3836 ( .IN1(n2168), .IN2(n2019), .QN(\ab[26][3] ) );
  NOR2X0 U3837 ( .IN1(A[26]), .IN2(n2094), .QN(\ab[26][31] ) );
  NOR2X0 U3838 ( .IN1(n2095), .IN2(n2018), .QN(\ab[26][30] ) );
  NOR2X0 U3839 ( .IN1(n1945), .IN2(n2018), .QN(\ab[26][2] ) );
  NOR2X0 U3840 ( .IN1(n2097), .IN2(n2018), .QN(\ab[26][29] ) );
  NOR2X0 U3841 ( .IN1(n2100), .IN2(n2018), .QN(\ab[26][28] ) );
  NOR2X0 U3842 ( .IN1(n2102), .IN2(n2018), .QN(\ab[26][27] ) );
  NOR2X0 U3843 ( .IN1(n2104), .IN2(n2018), .QN(\ab[26][26] ) );
  NOR2X0 U3844 ( .IN1(n2107), .IN2(n2018), .QN(\ab[26][25] ) );
  NOR2X0 U3845 ( .IN1(n2110), .IN2(n2018), .QN(\ab[26][24] ) );
  NOR2X0 U3846 ( .IN1(n2115), .IN2(n2018), .QN(\ab[26][23] ) );
  NOR2X0 U3847 ( .IN1(n2118), .IN2(n2018), .QN(\ab[26][22] ) );
  NOR2X0 U3848 ( .IN1(n2119), .IN2(n2018), .QN(\ab[26][21] ) );
  NOR2X0 U3849 ( .IN1(n2124), .IN2(n2018), .QN(\ab[26][20] ) );
  NOR2X0 U3850 ( .IN1(n2171), .IN2(n2017), .QN(\ab[26][1] ) );
  NOR2X0 U3851 ( .IN1(n2125), .IN2(n2017), .QN(\ab[26][19] ) );
  NOR2X0 U3852 ( .IN1(n2128), .IN2(n2017), .QN(\ab[26][18] ) );
  NOR2X0 U3853 ( .IN1(n2131), .IN2(n2017), .QN(\ab[26][17] ) );
  NOR2X0 U3854 ( .IN1(n2134), .IN2(n2017), .QN(\ab[26][16] ) );
  NOR2X0 U3855 ( .IN1(n2137), .IN2(n2017), .QN(\ab[26][15] ) );
  NOR2X0 U3856 ( .IN1(n2142), .IN2(n2017), .QN(\ab[26][14] ) );
  NOR2X0 U3857 ( .IN1(n2143), .IN2(n2017), .QN(\ab[26][13] ) );
  NOR2X0 U3858 ( .IN1(n1903), .IN2(n2017), .QN(\ab[26][12] ) );
  NOR2X0 U3859 ( .IN1(n2148), .IN2(n2017), .QN(\ab[26][11] ) );
  NOR2X0 U3860 ( .IN1(n2149), .IN2(n2017), .QN(\ab[26][10] ) );
  NOR2X0 U3861 ( .IN1(n2172), .IN2(n2017), .QN(\ab[26][0] ) );
  NOR2X0 U3862 ( .IN1(n2153), .IN2(n2022), .QN(\ab[25][9] ) );
  NOR2X0 U3863 ( .IN1(n2155), .IN2(n2022), .QN(\ab[25][8] ) );
  NOR2X0 U3864 ( .IN1(n2159), .IN2(n2022), .QN(\ab[25][7] ) );
  NOR2X0 U3865 ( .IN1(n2161), .IN2(n2022), .QN(\ab[25][6] ) );
  NOR2X0 U3866 ( .IN1(n2162), .IN2(n2022), .QN(\ab[25][5] ) );
  NOR2X0 U3867 ( .IN1(n2164), .IN2(n2022), .QN(\ab[25][4] ) );
  NOR2X0 U3868 ( .IN1(n2168), .IN2(n2022), .QN(\ab[25][3] ) );
  NOR2X0 U3869 ( .IN1(A[25]), .IN2(n2094), .QN(\ab[25][31] ) );
  NOR2X0 U3870 ( .IN1(n2096), .IN2(n2021), .QN(\ab[25][30] ) );
  NOR2X0 U3871 ( .IN1(n1946), .IN2(n2021), .QN(\ab[25][2] ) );
  NOR2X0 U3872 ( .IN1(n580), .IN2(n2021), .QN(\ab[25][29] ) );
  NOR2X0 U3873 ( .IN1(n2098), .IN2(n2021), .QN(\ab[25][28] ) );
  NOR2X0 U3874 ( .IN1(n2101), .IN2(n2021), .QN(\ab[25][27] ) );
  NOR2X0 U3875 ( .IN1(n2106), .IN2(n2021), .QN(\ab[25][26] ) );
  NOR2X0 U3876 ( .IN1(n2108), .IN2(n2021), .QN(\ab[25][25] ) );
  NOR2X0 U3877 ( .IN1(n2111), .IN2(n2021), .QN(\ab[25][24] ) );
  NOR2X0 U3878 ( .IN1(n2113), .IN2(n2021), .QN(\ab[25][23] ) );
  NOR2X0 U3879 ( .IN1(n2116), .IN2(n2021), .QN(\ab[25][22] ) );
  NOR2X0 U3880 ( .IN1(n2120), .IN2(n2021), .QN(\ab[25][21] ) );
  NOR2X0 U3881 ( .IN1(n2122), .IN2(n2021), .QN(\ab[25][20] ) );
  NOR2X0 U3882 ( .IN1(n2170), .IN2(n2020), .QN(\ab[25][1] ) );
  NOR2X0 U3883 ( .IN1(n2126), .IN2(n2020), .QN(\ab[25][19] ) );
  NOR2X0 U3884 ( .IN1(n2129), .IN2(n2020), .QN(\ab[25][18] ) );
  NOR2X0 U3885 ( .IN1(n2132), .IN2(n2020), .QN(\ab[25][17] ) );
  NOR2X0 U3886 ( .IN1(n2135), .IN2(n2020), .QN(\ab[25][16] ) );
  NOR2X0 U3887 ( .IN1(n2138), .IN2(n2020), .QN(\ab[25][15] ) );
  NOR2X0 U3888 ( .IN1(n2140), .IN2(n2020), .QN(\ab[25][14] ) );
  NOR2X0 U3889 ( .IN1(n2144), .IN2(n2020), .QN(\ab[25][13] ) );
  NOR2X0 U3890 ( .IN1(n1904), .IN2(n2020), .QN(\ab[25][12] ) );
  NOR2X0 U3891 ( .IN1(n2148), .IN2(n2020), .QN(\ab[25][11] ) );
  NOR2X0 U3892 ( .IN1(n2150), .IN2(n2020), .QN(\ab[25][10] ) );
  NOR2X0 U3893 ( .IN1(n2173), .IN2(n2020), .QN(\ab[25][0] ) );
  NOR2X0 U3894 ( .IN1(n2152), .IN2(n2025), .QN(\ab[24][9] ) );
  NOR2X0 U3895 ( .IN1(n2157), .IN2(n2025), .QN(\ab[24][8] ) );
  NOR2X0 U3896 ( .IN1(n2158), .IN2(n2025), .QN(\ab[24][7] ) );
  NOR2X0 U3897 ( .IN1(n2160), .IN2(n2025), .QN(\ab[24][6] ) );
  NOR2X0 U3898 ( .IN1(n2162), .IN2(n2025), .QN(\ab[24][5] ) );
  NOR2X0 U3899 ( .IN1(n2166), .IN2(n2025), .QN(\ab[24][4] ) );
  NOR2X0 U3900 ( .IN1(n2168), .IN2(n2025), .QN(\ab[24][3] ) );
  NOR2X0 U3901 ( .IN1(A[24]), .IN2(n2094), .QN(\ab[24][31] ) );
  NOR2X0 U3902 ( .IN1(n2095), .IN2(n2024), .QN(\ab[24][30] ) );
  NOR2X0 U3903 ( .IN1(n1945), .IN2(n2024), .QN(\ab[24][2] ) );
  NOR2X0 U3904 ( .IN1(n578), .IN2(n2024), .QN(\ab[24][29] ) );
  NOR2X0 U3905 ( .IN1(n2099), .IN2(n2024), .QN(\ab[24][28] ) );
  NOR2X0 U3906 ( .IN1(n2102), .IN2(n2024), .QN(\ab[24][27] ) );
  NOR2X0 U3907 ( .IN1(n2104), .IN2(n2024), .QN(\ab[24][26] ) );
  NOR2X0 U3908 ( .IN1(n2108), .IN2(n2024), .QN(\ab[24][25] ) );
  NOR2X0 U3909 ( .IN1(n2111), .IN2(n2024), .QN(\ab[24][24] ) );
  NOR2X0 U3910 ( .IN1(n2114), .IN2(n2024), .QN(\ab[24][23] ) );
  NOR2X0 U3911 ( .IN1(n2116), .IN2(n2024), .QN(\ab[24][22] ) );
  NOR2X0 U3912 ( .IN1(n2120), .IN2(n2024), .QN(\ab[24][21] ) );
  NOR2X0 U3913 ( .IN1(n2123), .IN2(n2024), .QN(\ab[24][20] ) );
  NOR2X0 U3914 ( .IN1(n2171), .IN2(n2023), .QN(\ab[24][1] ) );
  NOR2X0 U3915 ( .IN1(n2126), .IN2(n2023), .QN(\ab[24][19] ) );
  NOR2X0 U3916 ( .IN1(n2129), .IN2(n2023), .QN(\ab[24][18] ) );
  NOR2X0 U3917 ( .IN1(n2132), .IN2(n2023), .QN(\ab[24][17] ) );
  NOR2X0 U3918 ( .IN1(n2135), .IN2(n2023), .QN(\ab[24][16] ) );
  NOR2X0 U3919 ( .IN1(n2138), .IN2(n2023), .QN(\ab[24][15] ) );
  NOR2X0 U3920 ( .IN1(n2142), .IN2(n2023), .QN(\ab[24][14] ) );
  NOR2X0 U3921 ( .IN1(n2144), .IN2(n2023), .QN(\ab[24][13] ) );
  NOR2X0 U3922 ( .IN1(n2146), .IN2(n2023), .QN(\ab[24][12] ) );
  NOR2X0 U3923 ( .IN1(n2148), .IN2(n2023), .QN(\ab[24][11] ) );
  NOR2X0 U3924 ( .IN1(n2150), .IN2(n2023), .QN(\ab[24][10] ) );
  NOR2X0 U3925 ( .IN1(n2173), .IN2(n2023), .QN(\ab[24][0] ) );
  NOR2X0 U3926 ( .IN1(n2153), .IN2(n2028), .QN(\ab[23][9] ) );
  NOR2X0 U3927 ( .IN1(n2155), .IN2(n2028), .QN(\ab[23][8] ) );
  NOR2X0 U3928 ( .IN1(n2158), .IN2(n2028), .QN(\ab[23][7] ) );
  NOR2X0 U3929 ( .IN1(n2160), .IN2(n2028), .QN(\ab[23][6] ) );
  NOR2X0 U3930 ( .IN1(n2162), .IN2(n2028), .QN(\ab[23][5] ) );
  NOR2X0 U3931 ( .IN1(n2164), .IN2(n2028), .QN(\ab[23][4] ) );
  NOR2X0 U3932 ( .IN1(n2168), .IN2(n2028), .QN(\ab[23][3] ) );
  NOR2X0 U3933 ( .IN1(A[23]), .IN2(n2094), .QN(\ab[23][31] ) );
  NOR2X0 U3934 ( .IN1(n2096), .IN2(n2027), .QN(\ab[23][30] ) );
  NOR2X0 U3935 ( .IN1(n1946), .IN2(n2027), .QN(\ab[23][2] ) );
  NOR2X0 U3936 ( .IN1(n579), .IN2(n2027), .QN(\ab[23][29] ) );
  NOR2X0 U3937 ( .IN1(n2100), .IN2(n2027), .QN(\ab[23][28] ) );
  NOR2X0 U3938 ( .IN1(n2101), .IN2(n2027), .QN(\ab[23][27] ) );
  NOR2X0 U3939 ( .IN1(n2106), .IN2(n2027), .QN(\ab[23][26] ) );
  NOR2X0 U3940 ( .IN1(n2108), .IN2(n2027), .QN(\ab[23][25] ) );
  NOR2X0 U3941 ( .IN1(n2111), .IN2(n2027), .QN(\ab[23][24] ) );
  NOR2X0 U3942 ( .IN1(n2115), .IN2(n2027), .QN(\ab[23][23] ) );
  NOR2X0 U3943 ( .IN1(n2117), .IN2(n2027), .QN(\ab[23][22] ) );
  NOR2X0 U3944 ( .IN1(n2120), .IN2(n2027), .QN(\ab[23][21] ) );
  NOR2X0 U3945 ( .IN1(n2124), .IN2(n2027), .QN(\ab[23][20] ) );
  NOR2X0 U3946 ( .IN1(n2170), .IN2(n2026), .QN(\ab[23][1] ) );
  NOR2X0 U3947 ( .IN1(n2126), .IN2(n2026), .QN(\ab[23][19] ) );
  NOR2X0 U3948 ( .IN1(n2129), .IN2(n2026), .QN(\ab[23][18] ) );
  NOR2X0 U3949 ( .IN1(n2132), .IN2(n2026), .QN(\ab[23][17] ) );
  NOR2X0 U3950 ( .IN1(n2135), .IN2(n2026), .QN(\ab[23][16] ) );
  NOR2X0 U3951 ( .IN1(n2138), .IN2(n2026), .QN(\ab[23][15] ) );
  NOR2X0 U3952 ( .IN1(n2140), .IN2(n2026), .QN(\ab[23][14] ) );
  NOR2X0 U3953 ( .IN1(n2144), .IN2(n2026), .QN(\ab[23][13] ) );
  NOR2X0 U3954 ( .IN1(n1903), .IN2(n2026), .QN(\ab[23][12] ) );
  NOR2X0 U3955 ( .IN1(n2148), .IN2(n2026), .QN(\ab[23][11] ) );
  NOR2X0 U3956 ( .IN1(n2150), .IN2(n2026), .QN(\ab[23][10] ) );
  NOR2X0 U3957 ( .IN1(n2173), .IN2(n2026), .QN(\ab[23][0] ) );
  NOR2X0 U3958 ( .IN1(n2152), .IN2(n2031), .QN(\ab[22][9] ) );
  NOR2X0 U3959 ( .IN1(n2157), .IN2(n2031), .QN(\ab[22][8] ) );
  NOR2X0 U3960 ( .IN1(n2159), .IN2(n2031), .QN(\ab[22][7] ) );
  NOR2X0 U3961 ( .IN1(n2161), .IN2(n2031), .QN(\ab[22][6] ) );
  NOR2X0 U3962 ( .IN1(n2162), .IN2(n2031), .QN(\ab[22][5] ) );
  NOR2X0 U3963 ( .IN1(n2166), .IN2(n2031), .QN(\ab[22][4] ) );
  NOR2X0 U3964 ( .IN1(n2168), .IN2(n2031), .QN(\ab[22][3] ) );
  NOR2X0 U3965 ( .IN1(A[22]), .IN2(n2094), .QN(\ab[22][31] ) );
  NOR2X0 U3966 ( .IN1(n2095), .IN2(n2030), .QN(\ab[22][30] ) );
  NOR2X0 U3967 ( .IN1(n1945), .IN2(n2030), .QN(\ab[22][2] ) );
  NOR2X0 U3968 ( .IN1(n2097), .IN2(n2030), .QN(\ab[22][29] ) );
  NOR2X0 U3969 ( .IN1(n2098), .IN2(n2030), .QN(\ab[22][28] ) );
  NOR2X0 U3970 ( .IN1(n2102), .IN2(n2030), .QN(\ab[22][27] ) );
  NOR2X0 U3971 ( .IN1(n2104), .IN2(n2030), .QN(\ab[22][26] ) );
  NOR2X0 U3972 ( .IN1(n2108), .IN2(n2030), .QN(\ab[22][25] ) );
  NOR2X0 U3973 ( .IN1(n2111), .IN2(n2030), .QN(\ab[22][24] ) );
  NOR2X0 U3974 ( .IN1(n2113), .IN2(n2030), .QN(\ab[22][23] ) );
  NOR2X0 U3975 ( .IN1(n2118), .IN2(n2030), .QN(\ab[22][22] ) );
  NOR2X0 U3976 ( .IN1(n2120), .IN2(n2030), .QN(\ab[22][21] ) );
  NOR2X0 U3977 ( .IN1(n2122), .IN2(n2030), .QN(\ab[22][20] ) );
  NOR2X0 U3978 ( .IN1(n2171), .IN2(n2029), .QN(\ab[22][1] ) );
  NOR2X0 U3979 ( .IN1(n2126), .IN2(n2029), .QN(\ab[22][19] ) );
  NOR2X0 U3980 ( .IN1(n2129), .IN2(n2029), .QN(\ab[22][18] ) );
  NOR2X0 U3981 ( .IN1(n2135), .IN2(n2029), .QN(\ab[22][16] ) );
  NOR2X0 U3982 ( .IN1(n2138), .IN2(n2029), .QN(\ab[22][15] ) );
  NOR2X0 U3983 ( .IN1(n2142), .IN2(n2029), .QN(\ab[22][14] ) );
  NOR2X0 U3984 ( .IN1(n2144), .IN2(n2029), .QN(\ab[22][13] ) );
  NOR2X0 U3985 ( .IN1(n1904), .IN2(n2029), .QN(\ab[22][12] ) );
  NOR2X0 U3986 ( .IN1(n2148), .IN2(n2029), .QN(\ab[22][11] ) );
  NOR2X0 U3987 ( .IN1(n2150), .IN2(n2029), .QN(\ab[22][10] ) );
  NOR2X0 U3988 ( .IN1(n2173), .IN2(n2029), .QN(\ab[22][0] ) );
  NOR2X0 U3989 ( .IN1(n2153), .IN2(n2034), .QN(\ab[21][9] ) );
  NOR2X0 U3990 ( .IN1(n2155), .IN2(n2034), .QN(\ab[21][8] ) );
  NOR2X0 U3991 ( .IN1(n2158), .IN2(n2034), .QN(\ab[21][7] ) );
  NOR2X0 U3992 ( .IN1(n2160), .IN2(n2034), .QN(\ab[21][6] ) );
  NOR2X0 U3993 ( .IN1(n2162), .IN2(n2034), .QN(\ab[21][5] ) );
  NOR2X0 U3994 ( .IN1(n2164), .IN2(n2034), .QN(\ab[21][4] ) );
  NOR2X0 U3995 ( .IN1(n2168), .IN2(n2034), .QN(\ab[21][3] ) );
  NOR2X0 U3996 ( .IN1(A[21]), .IN2(n2094), .QN(\ab[21][31] ) );
  NOR2X0 U3997 ( .IN1(n2096), .IN2(n2033), .QN(\ab[21][30] ) );
  NOR2X0 U3998 ( .IN1(n1946), .IN2(n2033), .QN(\ab[21][2] ) );
  NOR2X0 U3999 ( .IN1(n580), .IN2(n2033), .QN(\ab[21][29] ) );
  NOR2X0 U4000 ( .IN1(n2099), .IN2(n2033), .QN(\ab[21][28] ) );
  NOR2X0 U4001 ( .IN1(n2101), .IN2(n2033), .QN(\ab[21][27] ) );
  NOR2X0 U4002 ( .IN1(n2106), .IN2(n2033), .QN(\ab[21][26] ) );
  NOR2X0 U4003 ( .IN1(n2108), .IN2(n2033), .QN(\ab[21][25] ) );
  NOR2X0 U4004 ( .IN1(n2111), .IN2(n2033), .QN(\ab[21][24] ) );
  NOR2X0 U4005 ( .IN1(n2114), .IN2(n2033), .QN(\ab[21][23] ) );
  NOR2X0 U4006 ( .IN1(n2116), .IN2(n2033), .QN(\ab[21][22] ) );
  NOR2X0 U4007 ( .IN1(n2120), .IN2(n2033), .QN(\ab[21][21] ) );
  NOR2X0 U4008 ( .IN1(n2123), .IN2(n2033), .QN(\ab[21][20] ) );
  NOR2X0 U4009 ( .IN1(n2170), .IN2(n2032), .QN(\ab[21][1] ) );
  NOR2X0 U4010 ( .IN1(n2126), .IN2(n2032), .QN(\ab[21][19] ) );
  NOR2X0 U4011 ( .IN1(n2129), .IN2(n2032), .QN(\ab[21][18] ) );
  NOR2X0 U4012 ( .IN1(n2132), .IN2(n2032), .QN(\ab[21][17] ) );
  NOR2X0 U4013 ( .IN1(n2135), .IN2(n2032), .QN(\ab[21][16] ) );
  NOR2X0 U4014 ( .IN1(n2138), .IN2(n2032), .QN(\ab[21][15] ) );
  NOR2X0 U4015 ( .IN1(n2140), .IN2(n2032), .QN(\ab[21][14] ) );
  NOR2X0 U4016 ( .IN1(n2144), .IN2(n2032), .QN(\ab[21][13] ) );
  NOR2X0 U4017 ( .IN1(n2146), .IN2(n2032), .QN(\ab[21][12] ) );
  NOR2X0 U4018 ( .IN1(n2148), .IN2(n2032), .QN(\ab[21][11] ) );
  NOR2X0 U4019 ( .IN1(n2150), .IN2(n2032), .QN(\ab[21][10] ) );
  NOR2X0 U4020 ( .IN1(n2173), .IN2(n2032), .QN(\ab[21][0] ) );
  NOR2X0 U4021 ( .IN1(n2152), .IN2(n2037), .QN(\ab[20][9] ) );
  NOR2X0 U4022 ( .IN1(n2157), .IN2(n2037), .QN(\ab[20][8] ) );
  NOR2X0 U4023 ( .IN1(n2158), .IN2(n2037), .QN(\ab[20][7] ) );
  NOR2X0 U4024 ( .IN1(n2160), .IN2(n2037), .QN(\ab[20][6] ) );
  NOR2X0 U4025 ( .IN1(n2162), .IN2(n2037), .QN(\ab[20][5] ) );
  NOR2X0 U4026 ( .IN1(n2166), .IN2(n2037), .QN(\ab[20][4] ) );
  NOR2X0 U4027 ( .IN1(n2168), .IN2(n2037), .QN(\ab[20][3] ) );
  NOR2X0 U4028 ( .IN1(A[20]), .IN2(n2094), .QN(\ab[20][31] ) );
  NOR2X0 U4029 ( .IN1(n2095), .IN2(n2036), .QN(\ab[20][30] ) );
  NOR2X0 U4030 ( .IN1(n1945), .IN2(n2036), .QN(\ab[20][2] ) );
  NOR2X0 U4031 ( .IN1(n578), .IN2(n2036), .QN(\ab[20][29] ) );
  NOR2X0 U4032 ( .IN1(n2100), .IN2(n2036), .QN(\ab[20][28] ) );
  NOR2X0 U4033 ( .IN1(n2102), .IN2(n2036), .QN(\ab[20][27] ) );
  NOR2X0 U4034 ( .IN1(n2104), .IN2(n2036), .QN(\ab[20][26] ) );
  NOR2X0 U4035 ( .IN1(n2108), .IN2(n2036), .QN(\ab[20][25] ) );
  NOR2X0 U4036 ( .IN1(n2111), .IN2(n2036), .QN(\ab[20][24] ) );
  NOR2X0 U4037 ( .IN1(n2115), .IN2(n2036), .QN(\ab[20][23] ) );
  NOR2X0 U4038 ( .IN1(n2117), .IN2(n2036), .QN(\ab[20][22] ) );
  NOR2X0 U4039 ( .IN1(n2120), .IN2(n2036), .QN(\ab[20][21] ) );
  NOR2X0 U4040 ( .IN1(n2124), .IN2(n2036), .QN(\ab[20][20] ) );
  NOR2X0 U4041 ( .IN1(n2171), .IN2(n2035), .QN(\ab[20][1] ) );
  NOR2X0 U4042 ( .IN1(n2126), .IN2(n2035), .QN(\ab[20][19] ) );
  NOR2X0 U4043 ( .IN1(n2129), .IN2(n2035), .QN(\ab[20][18] ) );
  NOR2X0 U4044 ( .IN1(n2132), .IN2(n2035), .QN(\ab[20][17] ) );
  NOR2X0 U4045 ( .IN1(n2135), .IN2(n2035), .QN(\ab[20][16] ) );
  NOR2X0 U4046 ( .IN1(n2138), .IN2(n2035), .QN(\ab[20][15] ) );
  NOR2X0 U4047 ( .IN1(n2142), .IN2(n2035), .QN(\ab[20][14] ) );
  NOR2X0 U4048 ( .IN1(n2144), .IN2(n2035), .QN(\ab[20][13] ) );
  NOR2X0 U4049 ( .IN1(n1903), .IN2(n2035), .QN(\ab[20][12] ) );
  NOR2X0 U4050 ( .IN1(n2148), .IN2(n2035), .QN(\ab[20][11] ) );
  NOR2X0 U4051 ( .IN1(n2150), .IN2(n2035), .QN(\ab[20][10] ) );
  NOR2X0 U4052 ( .IN1(n2173), .IN2(n2035), .QN(\ab[20][0] ) );
  NOR2X0 U4053 ( .IN1(n2154), .IN2(n2003), .QN(\ab[1][9] ) );
  NOR2X0 U4054 ( .IN1(n2156), .IN2(n2002), .QN(\ab[1][8] ) );
  NOR2X0 U4055 ( .IN1(n2232), .IN2(n2091), .QN(\ab[1][7] ) );
  NOR2X0 U4056 ( .IN1(n2233), .IN2(n2091), .QN(\ab[1][6] ) );
  NOR2X0 U4057 ( .IN1(n2234), .IN2(n2003), .QN(\ab[1][5] ) );
  NOR2X0 U4058 ( .IN1(n2165), .IN2(n2091), .QN(\ab[1][4] ) );
  NOR2X0 U4059 ( .IN1(n2236), .IN2(n721), .QN(\ab[1][3] ) );
  NOR2X0 U4060 ( .IN1(n2209), .IN2(n721), .QN(\ab[1][30] ) );
  NOR2X0 U4061 ( .IN1(n2237), .IN2(n2002), .QN(\ab[1][2] ) );
  NOR2X0 U4062 ( .IN1(n2210), .IN2(n721), .QN(\ab[1][29] ) );
  NOR2X0 U4063 ( .IN1(n2099), .IN2(n2003), .QN(\ab[1][28] ) );
  NOR2X0 U4064 ( .IN1(n2103), .IN2(n2002), .QN(\ab[1][27] ) );
  NOR2X0 U4065 ( .IN1(n2105), .IN2(n2091), .QN(\ab[1][26] ) );
  NOR2X0 U4066 ( .IN1(n2108), .IN2(n2091), .QN(\ab[1][25] ) );
  NOR2X0 U4067 ( .IN1(n2111), .IN2(n2003), .QN(\ab[1][24] ) );
  NOR2X0 U4068 ( .IN1(n2114), .IN2(n2002), .QN(\ab[1][23] ) );
  NOR2X0 U4069 ( .IN1(n2117), .IN2(n721), .QN(\ab[1][22] ) );
  NOR2X0 U4070 ( .IN1(n2120), .IN2(n2003), .QN(\ab[1][21] ) );
  NOR2X0 U4071 ( .IN1(n2123), .IN2(n2091), .QN(\ab[1][20] ) );
  NOR2X0 U4072 ( .IN1(n2238), .IN2(n721), .QN(\ab[1][1] ) );
  NOR2X0 U4073 ( .IN1(n2126), .IN2(n2002), .QN(\ab[1][19] ) );
  NOR2X0 U4074 ( .IN1(n2129), .IN2(n2002), .QN(\ab[1][18] ) );
  NOR2X0 U4075 ( .IN1(n2132), .IN2(n2090), .QN(\ab[1][17] ) );
  NOR2X0 U4076 ( .IN1(n2135), .IN2(n2003), .QN(\ab[1][16] ) );
  NOR2X0 U4077 ( .IN1(n2138), .IN2(n2002), .QN(\ab[1][15] ) );
  NOR2X0 U4078 ( .IN1(n2141), .IN2(n721), .QN(\ab[1][14] ) );
  NOR2X0 U4079 ( .IN1(n2144), .IN2(n2091), .QN(\ab[1][13] ) );
  NOR2X0 U4080 ( .IN1(n2227), .IN2(n2002), .QN(\ab[1][12] ) );
  NOR2X0 U4081 ( .IN1(n2228), .IN2(n721), .QN(\ab[1][11] ) );
  NOR2X0 U4082 ( .IN1(n2153), .IN2(n2040), .QN(\ab[19][9] ) );
  NOR2X0 U4083 ( .IN1(n2155), .IN2(n2040), .QN(\ab[19][8] ) );
  NOR2X0 U4084 ( .IN1(n2159), .IN2(n2040), .QN(\ab[19][7] ) );
  NOR2X0 U4085 ( .IN1(n2161), .IN2(n2040), .QN(\ab[19][6] ) );
  NOR2X0 U4086 ( .IN1(n2162), .IN2(n2040), .QN(\ab[19][5] ) );
  NOR2X0 U4087 ( .IN1(n2164), .IN2(n2040), .QN(\ab[19][4] ) );
  NOR2X0 U4088 ( .IN1(n2168), .IN2(n2040), .QN(\ab[19][3] ) );
  NOR2X0 U4089 ( .IN1(A[19]), .IN2(n2094), .QN(\ab[19][31] ) );
  NOR2X0 U4090 ( .IN1(n2096), .IN2(n2039), .QN(\ab[19][30] ) );
  NOR2X0 U4091 ( .IN1(n1946), .IN2(n2039), .QN(\ab[19][2] ) );
  NOR2X0 U4092 ( .IN1(n579), .IN2(n2039), .QN(\ab[19][29] ) );
  NOR2X0 U4093 ( .IN1(n2098), .IN2(n2039), .QN(\ab[19][28] ) );
  NOR2X0 U4094 ( .IN1(n2101), .IN2(n2039), .QN(\ab[19][27] ) );
  NOR2X0 U4095 ( .IN1(n2106), .IN2(n2039), .QN(\ab[19][26] ) );
  NOR2X0 U4096 ( .IN1(n2108), .IN2(n2039), .QN(\ab[19][25] ) );
  NOR2X0 U4097 ( .IN1(n2111), .IN2(n2039), .QN(\ab[19][24] ) );
  NOR2X0 U4098 ( .IN1(n2113), .IN2(n2039), .QN(\ab[19][23] ) );
  NOR2X0 U4099 ( .IN1(n2118), .IN2(n2039), .QN(\ab[19][22] ) );
  NOR2X0 U4100 ( .IN1(n2120), .IN2(n2039), .QN(\ab[19][21] ) );
  NOR2X0 U4101 ( .IN1(n2122), .IN2(n2039), .QN(\ab[19][20] ) );
  NOR2X0 U4102 ( .IN1(n2170), .IN2(n2038), .QN(\ab[19][1] ) );
  NOR2X0 U4103 ( .IN1(n2126), .IN2(n2038), .QN(\ab[19][19] ) );
  NOR2X0 U4104 ( .IN1(n2129), .IN2(n2038), .QN(\ab[19][18] ) );
  NOR2X0 U4105 ( .IN1(n2132), .IN2(n2038), .QN(\ab[19][17] ) );
  NOR2X0 U4106 ( .IN1(n2135), .IN2(n2038), .QN(\ab[19][16] ) );
  NOR2X0 U4107 ( .IN1(n2138), .IN2(n2038), .QN(\ab[19][15] ) );
  NOR2X0 U4108 ( .IN1(n2140), .IN2(n2038), .QN(\ab[19][14] ) );
  NOR2X0 U4109 ( .IN1(n2144), .IN2(n2038), .QN(\ab[19][13] ) );
  NOR2X0 U4110 ( .IN1(n1904), .IN2(n2038), .QN(\ab[19][12] ) );
  NOR2X0 U4111 ( .IN1(n2148), .IN2(n2038), .QN(\ab[19][11] ) );
  NOR2X0 U4112 ( .IN1(n2173), .IN2(n2038), .QN(\ab[19][0] ) );
  NOR2X0 U4113 ( .IN1(n2152), .IN2(n2043), .QN(\ab[18][9] ) );
  NOR2X0 U4114 ( .IN1(n2157), .IN2(n2043), .QN(\ab[18][8] ) );
  NOR2X0 U4115 ( .IN1(n2158), .IN2(n2043), .QN(\ab[18][7] ) );
  NOR2X0 U4116 ( .IN1(n2160), .IN2(n2043), .QN(\ab[18][6] ) );
  NOR2X0 U4117 ( .IN1(n2162), .IN2(n2043), .QN(\ab[18][5] ) );
  NOR2X0 U4118 ( .IN1(n2166), .IN2(n2043), .QN(\ab[18][4] ) );
  NOR2X0 U4119 ( .IN1(n2168), .IN2(n2043), .QN(\ab[18][3] ) );
  NOR2X0 U4120 ( .IN1(A[18]), .IN2(n2094), .QN(\ab[18][31] ) );
  NOR2X0 U4121 ( .IN1(n2095), .IN2(n2042), .QN(\ab[18][30] ) );
  NOR2X0 U4122 ( .IN1(n2169), .IN2(n2042), .QN(\ab[18][2] ) );
  NOR2X0 U4123 ( .IN1(n2097), .IN2(n2042), .QN(\ab[18][29] ) );
  NOR2X0 U4124 ( .IN1(n2099), .IN2(n2042), .QN(\ab[18][28] ) );
  NOR2X0 U4125 ( .IN1(n2102), .IN2(n2042), .QN(\ab[18][27] ) );
  NOR2X0 U4126 ( .IN1(n2104), .IN2(n2042), .QN(\ab[18][26] ) );
  NOR2X0 U4127 ( .IN1(n2108), .IN2(n2042), .QN(\ab[18][25] ) );
  NOR2X0 U4128 ( .IN1(n2111), .IN2(n2042), .QN(\ab[18][24] ) );
  NOR2X0 U4129 ( .IN1(n2114), .IN2(n2042), .QN(\ab[18][23] ) );
  NOR2X0 U4130 ( .IN1(n2116), .IN2(n2042), .QN(\ab[18][22] ) );
  NOR2X0 U4131 ( .IN1(n2120), .IN2(n2042), .QN(\ab[18][21] ) );
  NOR2X0 U4132 ( .IN1(n2123), .IN2(n2042), .QN(\ab[18][20] ) );
  NOR2X0 U4133 ( .IN1(n2171), .IN2(n2041), .QN(\ab[18][1] ) );
  NOR2X0 U4134 ( .IN1(n2126), .IN2(n2041), .QN(\ab[18][19] ) );
  NOR2X0 U4135 ( .IN1(n2129), .IN2(n2041), .QN(\ab[18][18] ) );
  NOR2X0 U4136 ( .IN1(n2132), .IN2(n2041), .QN(\ab[18][17] ) );
  NOR2X0 U4137 ( .IN1(n2135), .IN2(n2041), .QN(\ab[18][16] ) );
  NOR2X0 U4138 ( .IN1(n2138), .IN2(n2041), .QN(\ab[18][15] ) );
  NOR2X0 U4139 ( .IN1(n2142), .IN2(n2041), .QN(\ab[18][14] ) );
  NOR2X0 U4140 ( .IN1(n2144), .IN2(n2041), .QN(\ab[18][13] ) );
  NOR2X0 U4141 ( .IN1(n2146), .IN2(n2041), .QN(\ab[18][12] ) );
  NOR2X0 U4142 ( .IN1(n2148), .IN2(n2041), .QN(\ab[18][11] ) );
  NOR2X0 U4143 ( .IN1(n2150), .IN2(n2041), .QN(\ab[18][10] ) );
  NOR2X0 U4144 ( .IN1(n2173), .IN2(n2041), .QN(\ab[18][0] ) );
  NOR2X0 U4145 ( .IN1(n2152), .IN2(n2046), .QN(\ab[17][9] ) );
  NOR2X0 U4146 ( .IN1(n2155), .IN2(n2046), .QN(\ab[17][8] ) );
  NOR2X0 U4147 ( .IN1(n2158), .IN2(n2046), .QN(\ab[17][7] ) );
  NOR2X0 U4148 ( .IN1(n2160), .IN2(n2046), .QN(\ab[17][6] ) );
  NOR2X0 U4149 ( .IN1(n2162), .IN2(n2046), .QN(\ab[17][5] ) );
  NOR2X0 U4150 ( .IN1(n2164), .IN2(n2046), .QN(\ab[17][4] ) );
  NOR2X0 U4151 ( .IN1(n2168), .IN2(n2046), .QN(\ab[17][3] ) );
  NOR2X0 U4152 ( .IN1(A[17]), .IN2(n2094), .QN(\ab[17][31] ) );
  NOR2X0 U4153 ( .IN1(n2096), .IN2(n2045), .QN(\ab[17][30] ) );
  NOR2X0 U4154 ( .IN1(n1945), .IN2(n2045), .QN(\ab[17][2] ) );
  NOR2X0 U4155 ( .IN1(n580), .IN2(n2045), .QN(\ab[17][29] ) );
  NOR2X0 U4156 ( .IN1(n2100), .IN2(n2045), .QN(\ab[17][28] ) );
  NOR2X0 U4157 ( .IN1(n2101), .IN2(n2045), .QN(\ab[17][27] ) );
  NOR2X0 U4158 ( .IN1(n2106), .IN2(n2045), .QN(\ab[17][26] ) );
  NOR2X0 U4159 ( .IN1(n2108), .IN2(n2045), .QN(\ab[17][25] ) );
  NOR2X0 U4160 ( .IN1(n2111), .IN2(n2045), .QN(\ab[17][24] ) );
  NOR2X0 U4161 ( .IN1(n2115), .IN2(n2045), .QN(\ab[17][23] ) );
  NOR2X0 U4162 ( .IN1(n2117), .IN2(n2045), .QN(\ab[17][22] ) );
  NOR2X0 U4163 ( .IN1(n2120), .IN2(n2045), .QN(\ab[17][21] ) );
  NOR2X0 U4164 ( .IN1(n2124), .IN2(n2045), .QN(\ab[17][20] ) );
  NOR2X0 U4165 ( .IN1(n2170), .IN2(n2044), .QN(\ab[17][1] ) );
  NOR2X0 U4166 ( .IN1(n2126), .IN2(n2044), .QN(\ab[17][19] ) );
  NOR2X0 U4167 ( .IN1(n2129), .IN2(n2044), .QN(\ab[17][18] ) );
  NOR2X0 U4168 ( .IN1(n2132), .IN2(n2044), .QN(\ab[17][17] ) );
  NOR2X0 U4169 ( .IN1(n2135), .IN2(n2044), .QN(\ab[17][16] ) );
  NOR2X0 U4170 ( .IN1(n2138), .IN2(n2044), .QN(\ab[17][15] ) );
  NOR2X0 U4171 ( .IN1(n2140), .IN2(n2044), .QN(\ab[17][14] ) );
  NOR2X0 U4172 ( .IN1(n2144), .IN2(n2044), .QN(\ab[17][13] ) );
  NOR2X0 U4173 ( .IN1(n1903), .IN2(n2044), .QN(\ab[17][12] ) );
  NOR2X0 U4174 ( .IN1(n2148), .IN2(n2044), .QN(\ab[17][11] ) );
  NOR2X0 U4175 ( .IN1(n2150), .IN2(n2044), .QN(\ab[17][10] ) );
  NOR2X0 U4176 ( .IN1(n2153), .IN2(n2049), .QN(\ab[16][9] ) );
  NOR2X0 U4177 ( .IN1(n2157), .IN2(n2049), .QN(\ab[16][8] ) );
  NOR2X0 U4178 ( .IN1(n2159), .IN2(n2049), .QN(\ab[16][7] ) );
  NOR2X0 U4179 ( .IN1(n2161), .IN2(n2049), .QN(\ab[16][6] ) );
  NOR2X0 U4180 ( .IN1(n2162), .IN2(n2049), .QN(\ab[16][5] ) );
  NOR2X0 U4181 ( .IN1(n2166), .IN2(n2049), .QN(\ab[16][4] ) );
  NOR2X0 U4182 ( .IN1(n2168), .IN2(n2049), .QN(\ab[16][3] ) );
  NOR2X0 U4183 ( .IN1(A[16]), .IN2(n2094), .QN(\ab[16][31] ) );
  NOR2X0 U4184 ( .IN1(n2095), .IN2(n2048), .QN(\ab[16][30] ) );
  NOR2X0 U4185 ( .IN1(n1946), .IN2(n2048), .QN(\ab[16][2] ) );
  NOR2X0 U4186 ( .IN1(n578), .IN2(n2048), .QN(\ab[16][29] ) );
  NOR2X0 U4187 ( .IN1(n2098), .IN2(n2048), .QN(\ab[16][28] ) );
  NOR2X0 U4188 ( .IN1(n2102), .IN2(n2048), .QN(\ab[16][27] ) );
  NOR2X0 U4189 ( .IN1(n2104), .IN2(n2048), .QN(\ab[16][26] ) );
  NOR2X0 U4190 ( .IN1(n2108), .IN2(n2048), .QN(\ab[16][25] ) );
  NOR2X0 U4191 ( .IN1(n2111), .IN2(n2048), .QN(\ab[16][24] ) );
  NOR2X0 U4192 ( .IN1(n2113), .IN2(n2048), .QN(\ab[16][23] ) );
  NOR2X0 U4193 ( .IN1(n2118), .IN2(n2048), .QN(\ab[16][22] ) );
  NOR2X0 U4194 ( .IN1(n2120), .IN2(n2048), .QN(\ab[16][21] ) );
  NOR2X0 U4195 ( .IN1(n2122), .IN2(n2048), .QN(\ab[16][20] ) );
  NOR2X0 U4196 ( .IN1(n2171), .IN2(n2047), .QN(\ab[16][1] ) );
  NOR2X0 U4197 ( .IN1(n2126), .IN2(n2047), .QN(\ab[16][19] ) );
  NOR2X0 U4198 ( .IN1(n2129), .IN2(n2047), .QN(\ab[16][18] ) );
  NOR2X0 U4199 ( .IN1(n2132), .IN2(n2047), .QN(\ab[16][17] ) );
  NOR2X0 U4200 ( .IN1(n2135), .IN2(n2047), .QN(\ab[16][16] ) );
  NOR2X0 U4201 ( .IN1(n2138), .IN2(n2047), .QN(\ab[16][15] ) );
  NOR2X0 U4202 ( .IN1(n2142), .IN2(n2047), .QN(\ab[16][14] ) );
  NOR2X0 U4203 ( .IN1(n2144), .IN2(n2047), .QN(\ab[16][13] ) );
  NOR2X0 U4204 ( .IN1(n1904), .IN2(n2047), .QN(\ab[16][12] ) );
  NOR2X0 U4205 ( .IN1(n2148), .IN2(n2047), .QN(\ab[16][11] ) );
  NOR2X0 U4206 ( .IN1(n2150), .IN2(n2047), .QN(\ab[16][10] ) );
  NOR2X0 U4207 ( .IN1(n2173), .IN2(n2047), .QN(\ab[16][0] ) );
  NOR2X0 U4208 ( .IN1(n2152), .IN2(n2052), .QN(\ab[15][9] ) );
  NOR2X0 U4209 ( .IN1(n2155), .IN2(n2052), .QN(\ab[15][8] ) );
  NOR2X0 U4210 ( .IN1(n2158), .IN2(n2052), .QN(\ab[15][7] ) );
  NOR2X0 U4211 ( .IN1(n2160), .IN2(n2052), .QN(\ab[15][6] ) );
  NOR2X0 U4212 ( .IN1(n2162), .IN2(n2052), .QN(\ab[15][5] ) );
  NOR2X0 U4213 ( .IN1(n2164), .IN2(n2052), .QN(\ab[15][4] ) );
  NOR2X0 U4214 ( .IN1(n2168), .IN2(n2052), .QN(\ab[15][3] ) );
  NOR2X0 U4215 ( .IN1(A[15]), .IN2(n2094), .QN(\ab[15][31] ) );
  NOR2X0 U4216 ( .IN1(n2096), .IN2(n2051), .QN(\ab[15][30] ) );
  NOR2X0 U4217 ( .IN1(n2169), .IN2(n2051), .QN(\ab[15][2] ) );
  NOR2X0 U4218 ( .IN1(n579), .IN2(n2051), .QN(\ab[15][29] ) );
  NOR2X0 U4219 ( .IN1(n2099), .IN2(n2051), .QN(\ab[15][28] ) );
  NOR2X0 U4220 ( .IN1(n2101), .IN2(n2051), .QN(\ab[15][27] ) );
  NOR2X0 U4221 ( .IN1(n2106), .IN2(n2051), .QN(\ab[15][26] ) );
  NOR2X0 U4222 ( .IN1(n2108), .IN2(n2051), .QN(\ab[15][25] ) );
  NOR2X0 U4223 ( .IN1(n2111), .IN2(n2051), .QN(\ab[15][24] ) );
  NOR2X0 U4224 ( .IN1(n2114), .IN2(n2051), .QN(\ab[15][23] ) );
  NOR2X0 U4225 ( .IN1(n2116), .IN2(n2051), .QN(\ab[15][22] ) );
  NOR2X0 U4226 ( .IN1(n2120), .IN2(n2051), .QN(\ab[15][21] ) );
  NOR2X0 U4227 ( .IN1(n2123), .IN2(n2051), .QN(\ab[15][20] ) );
  NOR2X0 U4228 ( .IN1(n2170), .IN2(n2050), .QN(\ab[15][1] ) );
  NOR2X0 U4229 ( .IN1(n2126), .IN2(n2050), .QN(\ab[15][19] ) );
  NOR2X0 U4230 ( .IN1(n2129), .IN2(n2050), .QN(\ab[15][18] ) );
  NOR2X0 U4231 ( .IN1(n2132), .IN2(n2050), .QN(\ab[15][17] ) );
  NOR2X0 U4232 ( .IN1(n2135), .IN2(n2050), .QN(\ab[15][16] ) );
  NOR2X0 U4233 ( .IN1(n2138), .IN2(n2050), .QN(\ab[15][15] ) );
  NOR2X0 U4234 ( .IN1(n2140), .IN2(n2050), .QN(\ab[15][14] ) );
  NOR2X0 U4235 ( .IN1(n2144), .IN2(n2050), .QN(\ab[15][13] ) );
  NOR2X0 U4236 ( .IN1(n2146), .IN2(n2050), .QN(\ab[15][12] ) );
  NOR2X0 U4237 ( .IN1(n2148), .IN2(n2050), .QN(\ab[15][11] ) );
  NOR2X0 U4238 ( .IN1(n2150), .IN2(n2050), .QN(\ab[15][10] ) );
  NOR2X0 U4239 ( .IN1(n2153), .IN2(n2055), .QN(\ab[14][9] ) );
  NOR2X0 U4240 ( .IN1(n2157), .IN2(n2055), .QN(\ab[14][8] ) );
  NOR2X0 U4241 ( .IN1(n2158), .IN2(n2055), .QN(\ab[14][7] ) );
  NOR2X0 U4242 ( .IN1(n2160), .IN2(n2055), .QN(\ab[14][6] ) );
  NOR2X0 U4243 ( .IN1(n2162), .IN2(n2055), .QN(\ab[14][5] ) );
  NOR2X0 U4244 ( .IN1(n2166), .IN2(n2055), .QN(\ab[14][4] ) );
  NOR2X0 U4245 ( .IN1(n2168), .IN2(n2055), .QN(\ab[14][3] ) );
  NOR2X0 U4246 ( .IN1(A[14]), .IN2(n2094), .QN(\ab[14][31] ) );
  NOR2X0 U4247 ( .IN1(n2095), .IN2(n2054), .QN(\ab[14][30] ) );
  NOR2X0 U4248 ( .IN1(n1945), .IN2(n2054), .QN(\ab[14][2] ) );
  NOR2X0 U4249 ( .IN1(n2097), .IN2(n2054), .QN(\ab[14][29] ) );
  NOR2X0 U4250 ( .IN1(n2100), .IN2(n2054), .QN(\ab[14][28] ) );
  NOR2X0 U4251 ( .IN1(n2102), .IN2(n2054), .QN(\ab[14][27] ) );
  NOR2X0 U4252 ( .IN1(n2104), .IN2(n2054), .QN(\ab[14][26] ) );
  NOR2X0 U4253 ( .IN1(n2108), .IN2(n2054), .QN(\ab[14][25] ) );
  NOR2X0 U4254 ( .IN1(n2111), .IN2(n2054), .QN(\ab[14][24] ) );
  NOR2X0 U4255 ( .IN1(n2115), .IN2(n2054), .QN(\ab[14][23] ) );
  NOR2X0 U4256 ( .IN1(n2117), .IN2(n2054), .QN(\ab[14][22] ) );
  NOR2X0 U4257 ( .IN1(n2120), .IN2(n2054), .QN(\ab[14][21] ) );
  NOR2X0 U4258 ( .IN1(n2124), .IN2(n2054), .QN(\ab[14][20] ) );
  NOR2X0 U4259 ( .IN1(n2171), .IN2(n2053), .QN(\ab[14][1] ) );
  NOR2X0 U4260 ( .IN1(n2126), .IN2(n2053), .QN(\ab[14][19] ) );
  NOR2X0 U4261 ( .IN1(n2129), .IN2(n2053), .QN(\ab[14][18] ) );
  NOR2X0 U4262 ( .IN1(n2132), .IN2(n2053), .QN(\ab[14][17] ) );
  NOR2X0 U4263 ( .IN1(n2135), .IN2(n2053), .QN(\ab[14][16] ) );
  NOR2X0 U4264 ( .IN1(n2138), .IN2(n2053), .QN(\ab[14][15] ) );
  NOR2X0 U4265 ( .IN1(n2142), .IN2(n2053), .QN(\ab[14][14] ) );
  NOR2X0 U4266 ( .IN1(n2144), .IN2(n2053), .QN(\ab[14][13] ) );
  NOR2X0 U4267 ( .IN1(n1903), .IN2(n2053), .QN(\ab[14][12] ) );
  NOR2X0 U4268 ( .IN1(n2148), .IN2(n2053), .QN(\ab[14][11] ) );
  NOR2X0 U4269 ( .IN1(n2150), .IN2(n2053), .QN(\ab[14][10] ) );
  NOR2X0 U4270 ( .IN1(n2173), .IN2(n2053), .QN(\ab[14][0] ) );
  NOR2X0 U4271 ( .IN1(n2152), .IN2(n2058), .QN(\ab[13][9] ) );
  NOR2X0 U4272 ( .IN1(n2155), .IN2(n2058), .QN(\ab[13][8] ) );
  NOR2X0 U4273 ( .IN1(n2159), .IN2(n2058), .QN(\ab[13][7] ) );
  NOR2X0 U4274 ( .IN1(n2161), .IN2(n2058), .QN(\ab[13][6] ) );
  NOR2X0 U4275 ( .IN1(n2163), .IN2(n2058), .QN(\ab[13][5] ) );
  NOR2X0 U4276 ( .IN1(n2164), .IN2(n2058), .QN(\ab[13][4] ) );
  NOR2X0 U4277 ( .IN1(n2168), .IN2(n2058), .QN(\ab[13][3] ) );
  NOR2X0 U4278 ( .IN1(A[13]), .IN2(n2094), .QN(\ab[13][31] ) );
  NOR2X0 U4279 ( .IN1(n2096), .IN2(n2057), .QN(\ab[13][30] ) );
  NOR2X0 U4280 ( .IN1(n1946), .IN2(n2057), .QN(\ab[13][2] ) );
  NOR2X0 U4281 ( .IN1(n580), .IN2(n2057), .QN(\ab[13][29] ) );
  NOR2X0 U4282 ( .IN1(n2098), .IN2(n2057), .QN(\ab[13][28] ) );
  NOR2X0 U4283 ( .IN1(n2101), .IN2(n2057), .QN(\ab[13][27] ) );
  NOR2X0 U4284 ( .IN1(n2106), .IN2(n2057), .QN(\ab[13][26] ) );
  NOR2X0 U4285 ( .IN1(n2109), .IN2(n2057), .QN(\ab[13][25] ) );
  NOR2X0 U4286 ( .IN1(n2112), .IN2(n2057), .QN(\ab[13][24] ) );
  NOR2X0 U4287 ( .IN1(n2113), .IN2(n2057), .QN(\ab[13][23] ) );
  NOR2X0 U4288 ( .IN1(n2118), .IN2(n2057), .QN(\ab[13][22] ) );
  NOR2X0 U4289 ( .IN1(n2121), .IN2(n2057), .QN(\ab[13][21] ) );
  NOR2X0 U4290 ( .IN1(n2122), .IN2(n2057), .QN(\ab[13][20] ) );
  NOR2X0 U4291 ( .IN1(n2170), .IN2(n2056), .QN(\ab[13][1] ) );
  NOR2X0 U4292 ( .IN1(n2127), .IN2(n2056), .QN(\ab[13][19] ) );
  NOR2X0 U4293 ( .IN1(n2130), .IN2(n2056), .QN(\ab[13][18] ) );
  NOR2X0 U4294 ( .IN1(n2133), .IN2(n2056), .QN(\ab[13][17] ) );
  NOR2X0 U4295 ( .IN1(n2136), .IN2(n2056), .QN(\ab[13][16] ) );
  NOR2X0 U4296 ( .IN1(n2139), .IN2(n2056), .QN(\ab[13][15] ) );
  NOR2X0 U4297 ( .IN1(n2140), .IN2(n2056), .QN(\ab[13][14] ) );
  NOR2X0 U4298 ( .IN1(n2145), .IN2(n2056), .QN(\ab[13][13] ) );
  NOR2X0 U4299 ( .IN1(n1904), .IN2(n2056), .QN(\ab[13][12] ) );
  NOR2X0 U4300 ( .IN1(n2148), .IN2(n2056), .QN(\ab[13][11] ) );
  NOR2X0 U4301 ( .IN1(n2151), .IN2(n2056), .QN(\ab[13][10] ) );
  NOR2X0 U4302 ( .IN1(n2174), .IN2(n2056), .QN(\ab[13][0] ) );
  NOR2X0 U4303 ( .IN1(n2153), .IN2(n2061), .QN(\ab[12][9] ) );
  NOR2X0 U4304 ( .IN1(n2157), .IN2(n2061), .QN(\ab[12][8] ) );
  NOR2X0 U4305 ( .IN1(n2158), .IN2(n2061), .QN(\ab[12][7] ) );
  NOR2X0 U4306 ( .IN1(n2160), .IN2(n2061), .QN(\ab[12][6] ) );
  NOR2X0 U4307 ( .IN1(n2163), .IN2(n2061), .QN(\ab[12][5] ) );
  NOR2X0 U4308 ( .IN1(n2166), .IN2(n2061), .QN(\ab[12][4] ) );
  NOR2X0 U4309 ( .IN1(n2168), .IN2(n2061), .QN(\ab[12][3] ) );
  NOR2X0 U4310 ( .IN1(A[12]), .IN2(n2094), .QN(\ab[12][31] ) );
  NOR2X0 U4311 ( .IN1(n2095), .IN2(n2060), .QN(\ab[12][30] ) );
  NOR2X0 U4312 ( .IN1(n2169), .IN2(n2060), .QN(\ab[12][2] ) );
  NOR2X0 U4313 ( .IN1(n578), .IN2(n2060), .QN(\ab[12][29] ) );
  NOR2X0 U4314 ( .IN1(n2099), .IN2(n2060), .QN(\ab[12][28] ) );
  NOR2X0 U4315 ( .IN1(n2102), .IN2(n2060), .QN(\ab[12][27] ) );
  NOR2X0 U4316 ( .IN1(n2104), .IN2(n2060), .QN(\ab[12][26] ) );
  NOR2X0 U4317 ( .IN1(n2109), .IN2(n2060), .QN(\ab[12][25] ) );
  NOR2X0 U4318 ( .IN1(n2112), .IN2(n2060), .QN(\ab[12][24] ) );
  NOR2X0 U4319 ( .IN1(n2114), .IN2(n2060), .QN(\ab[12][23] ) );
  NOR2X0 U4320 ( .IN1(n2117), .IN2(n2060), .QN(\ab[12][22] ) );
  NOR2X0 U4321 ( .IN1(n2121), .IN2(n2060), .QN(\ab[12][21] ) );
  NOR2X0 U4322 ( .IN1(n2123), .IN2(n2060), .QN(\ab[12][20] ) );
  NOR2X0 U4323 ( .IN1(n2171), .IN2(n2059), .QN(\ab[12][1] ) );
  NOR2X0 U4324 ( .IN1(n2127), .IN2(n2059), .QN(\ab[12][19] ) );
  NOR2X0 U4325 ( .IN1(n2130), .IN2(n2059), .QN(\ab[12][18] ) );
  NOR2X0 U4326 ( .IN1(n2133), .IN2(n2059), .QN(\ab[12][17] ) );
  NOR2X0 U4327 ( .IN1(n2136), .IN2(n2059), .QN(\ab[12][16] ) );
  NOR2X0 U4328 ( .IN1(n2139), .IN2(n2059), .QN(\ab[12][15] ) );
  NOR2X0 U4329 ( .IN1(n2142), .IN2(n2059), .QN(\ab[12][14] ) );
  NOR2X0 U4330 ( .IN1(n2145), .IN2(n2059), .QN(\ab[12][13] ) );
  NOR2X0 U4331 ( .IN1(n2146), .IN2(n2059), .QN(\ab[12][12] ) );
  NOR2X0 U4332 ( .IN1(n2148), .IN2(n2059), .QN(\ab[12][11] ) );
  NOR2X0 U4333 ( .IN1(n2151), .IN2(n2059), .QN(\ab[12][10] ) );
  NOR2X0 U4334 ( .IN1(n2174), .IN2(n2059), .QN(\ab[12][0] ) );
  NOR2X0 U4335 ( .IN1(n2152), .IN2(n2064), .QN(\ab[11][9] ) );
  NOR2X0 U4336 ( .IN1(n2155), .IN2(n2064), .QN(\ab[11][8] ) );
  NOR2X0 U4337 ( .IN1(n2158), .IN2(n2064), .QN(\ab[11][7] ) );
  NOR2X0 U4338 ( .IN1(n2160), .IN2(n2064), .QN(\ab[11][6] ) );
  NOR2X0 U4339 ( .IN1(n2163), .IN2(n2064), .QN(\ab[11][5] ) );
  NOR2X0 U4340 ( .IN1(n2164), .IN2(n2064), .QN(\ab[11][4] ) );
  NOR2X0 U4341 ( .IN1(n2168), .IN2(n2064), .QN(\ab[11][3] ) );
  NOR2X0 U4342 ( .IN1(A[11]), .IN2(n2094), .QN(\ab[11][31] ) );
  NOR2X0 U4343 ( .IN1(n2096), .IN2(n2063), .QN(\ab[11][30] ) );
  NOR2X0 U4344 ( .IN1(n1945), .IN2(n2063), .QN(\ab[11][2] ) );
  NOR2X0 U4345 ( .IN1(n579), .IN2(n2063), .QN(\ab[11][29] ) );
  NOR2X0 U4346 ( .IN1(n2100), .IN2(n2063), .QN(\ab[11][28] ) );
  NOR2X0 U4347 ( .IN1(n2101), .IN2(n2063), .QN(\ab[11][27] ) );
  NOR2X0 U4348 ( .IN1(n2106), .IN2(n2063), .QN(\ab[11][26] ) );
  NOR2X0 U4349 ( .IN1(n2109), .IN2(n2063), .QN(\ab[11][25] ) );
  NOR2X0 U4350 ( .IN1(n2112), .IN2(n2063), .QN(\ab[11][24] ) );
  NOR2X0 U4351 ( .IN1(n2115), .IN2(n2063), .QN(\ab[11][23] ) );
  NOR2X0 U4352 ( .IN1(n2118), .IN2(n2063), .QN(\ab[11][22] ) );
  NOR2X0 U4353 ( .IN1(n2121), .IN2(n2063), .QN(\ab[11][21] ) );
  NOR2X0 U4354 ( .IN1(n2124), .IN2(n2063), .QN(\ab[11][20] ) );
  NOR2X0 U4355 ( .IN1(n2170), .IN2(n2062), .QN(\ab[11][1] ) );
  NOR2X0 U4356 ( .IN1(n2127), .IN2(n2062), .QN(\ab[11][19] ) );
  NOR2X0 U4357 ( .IN1(n2130), .IN2(n2062), .QN(\ab[11][18] ) );
  NOR2X0 U4358 ( .IN1(n2133), .IN2(n2062), .QN(\ab[11][17] ) );
  NOR2X0 U4359 ( .IN1(n2136), .IN2(n2062), .QN(\ab[11][16] ) );
  NOR2X0 U4360 ( .IN1(n2139), .IN2(n2062), .QN(\ab[11][15] ) );
  NOR2X0 U4361 ( .IN1(n2140), .IN2(n2062), .QN(\ab[11][14] ) );
  NOR2X0 U4362 ( .IN1(n2145), .IN2(n2062), .QN(\ab[11][13] ) );
  NOR2X0 U4363 ( .IN1(n1903), .IN2(n2062), .QN(\ab[11][12] ) );
  NOR2X0 U4364 ( .IN1(n2148), .IN2(n2062), .QN(\ab[11][11] ) );
  NOR2X0 U4365 ( .IN1(n2151), .IN2(n2062), .QN(\ab[11][10] ) );
  NOR2X0 U4366 ( .IN1(n2174), .IN2(n2062), .QN(\ab[11][0] ) );
  NOR2X0 U4367 ( .IN1(n2153), .IN2(n2067), .QN(\ab[10][9] ) );
  NOR2X0 U4368 ( .IN1(n2161), .IN2(n2067), .QN(\ab[10][6] ) );
  NOR2X0 U4369 ( .IN1(n2163), .IN2(n2067), .QN(\ab[10][5] ) );
  NOR2X0 U4370 ( .IN1(n2166), .IN2(n2067), .QN(\ab[10][4] ) );
  NOR2X0 U4371 ( .IN1(n2168), .IN2(n2067), .QN(\ab[10][3] ) );
  NOR2X0 U4372 ( .IN1(A[10]), .IN2(n2094), .QN(\ab[10][31] ) );
  NOR2X0 U4373 ( .IN1(n2095), .IN2(n2066), .QN(\ab[10][30] ) );
  NOR2X0 U4374 ( .IN1(n1946), .IN2(n2066), .QN(\ab[10][2] ) );
  NOR2X0 U4375 ( .IN1(n2097), .IN2(n2066), .QN(\ab[10][29] ) );
  NOR2X0 U4376 ( .IN1(n2098), .IN2(n2066), .QN(\ab[10][28] ) );
  NOR2X0 U4377 ( .IN1(n2102), .IN2(n2066), .QN(\ab[10][27] ) );
  NOR2X0 U4378 ( .IN1(n2104), .IN2(n2066), .QN(\ab[10][26] ) );
  NOR2X0 U4379 ( .IN1(n2109), .IN2(n2066), .QN(\ab[10][25] ) );
  NOR2X0 U4380 ( .IN1(n2112), .IN2(n2066), .QN(\ab[10][24] ) );
  NOR2X0 U4381 ( .IN1(n2113), .IN2(n2066), .QN(\ab[10][23] ) );
  NOR2X0 U4382 ( .IN1(n2116), .IN2(n2066), .QN(\ab[10][22] ) );
  NOR2X0 U4383 ( .IN1(n2121), .IN2(n2066), .QN(\ab[10][21] ) );
  NOR2X0 U4384 ( .IN1(n2122), .IN2(n2066), .QN(\ab[10][20] ) );
  NOR2X0 U4385 ( .IN1(n2171), .IN2(n2065), .QN(\ab[10][1] ) );
  NOR2X0 U4386 ( .IN1(n2127), .IN2(n2065), .QN(\ab[10][19] ) );
  NOR2X0 U4387 ( .IN1(n2130), .IN2(n2065), .QN(\ab[10][18] ) );
  NOR2X0 U4388 ( .IN1(n2133), .IN2(n2065), .QN(\ab[10][17] ) );
  NOR2X0 U4389 ( .IN1(n2136), .IN2(n2065), .QN(\ab[10][16] ) );
  NOR2X0 U4390 ( .IN1(n2139), .IN2(n2065), .QN(\ab[10][15] ) );
  NOR2X0 U4391 ( .IN1(n2142), .IN2(n2065), .QN(\ab[10][14] ) );
  NOR2X0 U4392 ( .IN1(n2145), .IN2(n2065), .QN(\ab[10][13] ) );
  NOR2X0 U4393 ( .IN1(n1904), .IN2(n2065), .QN(\ab[10][12] ) );
  NOR2X0 U4394 ( .IN1(n2148), .IN2(n2065), .QN(\ab[10][11] ) );
  NOR2X0 U4395 ( .IN1(n2151), .IN2(n2065), .QN(\ab[10][10] ) );
  NOR2X0 U4396 ( .IN1(n2174), .IN2(n2065), .QN(\ab[10][0] ) );
  NOR2X0 U4397 ( .IN1(n2154), .IN2(n2093), .QN(\ab[0][9] ) );
  NOR2X0 U4398 ( .IN1(n2156), .IN2(n2093), .QN(\ab[0][8] ) );
  NOR2X0 U4399 ( .IN1(n2159), .IN2(n2093), .QN(\ab[0][7] ) );
  NOR2X0 U4400 ( .IN1(n2161), .IN2(n2093), .QN(\ab[0][6] ) );
  NOR2X0 U4401 ( .IN1(n2163), .IN2(n2207), .QN(\ab[0][5] ) );
  NOR2X0 U4402 ( .IN1(n2165), .IN2(n2092), .QN(\ab[0][4] ) );
  NOR2X0 U4403 ( .IN1(n2167), .IN2(n2093), .QN(\ab[0][3] ) );
  NOR2X0 U4404 ( .IN1(n599), .IN2(n2208), .QN(\ab[0][31] ) );
  NOR2X0 U4405 ( .IN1(n2237), .IN2(n2207), .QN(\ab[0][2] ) );
  NOR2X0 U4406 ( .IN1(n2097), .IN2(n2093), .QN(\ab[0][29] ) );
  NOR2X0 U4407 ( .IN1(n2103), .IN2(n2092), .QN(\ab[0][27] ) );
  NOR2X0 U4408 ( .IN1(n2105), .IN2(n2093), .QN(\ab[0][26] ) );
  NOR2X0 U4409 ( .IN1(n2109), .IN2(n2093), .QN(\ab[0][25] ) );
  NOR2X0 U4410 ( .IN1(n2112), .IN2(n2093), .QN(\ab[0][24] ) );
  NOR2X0 U4411 ( .IN1(n2113), .IN2(n2093), .QN(\ab[0][23] ) );
  NOR2X0 U4412 ( .IN1(n2118), .IN2(n2207), .QN(\ab[0][22] ) );
  NOR2X0 U4413 ( .IN1(n2121), .IN2(n2093), .QN(\ab[0][21] ) );
  NOR2X0 U4414 ( .IN1(n2124), .IN2(n2092), .QN(\ab[0][20] ) );
  NOR2X0 U4415 ( .IN1(n2171), .IN2(n2093), .QN(\ab[0][1] ) );
  NOR2X0 U4416 ( .IN1(n2127), .IN2(n2207), .QN(\ab[0][19] ) );
  NOR2X0 U4417 ( .IN1(n2130), .IN2(n2207), .QN(\ab[0][18] ) );
  NOR2X0 U4418 ( .IN1(n2133), .IN2(n2207), .QN(\ab[0][17] ) );
  NOR2X0 U4419 ( .IN1(n2136), .IN2(n2207), .QN(\ab[0][16] ) );
  NOR2X0 U4420 ( .IN1(n2139), .IN2(n2207), .QN(\ab[0][15] ) );
  NOR2X0 U4421 ( .IN1(n2141), .IN2(n2207), .QN(\ab[0][14] ) );
  NOR2X0 U4422 ( .IN1(n2145), .IN2(n2207), .QN(\ab[0][13] ) );
  NOR2X0 U4423 ( .IN1(n2227), .IN2(n1971), .QN(\ab[0][12] ) );
  NOR2X0 U4424 ( .IN1(n2147), .IN2(n2093), .QN(\ab[0][11] ) );
  NOR2X0 U4425 ( .IN1(n2151), .IN2(n2207), .QN(\ab[0][10] ) );
  NOR2X0 U4426 ( .IN1(n2174), .IN2(n2207), .QN(PRODUCT[0]) );
endmodule


module VerilogMultiplier ( clk, rst, A, B, P );
  input [31:0] A;
  input [31:0] B;
  output [63:0] P;
  input clk, rst;
  wire   N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [31:0] B_reg;
  wire   [31:0] A_reg;

  DFFARX1 \A_reg_reg[31]  ( .D(A[31]), .CLK(clk), .RSTB(n19), .Q(A_reg[31]) );
  DFFARX1 \A_reg_reg[30]  ( .D(A[30]), .CLK(clk), .RSTB(n19), .Q(A_reg[30]) );
  DFFARX1 \A_reg_reg[29]  ( .D(A[29]), .CLK(clk), .RSTB(n19), .Q(A_reg[29]) );
  DFFARX1 \A_reg_reg[28]  ( .D(A[28]), .CLK(clk), .RSTB(n19), .Q(A_reg[28]) );
  DFFARX1 \A_reg_reg[27]  ( .D(A[27]), .CLK(clk), .RSTB(n19), .Q(A_reg[27]) );
  DFFARX1 \A_reg_reg[26]  ( .D(A[26]), .CLK(clk), .RSTB(n19), .Q(A_reg[26]) );
  DFFARX1 \A_reg_reg[25]  ( .D(A[25]), .CLK(clk), .RSTB(n19), .Q(A_reg[25]) );
  DFFARX1 \A_reg_reg[24]  ( .D(A[24]), .CLK(clk), .RSTB(n19), .Q(A_reg[24]) );
  DFFARX1 \A_reg_reg[23]  ( .D(A[23]), .CLK(clk), .RSTB(n18), .Q(A_reg[23]) );
  DFFARX1 \A_reg_reg[22]  ( .D(A[22]), .CLK(clk), .RSTB(n18), .Q(A_reg[22]) );
  DFFARX1 \A_reg_reg[21]  ( .D(A[21]), .CLK(clk), .RSTB(n18), .Q(A_reg[21]) );
  DFFARX1 \A_reg_reg[20]  ( .D(A[20]), .CLK(clk), .RSTB(n18), .Q(A_reg[20]) );
  DFFARX1 \A_reg_reg[19]  ( .D(A[19]), .CLK(clk), .RSTB(n18), .Q(A_reg[19]) );
  DFFARX1 \A_reg_reg[18]  ( .D(A[18]), .CLK(clk), .RSTB(n18), .Q(A_reg[18]) );
  DFFARX1 \A_reg_reg[17]  ( .D(A[17]), .CLK(clk), .RSTB(n18), .Q(A_reg[17]) );
  DFFARX1 \A_reg_reg[16]  ( .D(A[16]), .CLK(clk), .RSTB(n18), .Q(A_reg[16]) );
  DFFARX1 \A_reg_reg[15]  ( .D(A[15]), .CLK(clk), .RSTB(n18), .Q(A_reg[15]) );
  DFFARX1 \A_reg_reg[14]  ( .D(A[14]), .CLK(clk), .RSTB(n18), .Q(A_reg[14]) );
  DFFARX1 \A_reg_reg[13]  ( .D(A[13]), .CLK(clk), .RSTB(n17), .Q(A_reg[13]) );
  DFFARX1 \A_reg_reg[12]  ( .D(A[12]), .CLK(clk), .RSTB(n17), .Q(A_reg[12]) );
  DFFARX1 \A_reg_reg[11]  ( .D(A[11]), .CLK(clk), .RSTB(n17), .Q(A_reg[11]) );
  DFFARX1 \A_reg_reg[10]  ( .D(A[10]), .CLK(clk), .RSTB(n17), .Q(A_reg[10]) );
  DFFARX1 \A_reg_reg[9]  ( .D(A[9]), .CLK(clk), .RSTB(n17), .Q(A_reg[9]) );
  DFFARX1 \A_reg_reg[8]  ( .D(A[8]), .CLK(clk), .RSTB(n17), .Q(A_reg[8]) );
  DFFARX1 \A_reg_reg[7]  ( .D(A[7]), .CLK(clk), .RSTB(n17), .Q(A_reg[7]) );
  DFFARX1 \A_reg_reg[6]  ( .D(A[6]), .CLK(clk), .RSTB(n17), .Q(A_reg[6]) );
  DFFARX1 \A_reg_reg[5]  ( .D(A[5]), .CLK(clk), .RSTB(n17), .Q(A_reg[5]) );
  DFFARX1 \A_reg_reg[4]  ( .D(A[4]), .CLK(clk), .RSTB(n17), .Q(A_reg[4]) );
  DFFARX1 \A_reg_reg[3]  ( .D(A[3]), .CLK(clk), .RSTB(n16), .Q(A_reg[3]) );
  DFFARX1 \A_reg_reg[2]  ( .D(A[2]), .CLK(clk), .RSTB(n16), .Q(A_reg[2]) );
  DFFARX1 \A_reg_reg[1]  ( .D(A[1]), .CLK(clk), .RSTB(n16), .Q(A_reg[1]) );
  DFFARX1 \A_reg_reg[0]  ( .D(A[0]), .CLK(clk), .RSTB(n16), .Q(A_reg[0]) );
  DFFARX1 \P_reg_reg[63]  ( .D(N64), .CLK(clk), .RSTB(n16), .Q(P[63]) );
  DFFARX1 \P_reg_reg[62]  ( .D(N63), .CLK(clk), .RSTB(n16), .Q(P[62]) );
  DFFARX1 \P_reg_reg[61]  ( .D(N62), .CLK(clk), .RSTB(n16), .Q(P[61]) );
  DFFARX1 \P_reg_reg[60]  ( .D(N61), .CLK(clk), .RSTB(n16), .Q(P[60]) );
  DFFARX1 \P_reg_reg[59]  ( .D(N60), .CLK(clk), .RSTB(n16), .Q(P[59]) );
  DFFARX1 \P_reg_reg[58]  ( .D(N59), .CLK(clk), .RSTB(n16), .Q(P[58]) );
  DFFARX1 \P_reg_reg[57]  ( .D(N58), .CLK(clk), .RSTB(n15), .Q(P[57]) );
  DFFARX1 \P_reg_reg[56]  ( .D(N57), .CLK(clk), .RSTB(n15), .Q(P[56]) );
  DFFARX1 \P_reg_reg[55]  ( .D(N56), .CLK(clk), .RSTB(n15), .Q(P[55]) );
  DFFARX1 \P_reg_reg[54]  ( .D(N55), .CLK(clk), .RSTB(n15), .Q(P[54]) );
  DFFARX1 \P_reg_reg[53]  ( .D(N54), .CLK(clk), .RSTB(n15), .Q(P[53]) );
  DFFARX1 \P_reg_reg[52]  ( .D(N53), .CLK(clk), .RSTB(n15), .Q(P[52]) );
  DFFARX1 \P_reg_reg[51]  ( .D(N52), .CLK(clk), .RSTB(n15), .Q(P[51]) );
  DFFARX1 \P_reg_reg[50]  ( .D(N51), .CLK(clk), .RSTB(n15), .Q(P[50]) );
  DFFARX1 \P_reg_reg[49]  ( .D(N50), .CLK(clk), .RSTB(n15), .Q(P[49]) );
  DFFARX1 \P_reg_reg[48]  ( .D(N49), .CLK(clk), .RSTB(n15), .Q(P[48]) );
  DFFARX1 \P_reg_reg[47]  ( .D(N48), .CLK(clk), .RSTB(n14), .Q(P[47]) );
  DFFARX1 \P_reg_reg[46]  ( .D(N47), .CLK(clk), .RSTB(n14), .Q(P[46]) );
  DFFARX1 \P_reg_reg[45]  ( .D(N46), .CLK(clk), .RSTB(n14), .Q(P[45]) );
  DFFARX1 \P_reg_reg[44]  ( .D(N45), .CLK(clk), .RSTB(n14), .Q(P[44]) );
  DFFARX1 \P_reg_reg[43]  ( .D(N44), .CLK(clk), .RSTB(n14), .Q(P[43]) );
  DFFARX1 \P_reg_reg[42]  ( .D(N43), .CLK(clk), .RSTB(n14), .Q(P[42]) );
  DFFARX1 \P_reg_reg[41]  ( .D(N42), .CLK(clk), .RSTB(n14), .Q(P[41]) );
  DFFARX1 \P_reg_reg[40]  ( .D(N41), .CLK(clk), .RSTB(n14), .Q(P[40]) );
  DFFARX1 \P_reg_reg[39]  ( .D(N40), .CLK(clk), .RSTB(n14), .Q(P[39]) );
  DFFARX1 \P_reg_reg[38]  ( .D(N39), .CLK(clk), .RSTB(n14), .Q(P[38]) );
  DFFARX1 \P_reg_reg[37]  ( .D(N38), .CLK(clk), .RSTB(n13), .Q(P[37]) );
  DFFARX1 \P_reg_reg[36]  ( .D(N37), .CLK(clk), .RSTB(n13), .Q(P[36]) );
  DFFARX1 \P_reg_reg[35]  ( .D(N36), .CLK(clk), .RSTB(n13), .Q(P[35]) );
  DFFARX1 \P_reg_reg[34]  ( .D(N35), .CLK(clk), .RSTB(n13), .Q(P[34]) );
  DFFARX1 \P_reg_reg[33]  ( .D(N34), .CLK(clk), .RSTB(n13), .Q(P[33]) );
  DFFARX1 \P_reg_reg[32]  ( .D(N33), .CLK(clk), .RSTB(n13), .Q(P[32]) );
  DFFARX1 \P_reg_reg[31]  ( .D(N32), .CLK(clk), .RSTB(n13), .Q(P[31]) );
  DFFARX1 \P_reg_reg[30]  ( .D(N31), .CLK(clk), .RSTB(n13), .Q(P[30]) );
  DFFARX1 \P_reg_reg[29]  ( .D(N30), .CLK(clk), .RSTB(n13), .Q(P[29]) );
  DFFARX1 \P_reg_reg[28]  ( .D(N29), .CLK(clk), .RSTB(n13), .Q(P[28]) );
  DFFARX1 \P_reg_reg[27]  ( .D(N28), .CLK(clk), .RSTB(n12), .Q(P[27]) );
  DFFARX1 \P_reg_reg[26]  ( .D(N27), .CLK(clk), .RSTB(n12), .Q(P[26]) );
  DFFARX1 \P_reg_reg[25]  ( .D(N26), .CLK(clk), .RSTB(n12), .Q(P[25]) );
  DFFARX1 \P_reg_reg[24]  ( .D(N25), .CLK(clk), .RSTB(n12), .Q(P[24]) );
  DFFARX1 \P_reg_reg[23]  ( .D(N24), .CLK(clk), .RSTB(n12), .Q(P[23]) );
  DFFARX1 \P_reg_reg[22]  ( .D(N23), .CLK(clk), .RSTB(n12), .Q(P[22]) );
  DFFARX1 \P_reg_reg[21]  ( .D(N22), .CLK(clk), .RSTB(n12), .Q(P[21]) );
  DFFARX1 \P_reg_reg[20]  ( .D(N21), .CLK(clk), .RSTB(n12), .Q(P[20]) );
  DFFARX1 \P_reg_reg[19]  ( .D(N20), .CLK(clk), .RSTB(n12), .Q(P[19]) );
  DFFARX1 \P_reg_reg[18]  ( .D(N19), .CLK(clk), .RSTB(n12), .Q(P[18]) );
  DFFARX1 \P_reg_reg[17]  ( .D(N18), .CLK(clk), .RSTB(n11), .Q(P[17]) );
  DFFARX1 \P_reg_reg[16]  ( .D(N17), .CLK(clk), .RSTB(n11), .Q(P[16]) );
  DFFARX1 \P_reg_reg[15]  ( .D(N16), .CLK(clk), .RSTB(n11), .Q(P[15]) );
  DFFARX1 \P_reg_reg[14]  ( .D(N15), .CLK(clk), .RSTB(n11), .Q(P[14]) );
  DFFARX1 \P_reg_reg[13]  ( .D(N14), .CLK(clk), .RSTB(n11), .Q(P[13]) );
  DFFARX1 \P_reg_reg[12]  ( .D(N13), .CLK(clk), .RSTB(n11), .Q(P[12]) );
  DFFARX1 \P_reg_reg[11]  ( .D(N12), .CLK(clk), .RSTB(n11), .Q(P[11]) );
  DFFARX1 \P_reg_reg[10]  ( .D(N11), .CLK(clk), .RSTB(n11), .Q(P[10]) );
  DFFARX1 \P_reg_reg[9]  ( .D(N10), .CLK(clk), .RSTB(n11), .Q(P[9]) );
  DFFARX1 \P_reg_reg[8]  ( .D(N9), .CLK(clk), .RSTB(n11), .Q(P[8]) );
  DFFARX1 \P_reg_reg[7]  ( .D(N8), .CLK(clk), .RSTB(n10), .Q(P[7]) );
  DFFARX1 \P_reg_reg[6]  ( .D(N7), .CLK(clk), .RSTB(n10), .Q(P[6]) );
  DFFARX1 \P_reg_reg[5]  ( .D(N6), .CLK(clk), .RSTB(n10), .Q(P[5]) );
  DFFARX1 \P_reg_reg[4]  ( .D(N5), .CLK(clk), .RSTB(n10), .Q(P[4]) );
  DFFARX1 \P_reg_reg[3]  ( .D(N4), .CLK(clk), .RSTB(n10), .Q(P[3]) );
  DFFARX1 \P_reg_reg[2]  ( .D(N3), .CLK(clk), .RSTB(n10), .Q(P[2]) );
  DFFARX1 \P_reg_reg[1]  ( .D(N2), .CLK(clk), .RSTB(n10), .Q(P[1]) );
  DFFARX1 \P_reg_reg[0]  ( .D(N1), .CLK(clk), .RSTB(n10), .Q(P[0]) );
  DFFARX1 \B_reg_reg[31]  ( .D(B[31]), .CLK(clk), .RSTB(n10), .Q(B_reg[31]) );
  DFFARX1 \B_reg_reg[30]  ( .D(B[30]), .CLK(clk), .RSTB(n10), .Q(B_reg[30]) );
  DFFARX1 \B_reg_reg[29]  ( .D(B[29]), .CLK(clk), .RSTB(n9), .Q(B_reg[29]) );
  DFFARX1 \B_reg_reg[28]  ( .D(B[28]), .CLK(clk), .RSTB(n9), .Q(B_reg[28]) );
  DFFARX1 \B_reg_reg[27]  ( .D(B[27]), .CLK(clk), .RSTB(n9), .Q(B_reg[27]) );
  DFFARX1 \B_reg_reg[26]  ( .D(B[26]), .CLK(clk), .RSTB(n9), .Q(B_reg[26]) );
  DFFARX1 \B_reg_reg[25]  ( .D(B[25]), .CLK(clk), .RSTB(n9), .Q(B_reg[25]) );
  DFFARX1 \B_reg_reg[24]  ( .D(B[24]), .CLK(clk), .RSTB(n9), .Q(B_reg[24]) );
  DFFARX1 \B_reg_reg[23]  ( .D(B[23]), .CLK(clk), .RSTB(n9), .Q(B_reg[23]) );
  DFFARX1 \B_reg_reg[22]  ( .D(B[22]), .CLK(clk), .RSTB(n9), .Q(B_reg[22]) );
  DFFARX1 \B_reg_reg[21]  ( .D(B[21]), .CLK(clk), .RSTB(n9), .Q(B_reg[21]) );
  DFFARX1 \B_reg_reg[20]  ( .D(B[20]), .CLK(clk), .RSTB(n9), .Q(B_reg[20]) );
  DFFARX1 \B_reg_reg[19]  ( .D(B[19]), .CLK(clk), .RSTB(n8), .Q(B_reg[19]) );
  DFFARX1 \B_reg_reg[18]  ( .D(B[18]), .CLK(clk), .RSTB(n8), .Q(B_reg[18]) );
  DFFARX1 \B_reg_reg[17]  ( .D(B[17]), .CLK(clk), .RSTB(n8), .Q(B_reg[17]) );
  DFFARX1 \B_reg_reg[16]  ( .D(B[16]), .CLK(clk), .RSTB(n8), .Q(B_reg[16]) );
  DFFARX1 \B_reg_reg[15]  ( .D(B[15]), .CLK(clk), .RSTB(n8), .Q(B_reg[15]) );
  DFFARX1 \B_reg_reg[14]  ( .D(B[14]), .CLK(clk), .RSTB(n8), .Q(B_reg[14]) );
  DFFARX1 \B_reg_reg[13]  ( .D(B[13]), .CLK(clk), .RSTB(n8), .Q(B_reg[13]) );
  DFFARX1 \B_reg_reg[12]  ( .D(B[12]), .CLK(clk), .RSTB(n8), .Q(B_reg[12]) );
  DFFARX1 \B_reg_reg[11]  ( .D(B[11]), .CLK(clk), .RSTB(n8), .Q(B_reg[11]) );
  DFFARX1 \B_reg_reg[10]  ( .D(B[10]), .CLK(clk), .RSTB(n8), .Q(B_reg[10]) );
  DFFARX1 \B_reg_reg[9]  ( .D(B[9]), .CLK(clk), .RSTB(n7), .Q(B_reg[9]) );
  DFFARX1 \B_reg_reg[8]  ( .D(B[8]), .CLK(clk), .RSTB(n7), .Q(B_reg[8]) );
  DFFARX1 \B_reg_reg[7]  ( .D(B[7]), .CLK(clk), .RSTB(n7), .Q(B_reg[7]) );
  DFFARX1 \B_reg_reg[6]  ( .D(B[6]), .CLK(clk), .RSTB(n7), .Q(B_reg[6]) );
  DFFARX1 \B_reg_reg[5]  ( .D(B[5]), .CLK(clk), .RSTB(n7), .Q(B_reg[5]) );
  DFFARX1 \B_reg_reg[4]  ( .D(B[4]), .CLK(clk), .RSTB(n7), .Q(B_reg[4]) );
  DFFARX1 \B_reg_reg[3]  ( .D(B[3]), .CLK(clk), .RSTB(n7), .Q(B_reg[3]) );
  DFFARX1 \B_reg_reg[2]  ( .D(B[2]), .CLK(clk), .RSTB(n7), .Q(B_reg[2]) );
  DFFARX1 \B_reg_reg[1]  ( .D(B[1]), .CLK(clk), .RSTB(n7), .Q(B_reg[1]) );
  DFFARX1 \B_reg_reg[0]  ( .D(B[0]), .CLK(clk), .RSTB(n7), .Q(B_reg[0]) );
  VerilogMultiplier_DW02_mult_0 mult_21 ( .A(A_reg), .B(B_reg), .TC(1'b1), 
        .PRODUCT({N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4, N3, N2, N1}) );
  NBUFFX2 U4 ( .INP(n2), .Z(n7) );
  NBUFFX2 U5 ( .INP(n2), .Z(n8) );
  NBUFFX2 U6 ( .INP(n2), .Z(n9) );
  NBUFFX2 U7 ( .INP(n3), .Z(n10) );
  NBUFFX2 U8 ( .INP(n3), .Z(n11) );
  NBUFFX2 U9 ( .INP(n3), .Z(n12) );
  NBUFFX2 U10 ( .INP(n4), .Z(n13) );
  NBUFFX2 U11 ( .INP(n4), .Z(n14) );
  NBUFFX2 U12 ( .INP(n4), .Z(n15) );
  NBUFFX2 U13 ( .INP(n5), .Z(n16) );
  NBUFFX2 U14 ( .INP(n5), .Z(n17) );
  NBUFFX2 U15 ( .INP(n5), .Z(n18) );
  NBUFFX2 U16 ( .INP(n6), .Z(n19) );
  NBUFFX2 U17 ( .INP(n20), .Z(n6) );
  NBUFFX2 U18 ( .INP(n20), .Z(n2) );
  NBUFFX2 U19 ( .INP(n20), .Z(n3) );
  NBUFFX2 U20 ( .INP(n20), .Z(n4) );
  NBUFFX2 U21 ( .INP(n20), .Z(n5) );
  INVX0 U22 ( .INP(rst), .ZN(n20) );
endmodule

