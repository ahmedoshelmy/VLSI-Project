
module WallaceTreeMultiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160;
  wire   [63:1] carry;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  FA_X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  FA_X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  FA_X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  FA_X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  FA_X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FA_X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  FA_X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  FA_X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FA_X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_9 ( .A(B[9]), .B(A[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n58), .CO(carry[3]), .S(SUM[2]) );
  XOR2_X1 U1 ( .A(A[63]), .B(B[63]), .Z(n1) );
  XOR2_X1 U2 ( .A(carry[63]), .B(n1), .Z(SUM[63]) );
  XOR2_X1 U3 ( .A(A[30]), .B(B[30]), .Z(n2) );
  XOR2_X1 U4 ( .A(carry[30]), .B(n2), .Z(SUM[30]) );
  NAND2_X1 U5 ( .A1(carry[30]), .A2(A[30]), .ZN(n3) );
  NAND2_X1 U6 ( .A1(carry[30]), .A2(B[30]), .ZN(n4) );
  NAND2_X1 U7 ( .A1(A[30]), .A2(B[30]), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n3), .A2(n4), .A3(n5), .ZN(carry[31]) );
  XOR2_X1 U9 ( .A(B[31]), .B(A[31]), .Z(n6) );
  XOR2_X1 U10 ( .A(carry[31]), .B(n6), .Z(SUM[31]) );
  NAND2_X1 U11 ( .A1(carry[31]), .A2(B[31]), .ZN(n7) );
  NAND2_X1 U12 ( .A1(carry[31]), .A2(A[31]), .ZN(n8) );
  NAND2_X1 U13 ( .A1(B[31]), .A2(A[31]), .ZN(n9) );
  NAND3_X1 U14 ( .A1(n7), .A2(n8), .A3(n9), .ZN(carry[32]) );
  XOR2_X1 U15 ( .A(B[17]), .B(A[17]), .Z(n10) );
  XOR2_X1 U16 ( .A(carry[17]), .B(n10), .Z(SUM[17]) );
  NAND2_X1 U17 ( .A1(carry[17]), .A2(B[17]), .ZN(n11) );
  NAND2_X1 U18 ( .A1(carry[17]), .A2(A[17]), .ZN(n12) );
  NAND2_X1 U19 ( .A1(B[17]), .A2(A[17]), .ZN(n13) );
  NAND3_X1 U20 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[18]) );
  XOR2_X1 U21 ( .A(A[53]), .B(B[53]), .Z(n14) );
  XOR2_X1 U22 ( .A(carry[53]), .B(n14), .Z(SUM[53]) );
  NAND2_X1 U23 ( .A1(carry[53]), .A2(A[53]), .ZN(n15) );
  NAND2_X1 U24 ( .A1(carry[53]), .A2(B[53]), .ZN(n16) );
  NAND2_X1 U25 ( .A1(A[53]), .A2(B[53]), .ZN(n17) );
  NAND3_X1 U26 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[54]) );
  XOR2_X1 U27 ( .A(A[47]), .B(B[47]), .Z(n18) );
  XOR2_X1 U28 ( .A(carry[47]), .B(n18), .Z(SUM[47]) );
  NAND2_X1 U29 ( .A1(carry[47]), .A2(A[47]), .ZN(n19) );
  NAND2_X1 U30 ( .A1(carry[47]), .A2(B[47]), .ZN(n20) );
  NAND2_X1 U31 ( .A1(A[47]), .A2(B[47]), .ZN(n21) );
  NAND3_X1 U32 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[48]) );
  XOR2_X1 U33 ( .A(B[56]), .B(A[56]), .Z(n22) );
  XOR2_X1 U34 ( .A(carry[56]), .B(n22), .Z(SUM[56]) );
  NAND2_X1 U35 ( .A1(carry[56]), .A2(B[56]), .ZN(n23) );
  NAND2_X1 U36 ( .A1(carry[56]), .A2(A[56]), .ZN(n24) );
  NAND2_X1 U37 ( .A1(B[56]), .A2(A[56]), .ZN(n25) );
  NAND3_X1 U38 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[57]) );
  XOR2_X1 U39 ( .A(A[32]), .B(B[32]), .Z(n26) );
  XOR2_X1 U40 ( .A(carry[32]), .B(n26), .Z(SUM[32]) );
  NAND2_X1 U41 ( .A1(carry[32]), .A2(A[32]), .ZN(n27) );
  NAND2_X1 U42 ( .A1(carry[32]), .A2(B[32]), .ZN(n28) );
  NAND2_X1 U43 ( .A1(A[32]), .A2(B[32]), .ZN(n29) );
  NAND3_X1 U44 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[33]) );
  XOR2_X1 U45 ( .A(B[18]), .B(A[18]), .Z(n30) );
  XOR2_X1 U46 ( .A(carry[18]), .B(n30), .Z(SUM[18]) );
  NAND2_X1 U47 ( .A1(carry[18]), .A2(B[18]), .ZN(n31) );
  NAND2_X1 U48 ( .A1(carry[18]), .A2(A[18]), .ZN(n32) );
  NAND2_X1 U49 ( .A1(B[18]), .A2(A[18]), .ZN(n33) );
  NAND3_X1 U50 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[19]) );
  XOR2_X1 U51 ( .A(B[12]), .B(A[12]), .Z(n34) );
  XOR2_X1 U52 ( .A(carry[12]), .B(n34), .Z(SUM[12]) );
  NAND2_X1 U53 ( .A1(carry[12]), .A2(B[12]), .ZN(n35) );
  NAND2_X1 U54 ( .A1(carry[12]), .A2(A[12]), .ZN(n36) );
  NAND2_X1 U55 ( .A1(B[12]), .A2(A[12]), .ZN(n37) );
  NAND3_X1 U56 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[13]) );
  XOR2_X1 U57 ( .A(A[57]), .B(B[57]), .Z(n38) );
  XOR2_X1 U58 ( .A(carry[57]), .B(n38), .Z(SUM[57]) );
  NAND2_X1 U59 ( .A1(carry[57]), .A2(A[57]), .ZN(n39) );
  NAND2_X1 U60 ( .A1(carry[57]), .A2(B[57]), .ZN(n40) );
  NAND2_X1 U61 ( .A1(A[57]), .A2(B[57]), .ZN(n41) );
  NAND3_X1 U62 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[58]) );
  XOR2_X1 U63 ( .A(B[13]), .B(A[13]), .Z(n42) );
  XOR2_X1 U64 ( .A(carry[13]), .B(n42), .Z(SUM[13]) );
  NAND2_X1 U65 ( .A1(carry[13]), .A2(B[13]), .ZN(n43) );
  NAND2_X1 U66 ( .A1(carry[13]), .A2(A[13]), .ZN(n44) );
  NAND2_X1 U67 ( .A1(B[13]), .A2(A[13]), .ZN(n45) );
  NAND3_X1 U68 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[14]) );
  XOR2_X1 U69 ( .A(A[24]), .B(B[24]), .Z(n46) );
  XOR2_X1 U70 ( .A(carry[24]), .B(n46), .Z(SUM[24]) );
  NAND2_X1 U71 ( .A1(carry[24]), .A2(A[24]), .ZN(n47) );
  NAND2_X1 U72 ( .A1(carry[24]), .A2(B[24]), .ZN(n48) );
  NAND2_X1 U73 ( .A1(A[24]), .A2(B[24]), .ZN(n49) );
  NAND3_X1 U74 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[25]) );
  XOR2_X1 U75 ( .A(B[27]), .B(A[27]), .Z(n50) );
  XOR2_X1 U76 ( .A(carry[27]), .B(n50), .Z(SUM[27]) );
  NAND2_X1 U77 ( .A1(carry[27]), .A2(B[27]), .ZN(n51) );
  NAND2_X1 U78 ( .A1(carry[27]), .A2(A[27]), .ZN(n52) );
  NAND2_X1 U79 ( .A1(B[27]), .A2(A[27]), .ZN(n53) );
  NAND3_X1 U80 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[28]) );
  XOR2_X1 U81 ( .A(B[14]), .B(A[14]), .Z(n54) );
  XOR2_X1 U82 ( .A(carry[14]), .B(n54), .Z(SUM[14]) );
  NAND2_X1 U83 ( .A1(carry[14]), .A2(B[14]), .ZN(n55) );
  NAND2_X1 U84 ( .A1(carry[14]), .A2(A[14]), .ZN(n56) );
  NAND2_X1 U85 ( .A1(B[14]), .A2(A[14]), .ZN(n57) );
  NAND3_X1 U86 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[15]) );
  AND2_X1 U87 ( .A1(B[1]), .A2(A[1]), .ZN(n58) );
  XOR2_X1 U88 ( .A(B[28]), .B(A[28]), .Z(n59) );
  XOR2_X1 U89 ( .A(carry[28]), .B(n59), .Z(SUM[28]) );
  NAND2_X1 U90 ( .A1(carry[28]), .A2(B[28]), .ZN(n60) );
  NAND2_X1 U91 ( .A1(carry[28]), .A2(A[28]), .ZN(n61) );
  NAND2_X1 U92 ( .A1(B[28]), .A2(A[28]), .ZN(n62) );
  NAND3_X1 U93 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[29]) );
  XOR2_X1 U94 ( .A(A[45]), .B(B[45]), .Z(n63) );
  XOR2_X1 U95 ( .A(carry[45]), .B(n63), .Z(SUM[45]) );
  NAND2_X1 U96 ( .A1(carry[45]), .A2(A[45]), .ZN(n64) );
  NAND2_X1 U97 ( .A1(carry[45]), .A2(B[45]), .ZN(n65) );
  NAND2_X1 U98 ( .A1(A[45]), .A2(B[45]), .ZN(n66) );
  NAND3_X1 U99 ( .A1(n64), .A2(n65), .A3(n66), .ZN(carry[46]) );
  XOR2_X1 U100 ( .A(A[33]), .B(B[33]), .Z(n67) );
  XOR2_X1 U101 ( .A(carry[33]), .B(n67), .Z(SUM[33]) );
  NAND2_X1 U102 ( .A1(carry[33]), .A2(A[33]), .ZN(n68) );
  NAND2_X1 U103 ( .A1(carry[33]), .A2(B[33]), .ZN(n69) );
  NAND2_X1 U104 ( .A1(A[33]), .A2(B[33]), .ZN(n70) );
  NAND3_X1 U105 ( .A1(n68), .A2(n69), .A3(n70), .ZN(carry[34]) );
  XOR2_X1 U106 ( .A(B[15]), .B(A[15]), .Z(n71) );
  XOR2_X1 U107 ( .A(carry[15]), .B(n71), .Z(SUM[15]) );
  NAND2_X1 U108 ( .A1(carry[15]), .A2(B[15]), .ZN(n72) );
  NAND2_X1 U109 ( .A1(carry[15]), .A2(A[15]), .ZN(n73) );
  NAND2_X1 U110 ( .A1(B[15]), .A2(A[15]), .ZN(n74) );
  NAND3_X1 U111 ( .A1(n72), .A2(n73), .A3(n74), .ZN(carry[16]) );
  XOR2_X1 U112 ( .A(B[37]), .B(A[37]), .Z(n75) );
  XOR2_X1 U113 ( .A(n80), .B(n75), .Z(SUM[37]) );
  NAND2_X1 U114 ( .A1(n79), .A2(B[37]), .ZN(n76) );
  NAND2_X1 U115 ( .A1(carry[37]), .A2(A[37]), .ZN(n77) );
  NAND2_X1 U116 ( .A1(B[37]), .A2(A[37]), .ZN(n78) );
  NAND3_X1 U117 ( .A1(n76), .A2(n77), .A3(n78), .ZN(carry[38]) );
  NAND3_X1 U118 ( .A1(n90), .A2(n91), .A3(n92), .ZN(n79) );
  NAND3_X1 U119 ( .A1(n90), .A2(n91), .A3(n92), .ZN(n80) );
  XOR2_X1 U120 ( .A(A[8]), .B(B[8]), .Z(n81) );
  XOR2_X1 U121 ( .A(carry[8]), .B(n81), .Z(SUM[8]) );
  NAND2_X1 U122 ( .A1(carry[8]), .A2(A[8]), .ZN(n82) );
  NAND2_X1 U123 ( .A1(carry[8]), .A2(B[8]), .ZN(n83) );
  NAND2_X1 U124 ( .A1(A[8]), .A2(B[8]), .ZN(n84) );
  NAND3_X1 U125 ( .A1(n82), .A2(n84), .A3(n83), .ZN(carry[9]) );
  XOR2_X1 U126 ( .A(B[22]), .B(A[22]), .Z(n85) );
  XOR2_X1 U127 ( .A(carry[22]), .B(n85), .Z(SUM[22]) );
  NAND2_X1 U128 ( .A1(carry[22]), .A2(B[22]), .ZN(n86) );
  NAND2_X1 U129 ( .A1(carry[22]), .A2(A[22]), .ZN(n87) );
  NAND2_X1 U130 ( .A1(B[22]), .A2(A[22]), .ZN(n88) );
  NAND3_X1 U131 ( .A1(n86), .A2(n87), .A3(n88), .ZN(carry[23]) );
  XOR2_X1 U132 ( .A(B[36]), .B(A[36]), .Z(n89) );
  XOR2_X1 U133 ( .A(carry[36]), .B(n89), .Z(SUM[36]) );
  NAND2_X1 U134 ( .A1(carry[36]), .A2(B[36]), .ZN(n90) );
  NAND2_X1 U135 ( .A1(carry[36]), .A2(A[36]), .ZN(n91) );
  NAND2_X1 U136 ( .A1(B[36]), .A2(A[36]), .ZN(n92) );
  NAND3_X1 U137 ( .A1(n90), .A2(n91), .A3(n92), .ZN(carry[37]) );
  XOR2_X1 U138 ( .A(A[60]), .B(B[60]), .Z(n93) );
  XOR2_X1 U139 ( .A(carry[60]), .B(n93), .Z(SUM[60]) );
  NAND2_X1 U140 ( .A1(carry[60]), .A2(A[60]), .ZN(n94) );
  NAND2_X1 U141 ( .A1(carry[60]), .A2(B[60]), .ZN(n95) );
  NAND2_X1 U142 ( .A1(A[60]), .A2(B[60]), .ZN(n96) );
  NAND3_X1 U143 ( .A1(n94), .A2(n95), .A3(n96), .ZN(carry[61]) );
  XOR2_X1 U144 ( .A(A[48]), .B(B[48]), .Z(n97) );
  XOR2_X1 U145 ( .A(carry[48]), .B(n97), .Z(SUM[48]) );
  NAND2_X1 U146 ( .A1(carry[48]), .A2(A[48]), .ZN(n98) );
  NAND2_X1 U147 ( .A1(carry[48]), .A2(B[48]), .ZN(n99) );
  NAND2_X1 U148 ( .A1(A[48]), .A2(B[48]), .ZN(n100) );
  NAND3_X1 U149 ( .A1(n98), .A2(n99), .A3(n100), .ZN(carry[49]) );
  XOR2_X1 U150 ( .A(B[35]), .B(A[35]), .Z(n101) );
  XOR2_X1 U151 ( .A(carry[35]), .B(n101), .Z(SUM[35]) );
  NAND2_X1 U152 ( .A1(carry[35]), .A2(B[35]), .ZN(n102) );
  NAND2_X1 U153 ( .A1(carry[35]), .A2(A[35]), .ZN(n103) );
  NAND2_X1 U154 ( .A1(B[35]), .A2(A[35]), .ZN(n104) );
  NAND3_X1 U155 ( .A1(n102), .A2(n103), .A3(n104), .ZN(carry[36]) );
  XOR2_X1 U156 ( .A(B[21]), .B(A[21]), .Z(n105) );
  XOR2_X1 U157 ( .A(carry[21]), .B(n105), .Z(SUM[21]) );
  NAND2_X1 U158 ( .A1(carry[21]), .A2(B[21]), .ZN(n106) );
  NAND2_X1 U159 ( .A1(carry[21]), .A2(A[21]), .ZN(n107) );
  NAND2_X1 U160 ( .A1(B[21]), .A2(A[21]), .ZN(n108) );
  NAND3_X1 U161 ( .A1(n106), .A2(n107), .A3(n108), .ZN(carry[22]) );
  XOR2_X1 U162 ( .A(B[40]), .B(A[40]), .Z(n109) );
  XOR2_X1 U163 ( .A(carry[40]), .B(n109), .Z(SUM[40]) );
  NAND2_X1 U164 ( .A1(carry[40]), .A2(B[40]), .ZN(n110) );
  NAND2_X1 U165 ( .A1(carry[40]), .A2(A[40]), .ZN(n111) );
  NAND2_X1 U166 ( .A1(B[40]), .A2(A[40]), .ZN(n112) );
  NAND3_X1 U167 ( .A1(n110), .A2(n111), .A3(n112), .ZN(carry[41]) );
  XOR2_X1 U168 ( .A(B[19]), .B(A[19]), .Z(n113) );
  XOR2_X1 U169 ( .A(carry[19]), .B(n113), .Z(SUM[19]) );
  NAND2_X1 U170 ( .A1(carry[19]), .A2(B[19]), .ZN(n114) );
  NAND2_X1 U171 ( .A1(carry[19]), .A2(A[19]), .ZN(n115) );
  NAND2_X1 U172 ( .A1(B[19]), .A2(A[19]), .ZN(n116) );
  NAND3_X1 U173 ( .A1(n114), .A2(n115), .A3(n116), .ZN(carry[20]) );
  XOR2_X1 U174 ( .A(A[44]), .B(B[44]), .Z(n117) );
  XOR2_X1 U175 ( .A(carry[44]), .B(n117), .Z(SUM[44]) );
  NAND2_X1 U176 ( .A1(carry[44]), .A2(A[44]), .ZN(n118) );
  NAND2_X1 U177 ( .A1(carry[44]), .A2(B[44]), .ZN(n119) );
  NAND2_X1 U178 ( .A1(A[44]), .A2(B[44]), .ZN(n120) );
  NAND3_X1 U179 ( .A1(n118), .A2(n119), .A3(n120), .ZN(carry[45]) );
  XOR2_X1 U180 ( .A(A[59]), .B(B[59]), .Z(n121) );
  XOR2_X1 U181 ( .A(carry[59]), .B(n121), .Z(SUM[59]) );
  NAND2_X1 U182 ( .A1(carry[59]), .A2(A[59]), .ZN(n122) );
  NAND2_X1 U183 ( .A1(carry[59]), .A2(B[59]), .ZN(n123) );
  NAND2_X1 U184 ( .A1(A[59]), .A2(B[59]), .ZN(n124) );
  NAND3_X1 U185 ( .A1(n122), .A2(n123), .A3(n124), .ZN(carry[60]) );
  XOR2_X1 U186 ( .A(A[42]), .B(B[42]), .Z(n125) );
  XOR2_X1 U187 ( .A(carry[42]), .B(n125), .Z(SUM[42]) );
  NAND2_X1 U188 ( .A1(carry[42]), .A2(A[42]), .ZN(n126) );
  NAND2_X1 U189 ( .A1(carry[42]), .A2(B[42]), .ZN(n127) );
  NAND2_X1 U190 ( .A1(A[42]), .A2(B[42]), .ZN(n128) );
  NAND3_X1 U191 ( .A1(n126), .A2(n127), .A3(n128), .ZN(carry[43]) );
  XOR2_X1 U192 ( .A(A[62]), .B(B[62]), .Z(n129) );
  XOR2_X1 U193 ( .A(carry[62]), .B(n129), .Z(SUM[62]) );
  NAND2_X1 U194 ( .A1(carry[62]), .A2(A[62]), .ZN(n130) );
  NAND2_X1 U195 ( .A1(carry[62]), .A2(B[62]), .ZN(n131) );
  NAND2_X1 U196 ( .A1(A[62]), .A2(B[62]), .ZN(n132) );
  NAND3_X1 U197 ( .A1(n130), .A2(n131), .A3(n132), .ZN(carry[63]) );
  XOR2_X1 U198 ( .A(A[51]), .B(B[51]), .Z(n133) );
  XOR2_X1 U199 ( .A(carry[51]), .B(n133), .Z(SUM[51]) );
  NAND2_X1 U200 ( .A1(carry[51]), .A2(A[51]), .ZN(n134) );
  NAND2_X1 U201 ( .A1(carry[51]), .A2(B[51]), .ZN(n135) );
  NAND2_X1 U202 ( .A1(A[51]), .A2(B[51]), .ZN(n136) );
  NAND3_X1 U203 ( .A1(n134), .A2(n135), .A3(n136), .ZN(carry[52]) );
  XOR2_X1 U204 ( .A(B[39]), .B(A[39]), .Z(n137) );
  XOR2_X1 U205 ( .A(carry[39]), .B(n137), .Z(SUM[39]) );
  NAND2_X1 U206 ( .A1(carry[39]), .A2(B[39]), .ZN(n138) );
  NAND2_X1 U207 ( .A1(carry[39]), .A2(A[39]), .ZN(n139) );
  NAND2_X1 U208 ( .A1(B[39]), .A2(A[39]), .ZN(n140) );
  NAND3_X1 U209 ( .A1(n138), .A2(n139), .A3(n140), .ZN(carry[40]) );
  XOR2_X1 U210 ( .A(A[25]), .B(B[25]), .Z(n141) );
  XOR2_X1 U211 ( .A(carry[25]), .B(n141), .Z(SUM[25]) );
  NAND2_X1 U212 ( .A1(carry[25]), .A2(A[25]), .ZN(n142) );
  NAND2_X1 U213 ( .A1(carry[25]), .A2(B[25]), .ZN(n143) );
  NAND2_X1 U214 ( .A1(A[25]), .A2(B[25]), .ZN(n144) );
  NAND3_X1 U215 ( .A1(n142), .A2(n143), .A3(n144), .ZN(carry[26]) );
  XOR2_X1 U216 ( .A(B[10]), .B(A[10]), .Z(n145) );
  XOR2_X1 U217 ( .A(carry[10]), .B(n145), .Z(SUM[10]) );
  NAND2_X1 U218 ( .A1(carry[10]), .A2(B[10]), .ZN(n146) );
  NAND2_X1 U219 ( .A1(carry[10]), .A2(A[10]), .ZN(n147) );
  NAND2_X1 U220 ( .A1(B[10]), .A2(A[10]), .ZN(n148) );
  NAND3_X1 U221 ( .A1(n146), .A2(n147), .A3(n148), .ZN(carry[11]) );
  XOR2_X1 U222 ( .A(A[50]), .B(B[50]), .Z(n149) );
  XOR2_X1 U223 ( .A(carry[50]), .B(n149), .Z(SUM[50]) );
  NAND2_X1 U224 ( .A1(carry[50]), .A2(A[50]), .ZN(n150) );
  NAND2_X1 U225 ( .A1(carry[50]), .A2(B[50]), .ZN(n151) );
  NAND2_X1 U226 ( .A1(A[50]), .A2(B[50]), .ZN(n152) );
  NAND3_X1 U227 ( .A1(n151), .A2(n150), .A3(n152), .ZN(carry[51]) );
  XOR2_X1 U228 ( .A(A[54]), .B(B[54]), .Z(n153) );
  XOR2_X1 U229 ( .A(carry[54]), .B(n153), .Z(SUM[54]) );
  NAND2_X1 U230 ( .A1(carry[54]), .A2(A[54]), .ZN(n154) );
  NAND2_X1 U231 ( .A1(carry[54]), .A2(B[54]), .ZN(n155) );
  NAND2_X1 U232 ( .A1(A[54]), .A2(B[54]), .ZN(n156) );
  NAND3_X1 U233 ( .A1(n154), .A2(n155), .A3(n156), .ZN(carry[55]) );
  XOR2_X1 U234 ( .A(A[58]), .B(B[58]), .Z(n157) );
  XOR2_X1 U235 ( .A(carry[58]), .B(n157), .Z(SUM[58]) );
  NAND2_X1 U236 ( .A1(carry[58]), .A2(A[58]), .ZN(n158) );
  NAND2_X1 U237 ( .A1(carry[58]), .A2(B[58]), .ZN(n159) );
  NAND2_X1 U238 ( .A1(A[58]), .A2(B[58]), .ZN(n160) );
  NAND3_X1 U239 ( .A1(n158), .A2(n159), .A3(n160), .ZN(carry[59]) );
  XOR2_X1 U240 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
endmodule


module WallaceTreeMultiplier ( A, B, out, clk, rst );
  input [31:0] A;
  input [31:0] B;
  output [63:0] out;
  input clk, rst;
  wire   N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, \p[7][63] , \p[7][37] ,
         \p[7][36] , \p[7][35] , \p[7][34] , \p[7][33] , \p[7][32] ,
         \p[7][31] , \p[7][30] , \p[7][29] , \p[7][28] , \p[7][27] ,
         \p[7][26] , \p[7][25] , \p[7][24] , \p[7][23] , \p[7][22] ,
         \p[7][21] , \p[7][20] , \p[7][19] , \p[7][18] , \p[7][17] ,
         \p[7][16] , \p[7][15] , \p[7][14] , \p[7][13] , \p[7][12] ,
         \p[7][11] , \p[7][10] , \p[7][9] , \p[7][8] , \p[7][7] , \p[6][63] ,
         \p[6][36] , \p[6][35] , \p[6][34] , \p[6][33] , \p[6][32] ,
         \p[6][31] , \p[6][30] , \p[6][29] , \p[6][28] , \p[6][27] ,
         \p[6][26] , \p[6][25] , \p[6][24] , \p[6][23] , \p[6][22] ,
         \p[6][21] , \p[6][20] , \p[6][19] , \p[6][18] , \p[6][17] ,
         \p[6][16] , \p[6][15] , \p[6][14] , \p[6][13] , \p[6][12] ,
         \p[6][11] , \p[6][10] , \p[6][9] , \p[6][8] , \p[6][7] , \p[6][6] ,
         \p[5][63] , \p[5][35] , \p[5][34] , \p[5][33] , \p[5][32] ,
         \p[5][31] , \p[5][30] , \p[5][29] , \p[5][28] , \p[5][27] ,
         \p[5][26] , \p[5][25] , \p[5][24] , \p[5][23] , \p[5][22] ,
         \p[5][21] , \p[5][20] , \p[5][19] , \p[5][18] , \p[5][17] ,
         \p[5][16] , \p[5][15] , \p[5][14] , \p[5][13] , \p[5][12] ,
         \p[5][11] , \p[5][10] , \p[5][9] , \p[5][8] , \p[5][7] , \p[5][6] ,
         \p[5][5] , \p[4][63] , \p[4][34] , \p[4][33] , \p[4][32] , \p[4][31] ,
         \p[4][30] , \p[4][29] , \p[4][28] , \p[4][27] , \p[4][26] ,
         \p[4][25] , \p[4][24] , \p[4][23] , \p[4][22] , \p[4][21] ,
         \p[4][20] , \p[4][19] , \p[4][18] , \p[4][17] , \p[4][16] ,
         \p[4][15] , \p[4][14] , \p[4][13] , \p[4][12] , \p[4][11] ,
         \p[4][10] , \p[4][9] , \p[4][8] , \p[4][7] , \p[4][6] , \p[4][5] ,
         \p[4][4] , \p[3][63] , \p[3][33] , \p[3][32] , \p[3][31] , \p[3][30] ,
         \p[3][29] , \p[3][28] , \p[3][27] , \p[3][26] , \p[3][25] ,
         \p[3][24] , \p[3][23] , \p[3][22] , \p[3][21] , \p[3][20] ,
         \p[3][19] , \p[3][18] , \p[3][17] , \p[3][16] , \p[3][15] ,
         \p[3][14] , \p[3][13] , \p[3][12] , \p[3][11] , \p[3][10] , \p[3][9] ,
         \p[3][8] , \p[3][7] , \p[3][6] , \p[3][5] , \p[3][4] , \p[3][3] ,
         \p[2][63] , \p[2][32] , \p[2][31] , \p[2][30] , \p[2][29] ,
         \p[2][28] , \p[2][27] , \p[2][26] , \p[2][25] , \p[2][24] ,
         \p[2][23] , \p[2][22] , \p[2][21] , \p[2][20] , \p[2][19] ,
         \p[2][18] , \p[2][17] , \p[2][16] , \p[2][15] , \p[2][14] ,
         \p[2][13] , \p[2][12] , \p[2][11] , \p[2][10] , \p[2][9] , \p[2][8] ,
         \p[2][7] , \p[2][6] , \p[2][5] , \p[2][4] , \p[2][3] , \p[2][2] ,
         \p[1][63] , \p[1][31] , \p[1][30] , \p[1][29] , \p[1][28] ,
         \p[1][27] , \p[1][26] , \p[1][25] , \p[1][24] , \p[1][23] ,
         \p[1][22] , \p[1][21] , \p[1][20] , \p[1][19] , \p[1][18] ,
         \p[1][17] , \p[1][16] , \p[1][15] , \p[1][14] , \p[1][13] ,
         \p[1][12] , \p[1][11] , \p[1][10] , \p[1][9] , \p[1][8] , \p[1][7] ,
         \p[1][6] , \p[1][5] , \p[1][4] , \p[1][3] , \p[1][2] , \p[1][1] ,
         \p[0][63] , \p[0][30] , \p[0][29] , \p[0][28] , \p[0][27] ,
         \p[0][26] , \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] ,
         \p[0][21] , \p[0][20] , \p[0][19] , \p[0][18] , \p[0][17] ,
         \p[0][16] , \p[0][15] , \p[0][14] , \p[0][13] , \p[0][12] ,
         \p[0][11] , \p[0][10] , \p[0][9] , \p[0][8] , \p[0][7] , \p[0][6] ,
         \p[0][5] , \p[0][4] , \p[0][3] , \p[0][2] , \p[0][1] , \p[0][0] ,
         \p[63][63] , \p[62][63] , \p[61][63] , \p[60][63] , \p[59][63] ,
         \p[58][63] , \p[57][63] , \p[56][63] , \p[55][63] , \p[54][63] ,
         \p[53][63] , \p[52][63] , \p[51][63] , \p[50][63] , \p[49][63] ,
         \p[48][63] , \p[47][63] , \p[46][63] , \p[45][63] , \p[44][63] ,
         \p[43][63] , \p[42][63] , \p[41][63] , \p[40][63] , \p[39][63] ,
         \p[38][63] , \p[37][63] , \p[36][63] , \p[35][63] , \p[34][63] ,
         \p[33][63] , \p[32][63] , \p[30][63] , \p[30][60] , \p[30][59] ,
         \p[30][58] , \p[30][57] , \p[30][56] , \p[30][55] , \p[30][54] ,
         \p[30][53] , \p[30][52] , \p[30][51] , \p[30][50] , \p[30][49] ,
         \p[30][48] , \p[30][47] , \p[30][46] , \p[30][45] , \p[30][44] ,
         \p[30][43] , \p[30][42] , \p[30][41] , \p[30][40] , \p[30][39] ,
         \p[30][38] , \p[30][37] , \p[30][36] , \p[30][35] , \p[30][34] ,
         \p[30][33] , \p[30][32] , \p[30][31] , \p[30][30] , \p[29][63] ,
         \p[29][59] , \p[29][58] , \p[29][57] , \p[29][56] , \p[29][55] ,
         \p[29][54] , \p[29][53] , \p[29][52] , \p[29][51] , \p[29][50] ,
         \p[29][49] , \p[29][48] , \p[29][47] , \p[29][46] , \p[29][45] ,
         \p[29][44] , \p[29][43] , \p[29][42] , \p[29][41] , \p[29][40] ,
         \p[29][39] , \p[29][38] , \p[29][37] , \p[29][36] , \p[29][35] ,
         \p[29][34] , \p[29][33] , \p[29][32] , \p[29][31] , \p[29][30] ,
         \p[29][29] , \p[28][63] , \p[28][58] , \p[28][57] , \p[28][56] ,
         \p[28][55] , \p[28][54] , \p[28][53] , \p[28][52] , \p[28][51] ,
         \p[28][50] , \p[28][49] , \p[28][48] , \p[28][47] , \p[28][46] ,
         \p[28][45] , \p[28][44] , \p[28][43] , \p[28][42] , \p[28][41] ,
         \p[28][40] , \p[28][39] , \p[28][38] , \p[28][37] , \p[28][36] ,
         \p[28][35] , \p[28][34] , \p[28][33] , \p[28][32] , \p[28][31] ,
         \p[28][30] , \p[28][29] , \p[28][28] , \p[27][63] , \p[27][57] ,
         \p[27][56] , \p[27][55] , \p[27][54] , \p[27][53] , \p[27][52] ,
         \p[27][51] , \p[27][50] , \p[27][49] , \p[27][48] , \p[27][47] ,
         \p[27][46] , \p[27][45] , \p[27][44] , \p[27][43] , \p[27][42] ,
         \p[27][41] , \p[27][40] , \p[27][39] , \p[27][38] , \p[27][37] ,
         \p[27][36] , \p[27][35] , \p[27][34] , \p[27][33] , \p[27][32] ,
         \p[27][31] , \p[27][30] , \p[27][29] , \p[27][28] , \p[27][27] ,
         \p[26][63] , \p[26][56] , \p[26][55] , \p[26][54] , \p[26][53] ,
         \p[26][52] , \p[26][51] , \p[26][50] , \p[26][49] , \p[26][48] ,
         \p[26][47] , \p[26][46] , \p[26][45] , \p[26][44] , \p[26][43] ,
         \p[26][42] , \p[26][41] , \p[26][40] , \p[26][39] , \p[26][38] ,
         \p[26][37] , \p[26][36] , \p[26][35] , \p[26][34] , \p[26][33] ,
         \p[26][32] , \p[26][31] , \p[26][30] , \p[26][29] , \p[26][28] ,
         \p[26][27] , \p[26][26] , \p[25][63] , \p[25][55] , \p[25][54] ,
         \p[25][53] , \p[25][52] , \p[25][51] , \p[25][50] , \p[25][49] ,
         \p[25][48] , \p[25][47] , \p[25][46] , \p[25][45] , \p[25][44] ,
         \p[25][43] , \p[25][42] , \p[25][41] , \p[25][40] , \p[25][39] ,
         \p[25][38] , \p[25][37] , \p[25][36] , \p[25][35] , \p[25][34] ,
         \p[25][33] , \p[25][32] , \p[25][31] , \p[25][30] , \p[25][29] ,
         \p[25][28] , \p[25][27] , \p[25][26] , \p[25][25] , \p[24][63] ,
         \p[24][54] , \p[24][53] , \p[24][52] , \p[24][51] , \p[24][50] ,
         \p[24][49] , \p[24][48] , \p[24][47] , \p[24][46] , \p[24][45] ,
         \p[24][44] , \p[24][43] , \p[24][42] , \p[24][41] , \p[24][40] ,
         \p[24][39] , \p[24][38] , \p[24][37] , \p[24][36] , \p[24][35] ,
         \p[24][34] , \p[24][33] , \p[24][32] , \p[24][31] , \p[24][30] ,
         \p[24][29] , \p[24][28] , \p[24][27] , \p[24][26] , \p[24][25] ,
         \p[24][24] , \p[23][63] , \p[23][53] , \p[23][52] , \p[23][51] ,
         \p[23][50] , \p[23][49] , \p[23][48] , \p[23][47] , \p[23][46] ,
         \p[23][45] , \p[23][44] , \p[23][43] , \p[23][42] , \p[23][41] ,
         \p[23][40] , \p[23][39] , \p[23][38] , \p[23][37] , \p[23][36] ,
         \p[23][35] , \p[23][34] , \p[23][33] , \p[23][32] , \p[23][31] ,
         \p[23][30] , \p[23][29] , \p[23][28] , \p[23][27] , \p[23][26] ,
         \p[23][25] , \p[23][24] , \p[23][23] , \p[22][63] , \p[22][52] ,
         \p[22][51] , \p[22][50] , \p[22][49] , \p[22][48] , \p[22][47] ,
         \p[22][46] , \p[22][45] , \p[22][44] , \p[22][43] , \p[22][42] ,
         \p[22][41] , \p[22][40] , \p[22][39] , \p[22][38] , \p[22][37] ,
         \p[22][36] , \p[22][35] , \p[22][34] , \p[22][33] , \p[22][32] ,
         \p[22][31] , \p[22][30] , \p[22][29] , \p[22][28] , \p[22][27] ,
         \p[22][26] , \p[22][25] , \p[22][24] , \p[22][23] , \p[22][22] ,
         \p[21][63] , \p[21][51] , \p[21][50] , \p[21][49] , \p[21][48] ,
         \p[21][47] , \p[21][46] , \p[21][45] , \p[21][44] , \p[21][43] ,
         \p[21][42] , \p[21][41] , \p[21][40] , \p[21][39] , \p[21][38] ,
         \p[21][37] , \p[21][36] , \p[21][35] , \p[21][34] , \p[21][33] ,
         \p[21][32] , \p[21][31] , \p[21][30] , \p[21][29] , \p[21][28] ,
         \p[21][27] , \p[21][26] , \p[21][25] , \p[21][24] , \p[21][23] ,
         \p[21][22] , \p[21][21] , \p[20][63] , \p[20][50] , \p[20][49] ,
         \p[20][48] , \p[20][47] , \p[20][46] , \p[20][45] , \p[20][44] ,
         \p[20][43] , \p[20][42] , \p[20][41] , \p[20][40] , \p[20][39] ,
         \p[20][38] , \p[20][37] , \p[20][36] , \p[20][35] , \p[20][34] ,
         \p[20][33] , \p[20][32] , \p[20][31] , \p[20][30] , \p[20][29] ,
         \p[20][28] , \p[20][27] , \p[20][26] , \p[20][25] , \p[20][24] ,
         \p[20][23] , \p[20][22] , \p[20][21] , \p[20][20] , \p[19][63] ,
         \p[19][49] , \p[19][48] , \p[19][47] , \p[19][46] , \p[19][45] ,
         \p[19][44] , \p[19][43] , \p[19][42] , \p[19][41] , \p[19][40] ,
         \p[19][39] , \p[19][38] , \p[19][37] , \p[19][36] , \p[19][35] ,
         \p[19][34] , \p[19][33] , \p[19][32] , \p[19][31] , \p[19][30] ,
         \p[19][29] , \p[19][28] , \p[19][27] , \p[19][26] , \p[19][25] ,
         \p[19][24] , \p[19][23] , \p[19][22] , \p[19][21] , \p[19][20] ,
         \p[19][19] , \p[18][63] , \p[18][48] , \p[18][47] , \p[18][46] ,
         \p[18][45] , \p[18][44] , \p[18][43] , \p[18][42] , \p[18][41] ,
         \p[18][40] , \p[18][39] , \p[18][38] , \p[18][37] , \p[18][36] ,
         \p[18][35] , \p[18][34] , \p[18][33] , \p[18][32] , \p[18][31] ,
         \p[18][30] , \p[18][29] , \p[18][28] , \p[18][27] , \p[18][26] ,
         \p[18][25] , \p[18][24] , \p[18][23] , \p[18][22] , \p[18][21] ,
         \p[18][20] , \p[18][19] , \p[18][18] , \p[17][63] , \p[17][47] ,
         \p[17][46] , \p[17][45] , \p[17][44] , \p[17][43] , \p[17][42] ,
         \p[17][41] , \p[17][40] , \p[17][39] , \p[17][38] , \p[17][37] ,
         \p[17][36] , \p[17][35] , \p[17][34] , \p[17][33] , \p[17][32] ,
         \p[17][31] , \p[17][30] , \p[17][29] , \p[17][28] , \p[17][27] ,
         \p[17][26] , \p[17][25] , \p[17][24] , \p[17][23] , \p[17][22] ,
         \p[17][21] , \p[17][20] , \p[17][19] , \p[17][18] , \p[17][17] ,
         \p[16][63] , \p[16][46] , \p[16][45] , \p[16][44] , \p[16][43] ,
         \p[16][42] , \p[16][41] , \p[16][40] , \p[16][39] , \p[16][38] ,
         \p[16][37] , \p[16][36] , \p[16][35] , \p[16][34] , \p[16][33] ,
         \p[16][32] , \p[16][31] , \p[16][30] , \p[16][29] , \p[16][28] ,
         \p[16][27] , \p[16][26] , \p[16][25] , \p[16][24] , \p[16][23] ,
         \p[16][22] , \p[16][21] , \p[16][20] , \p[16][19] , \p[16][18] ,
         \p[16][17] , \p[16][16] , \p[15][63] , \p[15][45] , \p[15][44] ,
         \p[15][43] , \p[15][42] , \p[15][41] , \p[15][40] , \p[15][39] ,
         \p[15][38] , \p[15][37] , \p[15][36] , \p[15][35] , \p[15][34] ,
         \p[15][33] , \p[15][32] , \p[15][31] , \p[15][30] , \p[15][29] ,
         \p[15][28] , \p[15][27] , \p[15][26] , \p[15][25] , \p[15][24] ,
         \p[15][23] , \p[15][22] , \p[15][21] , \p[15][20] , \p[15][19] ,
         \p[15][18] , \p[15][17] , \p[15][16] , \p[15][15] , \p[14][63] ,
         \p[14][44] , \p[14][43] , \p[14][42] , \p[14][41] , \p[14][40] ,
         \p[14][39] , \p[14][38] , \p[14][37] , \p[14][36] , \p[14][35] ,
         \p[14][34] , \p[14][33] , \p[14][32] , \p[14][31] , \p[14][30] ,
         \p[14][29] , \p[14][28] , \p[14][27] , \p[14][26] , \p[14][25] ,
         \p[14][24] , \p[14][23] , \p[14][22] , \p[14][21] , \p[14][20] ,
         \p[14][19] , \p[14][18] , \p[14][17] , \p[14][16] , \p[14][15] ,
         \p[14][14] , \p[13][63] , \p[13][43] , \p[13][42] , \p[13][41] ,
         \p[13][40] , \p[13][39] , \p[13][38] , \p[13][37] , \p[13][36] ,
         \p[13][35] , \p[13][34] , \p[13][33] , \p[13][32] , \p[13][31] ,
         \p[13][30] , \p[13][29] , \p[13][28] , \p[13][27] , \p[13][26] ,
         \p[13][25] , \p[13][24] , \p[13][23] , \p[13][22] , \p[13][21] ,
         \p[13][20] , \p[13][19] , \p[13][18] , \p[13][17] , \p[13][16] ,
         \p[13][15] , \p[13][14] , \p[13][13] , \p[12][63] , \p[12][42] ,
         \p[12][41] , \p[12][40] , \p[12][39] , \p[12][38] , \p[12][37] ,
         \p[12][36] , \p[12][35] , \p[12][34] , \p[12][33] , \p[12][32] ,
         \p[12][31] , \p[12][30] , \p[12][29] , \p[12][28] , \p[12][27] ,
         \p[12][26] , \p[12][25] , \p[12][24] , \p[12][23] , \p[12][22] ,
         \p[12][21] , \p[12][20] , \p[12][19] , \p[12][18] , \p[12][17] ,
         \p[12][16] , \p[12][15] , \p[12][14] , \p[12][13] , \p[12][12] ,
         \p[11][63] , \p[11][41] , \p[11][40] , \p[11][39] , \p[11][38] ,
         \p[11][37] , \p[11][36] , \p[11][35] , \p[11][34] , \p[11][33] ,
         \p[11][32] , \p[11][31] , \p[11][30] , \p[11][29] , \p[11][28] ,
         \p[11][27] , \p[11][26] , \p[11][25] , \p[11][24] , \p[11][23] ,
         \p[11][22] , \p[11][21] , \p[11][20] , \p[11][19] , \p[11][18] ,
         \p[11][17] , \p[11][16] , \p[11][15] , \p[11][14] , \p[11][13] ,
         \p[11][12] , \p[11][11] , \p[10][63] , \p[10][40] , \p[10][39] ,
         \p[10][38] , \p[10][37] , \p[10][36] , \p[10][35] , \p[10][34] ,
         \p[10][33] , \p[10][32] , \p[10][31] , \p[10][30] , \p[10][29] ,
         \p[10][28] , \p[10][27] , \p[10][26] , \p[10][25] , \p[10][24] ,
         \p[10][23] , \p[10][22] , \p[10][21] , \p[10][20] , \p[10][19] ,
         \p[10][18] , \p[10][17] , \p[10][16] , \p[10][15] , \p[10][14] ,
         \p[10][13] , \p[10][12] , \p[10][11] , \p[10][10] , \p[9][63] ,
         \p[9][39] , \p[9][38] , \p[9][37] , \p[9][36] , \p[9][35] ,
         \p[9][34] , \p[9][33] , \p[9][32] , \p[9][31] , \p[9][30] ,
         \p[9][29] , \p[9][28] , \p[9][27] , \p[9][26] , \p[9][25] ,
         \p[9][24] , \p[9][23] , \p[9][22] , \p[9][21] , \p[9][20] ,
         \p[9][19] , \p[9][18] , \p[9][17] , \p[9][16] , \p[9][15] ,
         \p[9][14] , \p[9][13] , \p[9][12] , \p[9][11] , \p[9][10] , \p[9][9] ,
         \p[8][63] , \p[8][38] , \p[8][37] , \p[8][36] , \p[8][35] ,
         \p[8][34] , \p[8][33] , \p[8][32] , \p[8][31] , \p[8][30] ,
         \p[8][29] , \p[8][28] , \p[8][27] , \p[8][26] , \p[8][25] ,
         \p[8][24] , \p[8][23] , \p[8][22] , \p[8][21] , \p[8][20] ,
         \p[8][19] , \p[8][18] , \p[8][17] , \p[8][16] , \p[8][15] ,
         \p[8][14] , \p[8][13] , \p[8][12] , \p[8][11] , \p[8][10] , \p[8][9] ,
         \p[8][8] , \g[41][63] , \g[41][62] , \g[41][61] , \g[41][60] ,
         \g[41][59] , \g[41][58] , \g[41][57] , \g[41][56] , \g[41][55] ,
         \g[41][54] , \g[41][53] , \g[41][52] , \g[41][51] , \g[41][50] ,
         \g[41][49] , \g[41][48] , \g[41][47] , \g[41][46] , \g[41][45] ,
         \g[41][44] , \g[41][43] , \g[41][42] , \g[41][41] , \g[41][40] ,
         \g[41][39] , \g[41][38] , \g[41][37] , \g[41][36] , \g[41][35] ,
         \g[41][34] , \g[41][33] , \g[41][32] , \g[41][31] , \g[41][30] ,
         \g[41][29] , \g[41][28] , \g[41][27] , \g[41][26] , \g[41][25] ,
         \g[41][24] , \g[41][23] , \g[41][22] , \g[41][21] , \g[41][20] ,
         \g[41][19] , \g[41][18] , \g[41][17] , \g[41][16] , \g[41][15] ,
         \g[41][14] , \g[41][13] , \g[41][12] , \g[41][11] , \g[41][10] ,
         \g[41][9] , \g[41][8] , \g[41][7] , \g[41][6] , \g[41][5] ,
         \g[41][4] , \g[41][3] , \g[41][2] , \g[41][1] , \g[40][63] ,
         \g[40][62] , \g[40][61] , \g[40][60] , \g[40][59] , \g[40][58] ,
         \g[40][57] , \g[40][56] , \g[40][55] , \g[40][54] , \g[40][53] ,
         \g[40][52] , \g[40][51] , \g[40][50] , \g[40][49] , \g[40][48] ,
         \g[40][47] , \g[40][46] , \g[40][45] , \g[40][44] , \g[40][43] ,
         \g[40][42] , \g[40][41] , \g[40][40] , \g[40][39] , \g[40][38] ,
         \g[40][37] , \g[40][36] , \g[40][35] , \g[40][34] , \g[40][33] ,
         \g[40][32] , \g[40][31] , \g[40][30] , \g[40][29] , \g[40][28] ,
         \g[40][27] , \g[40][26] , \g[40][25] , \g[40][24] , \g[40][23] ,
         \g[40][22] , \g[40][21] , \g[40][20] , \g[40][19] , \g[40][18] ,
         \g[40][17] , \g[40][16] , \g[40][15] , \g[40][14] , \g[40][13] ,
         \g[40][12] , \g[40][11] , \g[40][10] , \g[40][9] , \g[40][8] ,
         \g[40][7] , \g[40][6] , \g[40][5] , \g[40][4] , \g[40][3] ,
         \g[40][2] , \g[40][1] , \g[39][63] , \g[39][62] , \g[39][61] ,
         \g[39][60] , \g[39][59] , \g[39][58] , \g[39][57] , \g[39][56] ,
         \g[39][55] , \g[39][54] , \g[39][53] , \g[39][52] , \g[39][51] ,
         \g[39][50] , \g[39][49] , \g[39][48] , \g[39][47] , \g[39][46] ,
         \g[39][45] , \g[39][44] , \g[39][43] , \g[39][42] , \g[39][41] ,
         \g[39][40] , \g[39][39] , \g[39][38] , \g[39][37] , \g[39][36] ,
         \g[39][35] , \g[39][34] , \g[39][33] , \g[39][32] , \g[39][31] ,
         \g[39][30] , \g[39][29] , \g[39][28] , \g[39][27] , \g[39][26] ,
         \g[39][25] , \g[39][24] , \g[39][23] , \g[39][22] , \g[39][21] ,
         \g[39][20] , \g[39][19] , \g[39][18] , \g[39][17] , \g[39][16] ,
         \g[39][15] , \g[39][14] , \g[39][13] , \g[39][12] , \g[39][11] ,
         \g[39][10] , \g[39][9] , \g[39][8] , \g[39][7] , \g[39][6] ,
         \g[39][5] , \g[39][4] , \g[39][3] , \g[39][2] , \g[39][1] ,
         \g[38][63] , \g[38][62] , \g[38][61] , \g[38][60] , \g[38][59] ,
         \g[38][58] , \g[38][57] , \g[38][56] , \g[38][55] , \g[38][54] ,
         \g[38][53] , \g[38][52] , \g[38][51] , \g[38][50] , \g[38][49] ,
         \g[38][48] , \g[38][47] , \g[38][46] , \g[38][45] , \g[38][44] ,
         \g[38][43] , \g[38][42] , \g[38][41] , \g[38][40] , \g[38][39] ,
         \g[38][38] , \g[38][37] , \g[38][36] , \g[38][35] , \g[38][34] ,
         \g[38][33] , \g[38][32] , \g[38][31] , \g[38][30] , \g[38][29] ,
         \g[38][28] , \g[38][27] , \g[38][26] , \g[38][25] , \g[38][24] ,
         \g[38][23] , \g[38][22] , \g[38][21] , \g[38][20] , \g[38][19] ,
         \g[38][18] , \g[38][17] , \g[38][16] , \g[38][15] , \g[38][14] ,
         \g[38][13] , \g[38][12] , \g[38][11] , \g[38][10] , \g[38][9] ,
         \g[38][8] , \g[38][7] , \g[38][6] , \g[38][5] , \g[38][4] ,
         \g[38][3] , \g[38][2] , \g[38][1] , \g[37][63] , \g[37][62] ,
         \g[37][61] , \g[37][60] , \g[37][59] , \g[37][58] , \g[37][57] ,
         \g[37][56] , \g[37][55] , \g[37][54] , \g[37][53] , \g[37][52] ,
         \g[37][51] , \g[37][50] , \g[37][49] , \g[37][48] , \g[37][47] ,
         \g[37][46] , \g[37][45] , \g[37][44] , \g[37][43] , \g[37][42] ,
         \g[37][41] , \g[37][40] , \g[37][39] , \g[37][38] , \g[37][37] ,
         \g[37][36] , \g[37][35] , \g[37][34] , \g[37][33] , \g[37][32] ,
         \g[37][31] , \g[37][30] , \g[37][29] , \g[37][28] , \g[37][27] ,
         \g[37][26] , \g[37][25] , \g[37][24] , \g[37][23] , \g[37][22] ,
         \g[37][21] , \g[37][20] , \g[37][19] , \g[37][18] , \g[37][17] ,
         \g[37][16] , \g[37][15] , \g[37][14] , \g[37][13] , \g[37][12] ,
         \g[37][11] , \g[37][10] , \g[37][9] , \g[37][8] , \g[37][7] ,
         \g[37][6] , \g[37][5] , \g[37][4] , \g[37][3] , \g[37][2] ,
         \g[37][1] , \g[36][63] , \g[36][62] , \g[36][61] , \g[36][60] ,
         \g[36][59] , \g[36][58] , \g[36][57] , \g[36][56] , \g[36][55] ,
         \g[36][54] , \g[36][53] , \g[36][52] , \g[36][51] , \g[36][50] ,
         \g[36][49] , \g[36][48] , \g[36][47] , \g[36][46] , \g[36][45] ,
         \g[36][44] , \g[36][43] , \g[36][42] , \g[36][41] , \g[36][40] ,
         \g[36][39] , \g[36][38] , \g[36][37] , \g[36][36] , \g[36][35] ,
         \g[36][34] , \g[36][33] , \g[36][32] , \g[36][31] , \g[36][30] ,
         \g[36][29] , \g[36][28] , \g[36][27] , \g[36][26] , \g[36][25] ,
         \g[36][24] , \g[36][23] , \g[36][22] , \g[36][21] , \g[36][20] ,
         \g[36][19] , \g[36][18] , \g[36][17] , \g[36][16] , \g[36][15] ,
         \g[36][14] , \g[36][13] , \g[36][12] , \g[36][11] , \g[36][10] ,
         \g[36][9] , \g[36][8] , \g[36][7] , \g[36][6] , \g[36][5] ,
         \g[36][4] , \g[36][3] , \g[36][2] , \g[36][1] , \g[35][63] ,
         \g[35][62] , \g[35][61] , \g[35][60] , \g[35][59] , \g[35][58] ,
         \g[35][57] , \g[35][56] , \g[35][55] , \g[35][54] , \g[35][53] ,
         \g[35][52] , \g[35][51] , \g[35][50] , \g[35][49] , \g[35][48] ,
         \g[35][47] , \g[35][46] , \g[35][45] , \g[35][44] , \g[35][43] ,
         \g[35][42] , \g[35][41] , \g[35][40] , \g[35][39] , \g[35][38] ,
         \g[35][37] , \g[35][36] , \g[35][35] , \g[35][34] , \g[35][33] ,
         \g[35][32] , \g[35][31] , \g[35][30] , \g[35][29] , \g[35][28] ,
         \g[35][27] , \g[35][26] , \g[35][25] , \g[35][24] , \g[35][23] ,
         \g[35][22] , \g[35][21] , \g[35][20] , \g[35][19] , \g[35][18] ,
         \g[35][17] , \g[35][16] , \g[35][15] , \g[35][14] , \g[35][13] ,
         \g[35][12] , \g[35][11] , \g[35][10] , \g[35][9] , \g[35][8] ,
         \g[35][7] , \g[35][6] , \g[35][5] , \g[35][4] , \g[35][3] ,
         \g[35][2] , \g[35][1] , \g[34][63] , \g[34][62] , \g[34][61] ,
         \g[34][60] , \g[34][59] , \g[34][58] , \g[34][57] , \g[34][56] ,
         \g[34][55] , \g[34][54] , \g[34][53] , \g[34][52] , \g[34][51] ,
         \g[34][50] , \g[34][49] , \g[34][48] , \g[34][47] , \g[34][46] ,
         \g[34][45] , \g[34][44] , \g[34][43] , \g[34][42] , \g[34][41] ,
         \g[34][40] , \g[34][39] , \g[34][38] , \g[34][37] , \g[34][36] ,
         \g[34][35] , \g[34][34] , \g[34][33] , \g[34][32] , \g[34][31] ,
         \g[34][30] , \g[34][29] , \g[34][28] , \g[34][27] , \g[34][26] ,
         \g[34][25] , \g[34][24] , \g[34][23] , \g[34][22] , \g[34][21] ,
         \g[34][20] , \g[34][19] , \g[34][18] , \g[34][17] , \g[34][16] ,
         \g[34][15] , \g[34][14] , \g[34][13] , \g[34][12] , \g[34][11] ,
         \g[34][10] , \g[34][9] , \g[34][8] , \g[34][7] , \g[34][6] ,
         \g[34][5] , \g[34][4] , \g[34][3] , \g[34][2] , \g[34][1] ,
         \g[33][63] , \g[33][62] , \g[33][61] , \g[33][60] , \g[33][59] ,
         \g[33][58] , \g[33][57] , \g[33][56] , \g[33][55] , \g[33][54] ,
         \g[33][53] , \g[33][52] , \g[33][51] , \g[33][50] , \g[33][49] ,
         \g[33][48] , \g[33][47] , \g[33][46] , \g[33][45] , \g[33][44] ,
         \g[33][43] , \g[33][42] , \g[33][41] , \g[33][40] , \g[33][39] ,
         \g[33][38] , \g[33][37] , \g[33][36] , \g[33][35] , \g[33][34] ,
         \g[33][33] , \g[33][32] , \g[33][31] , \g[33][30] , \g[33][29] ,
         \g[33][28] , \g[33][27] , \g[33][26] , \g[33][25] , \g[33][24] ,
         \g[33][23] , \g[33][22] , \g[33][21] , \g[33][20] , \g[33][19] ,
         \g[33][18] , \g[33][17] , \g[33][16] , \g[33][15] , \g[33][14] ,
         \g[33][13] , \g[33][12] , \g[33][11] , \g[33][10] , \g[33][9] ,
         \g[33][8] , \g[33][7] , \g[33][6] , \g[33][5] , \g[33][4] ,
         \g[33][3] , \g[33][2] , \g[33][1] , \g[32][63] , \g[32][62] ,
         \g[32][61] , \g[32][60] , \g[32][59] , \g[32][58] , \g[32][57] ,
         \g[32][56] , \g[32][55] , \g[32][54] , \g[32][53] , \g[32][52] ,
         \g[32][51] , \g[32][50] , \g[32][49] , \g[32][48] , \g[32][47] ,
         \g[32][46] , \g[32][45] , \g[32][44] , \g[32][43] , \g[32][42] ,
         \g[32][41] , \g[32][40] , \g[32][39] , \g[32][38] , \g[32][37] ,
         \g[32][36] , \g[32][35] , \g[32][34] , \g[32][33] , \g[32][32] ,
         \g[32][31] , \g[32][30] , \g[32][29] , \g[32][28] , \g[32][27] ,
         \g[32][26] , \g[32][25] , \g[32][24] , \g[32][23] , \g[32][22] ,
         \g[32][21] , \g[32][20] , \g[32][19] , \g[32][18] , \g[32][17] ,
         \g[32][16] , \g[32][15] , \g[32][14] , \g[32][13] , \g[32][12] ,
         \g[32][11] , \g[32][10] , \g[32][9] , \g[32][8] , \g[32][7] ,
         \g[32][6] , \g[32][5] , \g[32][4] , \g[32][3] , \g[32][2] ,
         \g[32][1] , \g[31][63] , \g[31][62] , \g[31][61] , \g[31][60] ,
         \g[31][59] , \g[31][58] , \g[31][57] , \g[31][56] , \g[31][55] ,
         \g[31][54] , \g[31][53] , \g[31][52] , \g[31][51] , \g[31][50] ,
         \g[31][49] , \g[31][48] , \g[31][47] , \g[31][46] , \g[31][45] ,
         \g[31][44] , \g[31][43] , \g[31][42] , \g[31][41] , \g[31][40] ,
         \g[31][39] , \g[31][38] , \g[31][37] , \g[31][36] , \g[31][35] ,
         \g[31][34] , \g[31][33] , \g[31][32] , \g[31][31] , \g[31][30] ,
         \g[31][29] , \g[31][28] , \g[31][27] , \g[31][26] , \g[31][25] ,
         \g[31][24] , \g[31][23] , \g[31][22] , \g[31][21] , \g[31][20] ,
         \g[31][19] , \g[31][18] , \g[31][17] , \g[31][16] , \g[31][15] ,
         \g[31][14] , \g[31][13] , \g[31][12] , \g[31][11] , \g[31][10] ,
         \g[31][9] , \g[31][8] , \g[31][7] , \g[31][6] , \g[31][5] ,
         \g[31][4] , \g[31][3] , \g[31][2] , \g[31][1] , \g[30][63] ,
         \g[30][62] , \g[30][61] , \g[30][60] , \g[30][59] , \g[30][58] ,
         \g[30][57] , \g[30][56] , \g[30][55] , \g[30][54] , \g[30][53] ,
         \g[30][52] , \g[30][51] , \g[30][50] , \g[30][49] , \g[30][48] ,
         \g[30][47] , \g[30][46] , \g[30][45] , \g[30][44] , \g[30][43] ,
         \g[30][42] , \g[30][41] , \g[30][40] , \g[30][39] , \g[30][38] ,
         \g[30][37] , \g[30][36] , \g[30][35] , \g[30][34] , \g[30][33] ,
         \g[30][32] , \g[30][31] , \g[30][30] , \g[30][29] , \g[30][28] ,
         \g[30][27] , \g[30][26] , \g[30][25] , \g[30][24] , \g[30][23] ,
         \g[30][22] , \g[30][21] , \g[30][20] , \g[30][19] , \g[30][18] ,
         \g[30][17] , \g[30][16] , \g[30][15] , \g[30][14] , \g[30][13] ,
         \g[30][12] , \g[30][11] , \g[30][10] , \g[30][9] , \g[30][8] ,
         \g[30][7] , \g[30][6] , \g[30][5] , \g[30][4] , \g[30][3] ,
         \g[30][2] , \g[30][1] , \g[29][63] , \g[29][62] , \g[29][61] ,
         \g[29][60] , \g[29][59] , \g[29][58] , \g[29][57] , \g[29][56] ,
         \g[29][55] , \g[29][54] , \g[29][53] , \g[29][52] , \g[29][51] ,
         \g[29][50] , \g[29][49] , \g[29][48] , \g[29][47] , \g[29][46] ,
         \g[29][45] , \g[29][44] , \g[29][43] , \g[29][42] , \g[29][41] ,
         \g[29][40] , \g[29][39] , \g[29][38] , \g[29][37] , \g[29][36] ,
         \g[29][35] , \g[29][34] , \g[29][33] , \g[29][32] , \g[29][31] ,
         \g[29][30] , \g[29][29] , \g[29][28] , \g[29][27] , \g[29][26] ,
         \g[29][25] , \g[29][24] , \g[29][23] , \g[29][22] , \g[29][21] ,
         \g[29][20] , \g[29][19] , \g[29][18] , \g[29][17] , \g[29][16] ,
         \g[29][15] , \g[29][14] , \g[29][13] , \g[29][12] , \g[29][11] ,
         \g[29][10] , \g[29][9] , \g[29][8] , \g[29][7] , \g[29][6] ,
         \g[29][5] , \g[29][4] , \g[29][3] , \g[29][2] , \g[29][1] ,
         \g[28][63] , \g[28][62] , \g[28][61] , \g[28][60] , \g[28][59] ,
         \g[28][58] , \g[28][57] , \g[28][56] , \g[28][55] , \g[28][54] ,
         \g[28][53] , \g[28][52] , \g[28][51] , \g[28][50] , \g[28][49] ,
         \g[28][48] , \g[28][47] , \g[28][46] , \g[28][45] , \g[28][44] ,
         \g[28][43] , \g[28][42] , \g[28][41] , \g[28][40] , \g[28][39] ,
         \g[28][38] , \g[28][37] , \g[28][36] , \g[28][35] , \g[28][34] ,
         \g[28][33] , \g[28][32] , \g[28][31] , \g[28][30] , \g[28][29] ,
         \g[28][28] , \g[28][27] , \g[28][26] , \g[28][25] , \g[28][24] ,
         \g[28][23] , \g[28][22] , \g[28][21] , \g[28][20] , \g[28][19] ,
         \g[28][18] , \g[28][17] , \g[28][16] , \g[28][15] , \g[28][14] ,
         \g[28][13] , \g[28][12] , \g[28][11] , \g[28][10] , \g[28][9] ,
         \g[28][8] , \g[28][7] , \g[28][6] , \g[28][5] , \g[28][4] ,
         \g[28][3] , \g[28][2] , \g[28][1] , \g[27][63] , \g[27][62] ,
         \g[27][61] , \g[27][60] , \g[27][59] , \g[27][58] , \g[27][57] ,
         \g[27][56] , \g[27][55] , \g[27][54] , \g[27][53] , \g[27][52] ,
         \g[27][51] , \g[27][50] , \g[27][49] , \g[27][48] , \g[27][47] ,
         \g[27][46] , \g[27][45] , \g[27][44] , \g[27][43] , \g[27][42] ,
         \g[27][41] , \g[27][40] , \g[27][39] , \g[27][38] , \g[27][37] ,
         \g[27][36] , \g[27][35] , \g[27][34] , \g[27][33] , \g[27][32] ,
         \g[27][31] , \g[27][30] , \g[27][29] , \g[27][28] , \g[27][27] ,
         \g[27][26] , \g[27][25] , \g[27][24] , \g[27][23] , \g[27][22] ,
         \g[27][21] , \g[27][20] , \g[27][19] , \g[27][18] , \g[27][17] ,
         \g[27][16] , \g[27][15] , \g[27][14] , \g[27][13] , \g[27][12] ,
         \g[27][11] , \g[27][10] , \g[27][9] , \g[27][8] , \g[27][7] ,
         \g[27][6] , \g[27][5] , \g[27][4] , \g[27][3] , \g[27][2] ,
         \g[27][1] , \g[26][63] , \g[26][62] , \g[26][61] , \g[26][60] ,
         \g[26][59] , \g[26][58] , \g[26][57] , \g[26][56] , \g[26][55] ,
         \g[26][54] , \g[26][53] , \g[26][52] , \g[26][51] , \g[26][50] ,
         \g[26][49] , \g[26][48] , \g[26][47] , \g[26][46] , \g[26][45] ,
         \g[26][44] , \g[26][43] , \g[26][42] , \g[26][41] , \g[26][40] ,
         \g[26][39] , \g[26][38] , \g[26][37] , \g[26][36] , \g[26][35] ,
         \g[26][34] , \g[26][33] , \g[26][32] , \g[26][31] , \g[26][30] ,
         \g[26][29] , \g[26][28] , \g[26][27] , \g[26][26] , \g[26][25] ,
         \g[26][24] , \g[26][23] , \g[26][22] , \g[26][21] , \g[26][20] ,
         \g[26][19] , \g[26][18] , \g[26][17] , \g[26][16] , \g[26][15] ,
         \g[26][14] , \g[26][13] , \g[26][12] , \g[26][11] , \g[26][10] ,
         \g[26][9] , \g[26][8] , \g[26][7] , \g[26][6] , \g[26][5] ,
         \g[26][4] , \g[26][3] , \g[26][2] , \g[26][1] , \g[25][63] ,
         \g[25][62] , \g[25][61] , \g[25][60] , \g[25][59] , \g[25][58] ,
         \g[25][57] , \g[25][56] , \g[25][55] , \g[25][54] , \g[25][53] ,
         \g[25][52] , \g[25][51] , \g[25][50] , \g[25][49] , \g[25][48] ,
         \g[25][47] , \g[25][46] , \g[25][45] , \g[25][44] , \g[25][43] ,
         \g[25][42] , \g[25][41] , \g[25][40] , \g[25][39] , \g[25][38] ,
         \g[25][37] , \g[25][36] , \g[25][35] , \g[25][34] , \g[25][33] ,
         \g[25][32] , \g[25][31] , \g[25][30] , \g[25][29] , \g[25][28] ,
         \g[25][27] , \g[25][26] , \g[25][25] , \g[25][24] , \g[25][23] ,
         \g[25][22] , \g[25][21] , \g[25][20] , \g[25][19] , \g[25][18] ,
         \g[25][17] , \g[25][16] , \g[25][15] , \g[25][14] , \g[25][13] ,
         \g[25][12] , \g[25][11] , \g[25][10] , \g[25][9] , \g[25][8] ,
         \g[25][7] , \g[25][6] , \g[25][5] , \g[25][4] , \g[25][3] ,
         \g[25][2] , \g[25][1] , \g[24][63] , \g[24][62] , \g[24][61] ,
         \g[24][60] , \g[24][59] , \g[24][58] , \g[24][57] , \g[24][56] ,
         \g[24][55] , \g[24][54] , \g[24][53] , \g[24][52] , \g[24][51] ,
         \g[24][50] , \g[24][49] , \g[24][48] , \g[24][47] , \g[24][46] ,
         \g[24][45] , \g[24][44] , \g[24][43] , \g[24][42] , \g[24][41] ,
         \g[24][40] , \g[24][39] , \g[24][38] , \g[24][37] , \g[24][36] ,
         \g[24][35] , \g[24][34] , \g[24][33] , \g[24][32] , \g[24][31] ,
         \g[24][30] , \g[24][29] , \g[24][28] , \g[24][27] , \g[24][26] ,
         \g[24][25] , \g[24][24] , \g[24][23] , \g[24][22] , \g[24][21] ,
         \g[24][20] , \g[24][19] , \g[24][18] , \g[24][17] , \g[24][16] ,
         \g[24][15] , \g[24][14] , \g[24][13] , \g[24][12] , \g[24][11] ,
         \g[24][10] , \g[24][9] , \g[24][8] , \g[24][7] , \g[24][6] ,
         \g[24][5] , \g[24][4] , \g[24][3] , \g[24][2] , \g[24][1] ,
         \g[23][63] , \g[23][62] , \g[23][61] , \g[23][60] , \g[23][59] ,
         \g[23][58] , \g[23][57] , \g[23][56] , \g[23][55] , \g[23][54] ,
         \g[23][53] , \g[23][52] , \g[23][51] , \g[23][50] , \g[23][49] ,
         \g[23][48] , \g[23][47] , \g[23][46] , \g[23][45] , \g[23][44] ,
         \g[23][43] , \g[23][42] , \g[23][41] , \g[23][40] , \g[23][39] ,
         \g[23][38] , \g[23][37] , \g[23][36] , \g[23][35] , \g[23][34] ,
         \g[23][33] , \g[23][32] , \g[23][31] , \g[23][30] , \g[23][29] ,
         \g[23][28] , \g[23][27] , \g[23][26] , \g[23][25] , \g[23][24] ,
         \g[23][23] , \g[23][22] , \g[23][21] , \g[23][20] , \g[23][19] ,
         \g[23][18] , \g[23][17] , \g[23][16] , \g[23][15] , \g[23][14] ,
         \g[23][13] , \g[23][12] , \g[23][11] , \g[23][10] , \g[23][9] ,
         \g[23][8] , \g[23][7] , \g[23][6] , \g[23][5] , \g[23][4] ,
         \g[23][3] , \g[23][2] , \g[23][1] , \g[22][63] , \g[22][62] ,
         \g[22][61] , \g[22][60] , \g[22][59] , \g[22][58] , \g[22][57] ,
         \g[22][56] , \g[22][55] , \g[22][54] , \g[22][53] , \g[22][52] ,
         \g[22][51] , \g[22][50] , \g[22][49] , \g[22][48] , \g[22][47] ,
         \g[22][46] , \g[22][45] , \g[22][44] , \g[22][43] , \g[22][42] ,
         \g[22][41] , \g[22][40] , \g[22][39] , \g[22][38] , \g[22][37] ,
         \g[22][36] , \g[22][35] , \g[22][34] , \g[22][33] , \g[22][32] ,
         \g[22][31] , \g[22][30] , \g[22][29] , \g[22][28] , \g[22][27] ,
         \g[22][26] , \g[22][25] , \g[22][24] , \g[22][23] , \g[22][22] ,
         \g[22][21] , \g[22][20] , \g[22][19] , \g[22][18] , \g[22][17] ,
         \g[22][16] , \g[22][15] , \g[22][14] , \g[22][13] , \g[22][12] ,
         \g[22][11] , \g[22][10] , \g[22][9] , \g[22][8] , \g[22][7] ,
         \g[22][6] , \g[22][5] , \g[22][4] , \g[22][3] , \g[22][2] ,
         \g[22][1] , \g[21][63] , \g[21][62] , \g[21][61] , \g[21][60] ,
         \g[21][59] , \g[21][58] , \g[21][57] , \g[21][56] , \g[21][55] ,
         \g[21][54] , \g[21][53] , \g[21][52] , \g[21][51] , \g[21][50] ,
         \g[21][49] , \g[21][48] , \g[21][47] , \g[21][46] , \g[21][45] ,
         \g[21][44] , \g[21][43] , \g[21][42] , \g[21][41] , \g[21][40] ,
         \g[21][39] , \g[21][38] , \g[21][37] , \g[21][36] , \g[21][35] ,
         \g[21][34] , \g[21][33] , \g[21][32] , \g[21][31] , \g[21][30] ,
         \g[21][29] , \g[21][28] , \g[21][27] , \g[21][26] , \g[21][25] ,
         \g[21][24] , \g[21][23] , \g[21][22] , \g[21][21] , \g[21][20] ,
         \g[21][19] , \g[21][18] , \g[21][17] , \g[21][16] , \g[21][15] ,
         \g[21][14] , \g[21][13] , \g[21][12] , \g[21][11] , \g[21][10] ,
         \g[21][9] , \g[21][8] , \g[21][7] , \g[21][6] , \g[21][5] ,
         \g[21][4] , \g[21][3] , \g[21][2] , \g[21][1] , \g[20][63] ,
         \g[20][62] , \g[20][61] , \g[20][60] , \g[20][59] , \g[20][58] ,
         \g[20][57] , \g[20][56] , \g[20][55] , \g[20][54] , \g[20][53] ,
         \g[20][52] , \g[20][51] , \g[20][50] , \g[20][49] , \g[20][48] ,
         \g[20][47] , \g[20][46] , \g[20][45] , \g[20][44] , \g[20][43] ,
         \g[20][42] , \g[20][41] , \g[20][40] , \g[20][39] , \g[20][38] ,
         \g[20][37] , \g[20][36] , \g[20][35] , \g[20][34] , \g[20][33] ,
         \g[20][32] , \g[20][31] , \g[20][30] , \g[20][29] , \g[20][28] ,
         \g[20][27] , \g[20][26] , \g[20][25] , \g[20][24] , \g[20][23] ,
         \g[20][22] , \g[20][21] , \g[20][20] , \g[20][19] , \g[20][18] ,
         \g[20][17] , \g[20][16] , \g[20][15] , \g[20][14] , \g[20][13] ,
         \g[20][12] , \g[20][11] , \g[20][10] , \g[20][9] , \g[20][8] ,
         \g[20][7] , \g[20][6] , \g[20][5] , \g[20][4] , \g[20][3] ,
         \g[20][2] , \g[20][1] , \g[20][0] , \g[19][63] , \g[19][62] ,
         \g[19][61] , \g[19][60] , \g[19][59] , \g[19][58] , \g[19][57] ,
         \g[19][56] , \g[19][55] , \g[19][54] , \g[19][53] , \g[19][52] ,
         \g[19][51] , \g[19][50] , \g[19][49] , \g[19][48] , \g[19][47] ,
         \g[19][46] , \g[19][45] , \g[19][44] , \g[19][43] , \g[19][42] ,
         \g[19][41] , \g[19][40] , \g[19][39] , \g[19][38] , \g[19][37] ,
         \g[19][36] , \g[19][35] , \g[19][34] , \g[19][33] , \g[19][32] ,
         \g[19][31] , \g[19][30] , \g[19][29] , \g[19][28] , \g[19][27] ,
         \g[19][26] , \g[19][25] , \g[19][24] , \g[19][23] , \g[19][22] ,
         \g[19][21] , \g[19][20] , \g[19][19] , \g[19][18] , \g[19][17] ,
         \g[19][16] , \g[19][15] , \g[19][14] , \g[19][13] , \g[19][12] ,
         \g[19][11] , \g[19][10] , \g[19][9] , \g[19][8] , \g[19][7] ,
         \g[19][6] , \g[19][5] , \g[19][4] , \g[19][3] , \g[19][2] ,
         \g[19][1] , \g[19][0] , \g[18][63] , \g[18][62] , \g[18][61] ,
         \g[18][60] , \g[18][59] , \g[18][58] , \g[18][57] , \g[18][56] ,
         \g[18][55] , \g[18][54] , \g[18][53] , \g[18][52] , \g[18][51] ,
         \g[18][50] , \g[18][49] , \g[18][48] , \g[18][47] , \g[18][46] ,
         \g[18][45] , \g[18][44] , \g[18][43] , \g[18][42] , \g[18][41] ,
         \g[18][40] , \g[18][39] , \g[18][38] , \g[18][37] , \g[18][36] ,
         \g[18][35] , \g[18][34] , \g[18][33] , \g[18][32] , \g[18][31] ,
         \g[18][30] , \g[18][29] , \g[18][28] , \g[18][27] , \g[18][26] ,
         \g[18][25] , \g[18][24] , \g[18][23] , \g[18][22] , \g[18][21] ,
         \g[18][20] , \g[18][19] , \g[18][18] , \g[18][17] , \g[18][16] ,
         \g[18][15] , \g[18][14] , \g[18][13] , \g[18][12] , \g[18][11] ,
         \g[18][10] , \g[18][9] , \g[18][8] , \g[18][7] , \g[18][6] ,
         \g[18][5] , \g[18][4] , \g[18][3] , \g[18][2] , \g[18][1] ,
         \g[18][0] , \g[17][63] , \g[17][62] , \g[17][61] , \g[17][60] ,
         \g[17][59] , \g[17][58] , \g[17][57] , \g[17][56] , \g[17][55] ,
         \g[17][54] , \g[17][53] , \g[17][52] , \g[17][51] , \g[17][50] ,
         \g[17][49] , \g[17][48] , \g[17][47] , \g[17][46] , \g[17][45] ,
         \g[17][44] , \g[17][43] , \g[17][42] , \g[17][41] , \g[17][40] ,
         \g[17][39] , \g[17][38] , \g[17][37] , \g[17][36] , \g[17][35] ,
         \g[17][34] , \g[17][33] , \g[17][32] , \g[17][31] , \g[17][30] ,
         \g[17][29] , \g[17][28] , \g[17][27] , \g[17][26] , \g[17][25] ,
         \g[17][24] , \g[17][23] , \g[17][22] , \g[17][21] , \g[17][20] ,
         \g[17][19] , \g[17][18] , \g[17][17] , \g[17][16] , \g[17][15] ,
         \g[17][14] , \g[17][13] , \g[17][12] , \g[17][11] , \g[17][10] ,
         \g[17][9] , \g[17][8] , \g[17][7] , \g[17][6] , \g[17][5] ,
         \g[17][4] , \g[17][3] , \g[17][2] , \g[17][1] , \g[17][0] ,
         \g[16][63] , \g[16][62] , \g[16][61] , \g[16][60] , \g[16][59] ,
         \g[16][58] , \g[16][57] , \g[16][56] , \g[16][55] , \g[16][54] ,
         \g[16][53] , \g[16][52] , \g[16][51] , \g[16][50] , \g[16][49] ,
         \g[16][48] , \g[16][47] , \g[16][46] , \g[16][45] , \g[16][44] ,
         \g[16][43] , \g[16][42] , \g[16][41] , \g[16][40] , \g[16][39] ,
         \g[16][38] , \g[16][37] , \g[16][36] , \g[16][35] , \g[16][34] ,
         \g[16][33] , \g[16][32] , \g[16][31] , \g[16][30] , \g[16][29] ,
         \g[16][28] , \g[16][27] , \g[16][26] , \g[16][25] , \g[16][24] ,
         \g[16][23] , \g[16][22] , \g[16][21] , \g[16][20] , \g[16][19] ,
         \g[16][18] , \g[16][17] , \g[16][16] , \g[16][15] , \g[16][14] ,
         \g[16][13] , \g[16][12] , \g[16][11] , \g[16][10] , \g[16][9] ,
         \g[16][8] , \g[16][7] , \g[16][6] , \g[16][5] , \g[16][4] ,
         \g[16][3] , \g[16][2] , \g[16][1] , \g[16][0] , \g[15][63] ,
         \g[15][62] , \g[15][61] , \g[15][60] , \g[15][59] , \g[15][58] ,
         \g[15][57] , \g[15][56] , \g[15][55] , \g[15][54] , \g[15][53] ,
         \g[15][52] , \g[15][51] , \g[15][50] , \g[15][49] , \g[15][48] ,
         \g[15][47] , \g[15][46] , \g[15][45] , \g[15][44] , \g[15][43] ,
         \g[15][42] , \g[15][41] , \g[15][40] , \g[15][39] , \g[15][38] ,
         \g[15][37] , \g[15][36] , \g[15][35] , \g[15][34] , \g[15][33] ,
         \g[15][32] , \g[15][31] , \g[15][30] , \g[15][29] , \g[15][28] ,
         \g[15][27] , \g[15][26] , \g[15][25] , \g[15][24] , \g[15][23] ,
         \g[15][22] , \g[15][21] , \g[15][20] , \g[15][19] , \g[15][18] ,
         \g[15][17] , \g[15][16] , \g[15][15] , \g[15][14] , \g[15][13] ,
         \g[15][12] , \g[15][11] , \g[15][10] , \g[15][9] , \g[15][8] ,
         \g[15][7] , \g[15][6] , \g[15][5] , \g[15][4] , \g[15][3] ,
         \g[15][2] , \g[15][1] , \g[15][0] , \g[14][63] , \g[14][62] ,
         \g[14][61] , \g[14][60] , \g[14][59] , \g[14][58] , \g[14][57] ,
         \g[14][56] , \g[14][55] , \g[14][54] , \g[14][53] , \g[14][52] ,
         \g[14][51] , \g[14][50] , \g[14][49] , \g[14][48] , \g[14][47] ,
         \g[14][46] , \g[14][45] , \g[14][44] , \g[14][43] , \g[14][42] ,
         \g[14][41] , \g[14][40] , \g[14][39] , \g[14][38] , \g[14][37] ,
         \g[14][36] , \g[14][35] , \g[14][34] , \g[14][33] , \g[14][32] ,
         \g[14][31] , \g[14][30] , \g[14][29] , \g[14][28] , \g[14][27] ,
         \g[14][26] , \g[14][25] , \g[14][24] , \g[14][23] , \g[14][22] ,
         \g[14][21] , \g[14][20] , \g[14][19] , \g[14][18] , \g[14][17] ,
         \g[14][16] , \g[14][15] , \g[14][14] , \g[14][13] , \g[14][12] ,
         \g[14][11] , \g[14][10] , \g[14][9] , \g[14][8] , \g[14][7] ,
         \g[14][6] , \g[14][5] , \g[14][4] , \g[14][3] , \g[14][2] ,
         \g[14][1] , \g[14][0] , \g[13][63] , \g[13][62] , \g[13][61] ,
         \g[13][60] , \g[13][59] , \g[13][58] , \g[13][57] , \g[13][56] ,
         \g[13][55] , \g[13][54] , \g[13][53] , \g[13][52] , \g[13][51] ,
         \g[13][50] , \g[13][49] , \g[13][48] , \g[13][47] , \g[13][46] ,
         \g[13][45] , \g[13][44] , \g[13][43] , \g[13][42] , \g[13][41] ,
         \g[13][40] , \g[13][39] , \g[13][38] , \g[13][37] , \g[13][36] ,
         \g[13][35] , \g[13][34] , \g[13][33] , \g[13][32] , \g[13][31] ,
         \g[13][30] , \g[13][29] , \g[13][28] , \g[13][27] , \g[13][26] ,
         \g[13][25] , \g[13][24] , \g[13][23] , \g[13][22] , \g[13][21] ,
         \g[13][20] , \g[13][19] , \g[13][18] , \g[13][17] , \g[13][16] ,
         \g[13][15] , \g[13][14] , \g[13][13] , \g[13][12] , \g[13][11] ,
         \g[13][10] , \g[13][9] , \g[13][8] , \g[13][7] , \g[13][6] ,
         \g[13][5] , \g[13][4] , \g[13][3] , \g[13][2] , \g[13][1] ,
         \g[13][0] , \g[12][63] , \g[12][62] , \g[12][61] , \g[12][60] ,
         \g[12][59] , \g[12][58] , \g[12][57] , \g[12][56] , \g[12][55] ,
         \g[12][54] , \g[12][53] , \g[12][52] , \g[12][51] , \g[12][50] ,
         \g[12][49] , \g[12][48] , \g[12][47] , \g[12][46] , \g[12][45] ,
         \g[12][44] , \g[12][43] , \g[12][42] , \g[12][41] , \g[12][40] ,
         \g[12][39] , \g[12][38] , \g[12][37] , \g[12][36] , \g[12][35] ,
         \g[12][34] , \g[12][33] , \g[12][32] , \g[12][31] , \g[12][30] ,
         \g[12][29] , \g[12][28] , \g[12][27] , \g[12][26] , \g[12][25] ,
         \g[12][24] , \g[12][23] , \g[12][22] , \g[12][21] , \g[12][20] ,
         \g[12][19] , \g[12][18] , \g[12][17] , \g[12][16] , \g[12][15] ,
         \g[12][14] , \g[12][13] , \g[12][12] , \g[12][11] , \g[12][10] ,
         \g[12][9] , \g[12][8] , \g[12][7] , \g[12][6] , \g[12][5] ,
         \g[12][4] , \g[12][3] , \g[12][2] , \g[12][1] , \g[12][0] ,
         \g[11][63] , \g[11][62] , \g[11][61] , \g[11][60] , \g[11][59] ,
         \g[11][58] , \g[11][57] , \g[11][56] , \g[11][55] , \g[11][54] ,
         \g[11][53] , \g[11][52] , \g[11][51] , \g[11][50] , \g[11][49] ,
         \g[11][48] , \g[11][47] , \g[11][46] , \g[11][45] , \g[11][44] ,
         \g[11][43] , \g[11][42] , \g[11][41] , \g[11][40] , \g[11][39] ,
         \g[11][38] , \g[11][37] , \g[11][36] , \g[11][35] , \g[11][34] ,
         \g[11][33] , \g[11][32] , \g[11][31] , \g[11][30] , \g[11][29] ,
         \g[11][28] , \g[11][27] , \g[11][26] , \g[11][25] , \g[11][24] ,
         \g[11][23] , \g[11][22] , \g[11][21] , \g[11][20] , \g[11][19] ,
         \g[11][18] , \g[11][17] , \g[11][16] , \g[11][15] , \g[11][14] ,
         \g[11][13] , \g[11][12] , \g[11][11] , \g[11][10] , \g[11][9] ,
         \g[11][8] , \g[11][7] , \g[11][6] , \g[11][5] , \g[11][4] ,
         \g[11][3] , \g[11][2] , \g[11][1] , \g[11][0] , \g[10][63] ,
         \g[10][62] , \g[10][61] , \g[10][60] , \g[10][59] , \g[10][58] ,
         \g[10][57] , \g[10][56] , \g[10][55] , \g[10][54] , \g[10][53] ,
         \g[10][52] , \g[10][51] , \g[10][50] , \g[10][49] , \g[10][48] ,
         \g[10][47] , \g[10][46] , \g[10][45] , \g[10][44] , \g[10][43] ,
         \g[10][42] , \g[10][41] , \g[10][40] , \g[10][39] , \g[10][38] ,
         \g[10][37] , \g[10][36] , \g[10][35] , \g[10][34] , \g[10][33] ,
         \g[10][32] , \g[10][31] , \g[10][30] , \g[10][29] , \g[10][28] ,
         \g[10][27] , \g[10][26] , \g[10][25] , \g[10][24] , \g[10][23] ,
         \g[10][22] , \g[10][21] , \g[10][20] , \g[10][19] , \g[10][18] ,
         \g[10][17] , \g[10][16] , \g[10][15] , \g[10][14] , \g[10][13] ,
         \g[10][12] , \g[10][11] , \g[10][10] , \g[10][9] , \g[10][8] ,
         \g[10][7] , \g[10][6] , \g[10][5] , \g[10][4] , \g[10][3] ,
         \g[10][2] , \g[10][1] , \g[10][0] , \g[9][63] , \g[9][62] ,
         \g[9][61] , \g[9][60] , \g[9][59] , \g[9][58] , \g[9][57] ,
         \g[9][56] , \g[9][55] , \g[9][54] , \g[9][53] , \g[9][52] ,
         \g[9][51] , \g[9][50] , \g[9][49] , \g[9][48] , \g[9][47] ,
         \g[9][46] , \g[9][45] , \g[9][44] , \g[9][43] , \g[9][42] ,
         \g[9][41] , \g[9][40] , \g[9][39] , \g[9][38] , \g[9][37] ,
         \g[9][36] , \g[9][35] , \g[9][34] , \g[9][33] , \g[9][32] ,
         \g[9][31] , \g[9][30] , \g[9][29] , \g[9][28] , \g[9][27] ,
         \g[9][26] , \g[9][25] , \g[9][24] , \g[9][23] , \g[9][22] ,
         \g[9][21] , \g[9][20] , \g[9][19] , \g[9][18] , \g[9][17] ,
         \g[9][16] , \g[9][15] , \g[9][14] , \g[9][13] , \g[9][12] ,
         \g[9][11] , \g[9][10] , \g[9][9] , \g[9][8] , \g[9][7] , \g[9][6] ,
         \g[9][5] , \g[9][4] , \g[9][3] , \g[9][2] , \g[9][1] , \g[9][0] ,
         \g[8][63] , \g[8][62] , \g[8][61] , \g[8][60] , \g[8][59] ,
         \g[8][58] , \g[8][57] , \g[8][56] , \g[8][55] , \g[8][54] ,
         \g[8][53] , \g[8][52] , \g[8][51] , \g[8][50] , \g[8][49] ,
         \g[8][48] , \g[8][47] , \g[8][46] , \g[8][45] , \g[8][44] ,
         \g[8][43] , \g[8][42] , \g[8][41] , \g[8][40] , \g[8][39] ,
         \g[8][38] , \g[8][37] , \g[8][36] , \g[8][35] , \g[8][34] ,
         \g[8][33] , \g[8][32] , \g[8][31] , \g[8][30] , \g[8][29] ,
         \g[8][28] , \g[8][27] , \g[8][26] , \g[8][25] , \g[8][24] ,
         \g[8][23] , \g[8][22] , \g[8][21] , \g[8][20] , \g[8][19] ,
         \g[8][18] , \g[8][17] , \g[8][16] , \g[8][15] , \g[8][14] ,
         \g[8][13] , \g[8][12] , \g[8][11] , \g[8][10] , \g[8][9] , \g[8][8] ,
         \g[8][7] , \g[8][6] , \g[8][5] , \g[8][4] , \g[8][3] , \g[8][2] ,
         \g[8][1] , \g[8][0] , \g[7][63] , \g[7][62] , \g[7][61] , \g[7][60] ,
         \g[7][59] , \g[7][58] , \g[7][57] , \g[7][56] , \g[7][55] ,
         \g[7][54] , \g[7][53] , \g[7][52] , \g[7][51] , \g[7][50] ,
         \g[7][49] , \g[7][48] , \g[7][47] , \g[7][46] , \g[7][45] ,
         \g[7][44] , \g[7][43] , \g[7][42] , \g[7][41] , \g[7][40] ,
         \g[7][39] , \g[7][38] , \g[7][37] , \g[7][36] , \g[7][35] ,
         \g[7][34] , \g[7][33] , \g[7][32] , \g[7][31] , \g[7][30] ,
         \g[7][29] , \g[7][28] , \g[7][27] , \g[7][26] , \g[7][25] ,
         \g[7][24] , \g[7][23] , \g[7][22] , \g[7][21] , \g[7][20] ,
         \g[7][19] , \g[7][18] , \g[7][17] , \g[7][16] , \g[7][15] ,
         \g[7][14] , \g[7][13] , \g[7][12] , \g[7][11] , \g[7][10] , \g[7][9] ,
         \g[7][8] , \g[7][7] , \g[7][6] , \g[7][5] , \g[7][4] , \g[7][3] ,
         \g[7][2] , \g[7][1] , \g[7][0] , \g[6][63] , \g[6][62] , \g[6][61] ,
         \g[6][60] , \g[6][59] , \g[6][58] , \g[6][57] , \g[6][56] ,
         \g[6][55] , \g[6][54] , \g[6][53] , \g[6][52] , \g[6][51] ,
         \g[6][50] , \g[6][49] , \g[6][48] , \g[6][47] , \g[6][46] ,
         \g[6][45] , \g[6][44] , \g[6][43] , \g[6][42] , \g[6][41] ,
         \g[6][40] , \g[6][39] , \g[6][38] , \g[6][37] , \g[6][36] ,
         \g[6][35] , \g[6][34] , \g[6][33] , \g[6][32] , \g[6][31] ,
         \g[6][30] , \g[6][29] , \g[6][28] , \g[6][27] , \g[6][26] ,
         \g[6][25] , \g[6][24] , \g[6][23] , \g[6][22] , \g[6][21] ,
         \g[6][20] , \g[6][19] , \g[6][18] , \g[6][17] , \g[6][16] ,
         \g[6][15] , \g[6][14] , \g[6][13] , \g[6][12] , \g[6][11] ,
         \g[6][10] , \g[6][9] , \g[6][8] , \g[6][7] , \g[6][6] , \g[6][5] ,
         \g[6][4] , \g[6][3] , \g[6][2] , \g[6][1] , \g[6][0] , \g[5][63] ,
         \g[5][62] , \g[5][61] , \g[5][60] , \g[5][59] , \g[5][58] ,
         \g[5][57] , \g[5][56] , \g[5][55] , \g[5][54] , \g[5][53] ,
         \g[5][52] , \g[5][51] , \g[5][50] , \g[5][49] , \g[5][48] ,
         \g[5][47] , \g[5][46] , \g[5][45] , \g[5][44] , \g[5][43] ,
         \g[5][42] , \g[5][41] , \g[5][40] , \g[5][39] , \g[5][38] ,
         \g[5][37] , \g[5][36] , \g[5][35] , \g[5][34] , \g[5][33] ,
         \g[5][32] , \g[5][31] , \g[5][30] , \g[5][29] , \g[5][28] ,
         \g[5][27] , \g[5][26] , \g[5][25] , \g[5][24] , \g[5][23] ,
         \g[5][22] , \g[5][21] , \g[5][20] , \g[5][19] , \g[5][18] ,
         \g[5][17] , \g[5][16] , \g[5][15] , \g[5][14] , \g[5][13] ,
         \g[5][12] , \g[5][11] , \g[5][10] , \g[5][9] , \g[5][8] , \g[5][7] ,
         \g[5][6] , \g[5][5] , \g[5][4] , \g[5][3] , \g[5][2] , \g[5][1] ,
         \g[5][0] , \g[4][63] , \g[4][62] , \g[4][61] , \g[4][60] , \g[4][59] ,
         \g[4][58] , \g[4][57] , \g[4][56] , \g[4][55] , \g[4][54] ,
         \g[4][53] , \g[4][52] , \g[4][51] , \g[4][50] , \g[4][49] ,
         \g[4][48] , \g[4][47] , \g[4][46] , \g[4][45] , \g[4][44] ,
         \g[4][43] , \g[4][42] , \g[4][41] , \g[4][40] , \g[4][39] ,
         \g[4][38] , \g[4][37] , \g[4][36] , \g[4][35] , \g[4][34] ,
         \g[4][33] , \g[4][32] , \g[4][31] , \g[4][30] , \g[4][29] ,
         \g[4][28] , \g[4][27] , \g[4][26] , \g[4][25] , \g[4][24] ,
         \g[4][23] , \g[4][22] , \g[4][21] , \g[4][20] , \g[4][19] ,
         \g[4][18] , \g[4][17] , \g[4][16] , \g[4][15] , \g[4][14] ,
         \g[4][13] , \g[4][12] , \g[4][11] , \g[4][10] , \g[4][9] , \g[4][8] ,
         \g[4][7] , \g[4][6] , \g[4][5] , \g[4][4] , \g[4][3] , \g[4][2] ,
         \g[4][1] , \g[4][0] , \g[3][63] , \g[3][62] , \g[3][61] , \g[3][60] ,
         \g[3][59] , \g[3][58] , \g[3][57] , \g[3][56] , \g[3][55] ,
         \g[3][54] , \g[3][53] , \g[3][52] , \g[3][51] , \g[3][50] ,
         \g[3][49] , \g[3][48] , \g[3][47] , \g[3][46] , \g[3][45] ,
         \g[3][44] , \g[3][43] , \g[3][42] , \g[3][41] , \g[3][40] ,
         \g[3][39] , \g[3][38] , \g[3][37] , \g[3][36] , \g[3][35] ,
         \g[3][34] , \g[3][33] , \g[3][32] , \g[3][31] , \g[3][30] ,
         \g[3][29] , \g[3][28] , \g[3][27] , \g[3][26] , \g[3][25] ,
         \g[3][24] , \g[3][23] , \g[3][22] , \g[3][21] , \g[3][20] ,
         \g[3][19] , \g[3][18] , \g[3][17] , \g[3][16] , \g[3][15] ,
         \g[3][14] , \g[3][13] , \g[3][12] , \g[3][11] , \g[3][10] , \g[3][9] ,
         \g[3][8] , \g[3][7] , \g[3][6] , \g[3][5] , \g[3][4] , \g[3][3] ,
         \g[3][2] , \g[3][1] , \g[3][0] , \g[2][63] , \g[2][62] , \g[2][61] ,
         \g[2][60] , \g[2][59] , \g[2][58] , \g[2][57] , \g[2][56] ,
         \g[2][55] , \g[2][54] , \g[2][53] , \g[2][52] , \g[2][51] ,
         \g[2][50] , \g[2][49] , \g[2][48] , \g[2][47] , \g[2][46] ,
         \g[2][45] , \g[2][44] , \g[2][43] , \g[2][42] , \g[2][41] ,
         \g[2][40] , \g[2][39] , \g[2][38] , \g[2][37] , \g[2][36] ,
         \g[2][35] , \g[2][34] , \g[2][33] , \g[2][32] , \g[2][31] ,
         \g[2][30] , \g[2][29] , \g[2][28] , \g[2][27] , \g[2][26] ,
         \g[2][25] , \g[2][24] , \g[2][23] , \g[2][22] , \g[2][21] ,
         \g[2][20] , \g[2][19] , \g[2][18] , \g[2][17] , \g[2][16] ,
         \g[2][15] , \g[2][14] , \g[2][13] , \g[2][12] , \g[2][11] ,
         \g[2][10] , \g[2][9] , \g[2][8] , \g[2][7] , \g[2][6] , \g[2][5] ,
         \g[2][4] , \g[2][3] , \g[2][2] , \g[2][1] , \g[2][0] , \g[1][63] ,
         \g[1][62] , \g[1][61] , \g[1][60] , \g[1][59] , \g[1][58] ,
         \g[1][57] , \g[1][56] , \g[1][55] , \g[1][54] , \g[1][53] ,
         \g[1][52] , \g[1][51] , \g[1][50] , \g[1][49] , \g[1][48] ,
         \g[1][47] , \g[1][46] , \g[1][45] , \g[1][44] , \g[1][43] ,
         \g[1][42] , \g[1][41] , \g[1][40] , \g[1][39] , \g[1][38] ,
         \g[1][37] , \g[1][36] , \g[1][35] , \g[1][34] , \g[1][33] ,
         \g[1][32] , \g[1][31] , \g[1][30] , \g[1][29] , \g[1][28] ,
         \g[1][27] , \g[1][26] , \g[1][25] , \g[1][24] , \g[1][23] ,
         \g[1][22] , \g[1][21] , \g[1][20] , \g[1][19] , \g[1][18] ,
         \g[1][17] , \g[1][16] , \g[1][15] , \g[1][14] , \g[1][13] ,
         \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] ,
         \g[1][6] , \g[1][5] , \g[1][4] , \g[1][3] , \g[1][2] , \g[1][1] ,
         \g[1][0] , \g[0][63] , \g[0][62] , \g[0][61] , \g[0][60] , \g[0][59] ,
         \g[0][58] , \g[0][57] , \g[0][56] , \g[0][55] , \g[0][54] ,
         \g[0][53] , \g[0][52] , \g[0][51] , \g[0][50] , \g[0][49] ,
         \g[0][48] , \g[0][47] , \g[0][46] , \g[0][45] , \g[0][44] ,
         \g[0][43] , \g[0][42] , \g[0][41] , \g[0][40] , \g[0][39] ,
         \g[0][38] , \g[0][37] , \g[0][36] , \g[0][35] , \g[0][34] ,
         \g[0][33] , \g[0][32] , \g[0][31] , \g[0][30] , \g[0][29] ,
         \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] , \g[0][24] ,
         \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , \g[0][19] ,
         \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] ,
         \g[0][13] , \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] ,
         \g[0][7] , \g[0][6] , \g[0][5] , \g[0][4] , \g[0][3] , \g[0][2] ,
         \g[0][1] , \g[0][0] , \g2[27][63] , \g2[27][62] , \g2[27][61] ,
         \g2[27][60] , \g2[27][59] , \g2[27][58] , \g2[27][57] , \g2[27][56] ,
         \g2[27][55] , \g2[27][54] , \g2[27][53] , \g2[27][52] , \g2[27][51] ,
         \g2[27][50] , \g2[27][49] , \g2[27][48] , \g2[27][47] , \g2[27][46] ,
         \g2[27][45] , \g2[27][44] , \g2[27][43] , \g2[27][42] , \g2[27][41] ,
         \g2[27][40] , \g2[27][39] , \g2[27][38] , \g2[27][37] , \g2[27][36] ,
         \g2[27][35] , \g2[27][34] , \g2[27][33] , \g2[27][32] , \g2[27][31] ,
         \g2[27][30] , \g2[27][29] , \g2[27][28] , \g2[27][27] , \g2[27][26] ,
         \g2[27][25] , \g2[27][24] , \g2[27][23] , \g2[27][22] , \g2[27][21] ,
         \g2[27][20] , \g2[27][19] , \g2[27][18] , \g2[27][17] , \g2[27][16] ,
         \g2[27][15] , \g2[27][14] , \g2[27][13] , \g2[27][12] , \g2[27][11] ,
         \g2[27][10] , \g2[27][9] , \g2[27][8] , \g2[27][7] , \g2[27][6] ,
         \g2[27][5] , \g2[27][4] , \g2[27][3] , \g2[27][2] , \g2[27][1] ,
         \g2[26][63] , \g2[26][62] , \g2[26][61] , \g2[26][60] , \g2[26][59] ,
         \g2[26][58] , \g2[26][57] , \g2[26][56] , \g2[26][55] , \g2[26][54] ,
         \g2[26][53] , \g2[26][52] , \g2[26][51] , \g2[26][50] , \g2[26][49] ,
         \g2[26][48] , \g2[26][47] , \g2[26][46] , \g2[26][45] , \g2[26][44] ,
         \g2[26][43] , \g2[26][42] , \g2[26][41] , \g2[26][40] , \g2[26][39] ,
         \g2[26][38] , \g2[26][37] , \g2[26][36] , \g2[26][35] , \g2[26][34] ,
         \g2[26][33] , \g2[26][32] , \g2[26][31] , \g2[26][30] , \g2[26][29] ,
         \g2[26][28] , \g2[26][27] , \g2[26][26] , \g2[26][25] , \g2[26][24] ,
         \g2[26][23] , \g2[26][22] , \g2[26][21] , \g2[26][20] , \g2[26][19] ,
         \g2[26][18] , \g2[26][17] , \g2[26][16] , \g2[26][15] , \g2[26][14] ,
         \g2[26][13] , \g2[26][12] , \g2[26][11] , \g2[26][10] , \g2[26][9] ,
         \g2[26][8] , \g2[26][7] , \g2[26][6] , \g2[26][5] , \g2[26][4] ,
         \g2[26][3] , \g2[26][2] , \g2[26][1] , \g2[25][63] , \g2[25][62] ,
         \g2[25][61] , \g2[25][60] , \g2[25][59] , \g2[25][58] , \g2[25][57] ,
         \g2[25][56] , \g2[25][55] , \g2[25][54] , \g2[25][53] , \g2[25][52] ,
         \g2[25][51] , \g2[25][50] , \g2[25][49] , \g2[25][48] , \g2[25][47] ,
         \g2[25][46] , \g2[25][45] , \g2[25][44] , \g2[25][43] , \g2[25][42] ,
         \g2[25][41] , \g2[25][40] , \g2[25][39] , \g2[25][38] , \g2[25][37] ,
         \g2[25][36] , \g2[25][35] , \g2[25][34] , \g2[25][33] , \g2[25][32] ,
         \g2[25][31] , \g2[25][30] , \g2[25][29] , \g2[25][28] , \g2[25][27] ,
         \g2[25][26] , \g2[25][25] , \g2[25][24] , \g2[25][23] , \g2[25][22] ,
         \g2[25][21] , \g2[25][20] , \g2[25][19] , \g2[25][18] , \g2[25][17] ,
         \g2[25][16] , \g2[25][15] , \g2[25][14] , \g2[25][13] , \g2[25][12] ,
         \g2[25][11] , \g2[25][10] , \g2[25][9] , \g2[25][8] , \g2[25][7] ,
         \g2[25][6] , \g2[25][5] , \g2[25][4] , \g2[25][3] , \g2[25][2] ,
         \g2[25][1] , \g2[24][63] , \g2[24][62] , \g2[24][61] , \g2[24][60] ,
         \g2[24][59] , \g2[24][58] , \g2[24][57] , \g2[24][56] , \g2[24][55] ,
         \g2[24][54] , \g2[24][53] , \g2[24][52] , \g2[24][51] , \g2[24][50] ,
         \g2[24][49] , \g2[24][48] , \g2[24][47] , \g2[24][46] , \g2[24][45] ,
         \g2[24][44] , \g2[24][43] , \g2[24][42] , \g2[24][41] , \g2[24][40] ,
         \g2[24][39] , \g2[24][38] , \g2[24][37] , \g2[24][36] , \g2[24][35] ,
         \g2[24][34] , \g2[24][33] , \g2[24][32] , \g2[24][31] , \g2[24][30] ,
         \g2[24][29] , \g2[24][28] , \g2[24][27] , \g2[24][26] , \g2[24][25] ,
         \g2[24][24] , \g2[24][23] , \g2[24][22] , \g2[24][21] , \g2[24][20] ,
         \g2[24][19] , \g2[24][18] , \g2[24][17] , \g2[24][16] , \g2[24][15] ,
         \g2[24][14] , \g2[24][13] , \g2[24][12] , \g2[24][11] , \g2[24][10] ,
         \g2[24][9] , \g2[24][8] , \g2[24][7] , \g2[24][6] , \g2[24][5] ,
         \g2[24][4] , \g2[24][3] , \g2[24][2] , \g2[24][1] , \g2[23][63] ,
         \g2[23][62] , \g2[23][61] , \g2[23][60] , \g2[23][59] , \g2[23][58] ,
         \g2[23][57] , \g2[23][56] , \g2[23][55] , \g2[23][54] , \g2[23][53] ,
         \g2[23][52] , \g2[23][51] , \g2[23][50] , \g2[23][49] , \g2[23][48] ,
         \g2[23][47] , \g2[23][46] , \g2[23][45] , \g2[23][44] , \g2[23][43] ,
         \g2[23][42] , \g2[23][41] , \g2[23][40] , \g2[23][39] , \g2[23][38] ,
         \g2[23][37] , \g2[23][36] , \g2[23][35] , \g2[23][34] , \g2[23][33] ,
         \g2[23][32] , \g2[23][31] , \g2[23][30] , \g2[23][29] , \g2[23][28] ,
         \g2[23][27] , \g2[23][26] , \g2[23][25] , \g2[23][24] , \g2[23][23] ,
         \g2[23][22] , \g2[23][21] , \g2[23][20] , \g2[23][19] , \g2[23][18] ,
         \g2[23][17] , \g2[23][16] , \g2[23][15] , \g2[23][14] , \g2[23][13] ,
         \g2[23][12] , \g2[23][11] , \g2[23][10] , \g2[23][9] , \g2[23][8] ,
         \g2[23][7] , \g2[23][6] , \g2[23][5] , \g2[23][4] , \g2[23][3] ,
         \g2[23][2] , \g2[23][1] , \g2[22][63] , \g2[22][62] , \g2[22][61] ,
         \g2[22][60] , \g2[22][59] , \g2[22][58] , \g2[22][57] , \g2[22][56] ,
         \g2[22][55] , \g2[22][54] , \g2[22][53] , \g2[22][52] , \g2[22][51] ,
         \g2[22][50] , \g2[22][49] , \g2[22][48] , \g2[22][47] , \g2[22][46] ,
         \g2[22][45] , \g2[22][44] , \g2[22][43] , \g2[22][42] , \g2[22][41] ,
         \g2[22][40] , \g2[22][39] , \g2[22][38] , \g2[22][37] , \g2[22][36] ,
         \g2[22][35] , \g2[22][34] , \g2[22][33] , \g2[22][32] , \g2[22][31] ,
         \g2[22][30] , \g2[22][29] , \g2[22][28] , \g2[22][27] , \g2[22][26] ,
         \g2[22][25] , \g2[22][24] , \g2[22][23] , \g2[22][22] , \g2[22][21] ,
         \g2[22][20] , \g2[22][19] , \g2[22][18] , \g2[22][17] , \g2[22][16] ,
         \g2[22][15] , \g2[22][14] , \g2[22][13] , \g2[22][12] , \g2[22][11] ,
         \g2[22][10] , \g2[22][9] , \g2[22][8] , \g2[22][7] , \g2[22][6] ,
         \g2[22][5] , \g2[22][4] , \g2[22][3] , \g2[22][2] , \g2[22][1] ,
         \g2[21][63] , \g2[21][62] , \g2[21][61] , \g2[21][60] , \g2[21][59] ,
         \g2[21][58] , \g2[21][57] , \g2[21][56] , \g2[21][55] , \g2[21][54] ,
         \g2[21][53] , \g2[21][52] , \g2[21][51] , \g2[21][50] , \g2[21][49] ,
         \g2[21][48] , \g2[21][47] , \g2[21][46] , \g2[21][45] , \g2[21][44] ,
         \g2[21][43] , \g2[21][42] , \g2[21][41] , \g2[21][40] , \g2[21][39] ,
         \g2[21][38] , \g2[21][37] , \g2[21][36] , \g2[21][35] , \g2[21][34] ,
         \g2[21][33] , \g2[21][32] , \g2[21][31] , \g2[21][30] , \g2[21][29] ,
         \g2[21][28] , \g2[21][27] , \g2[21][26] , \g2[21][25] , \g2[21][24] ,
         \g2[21][23] , \g2[21][22] , \g2[21][21] , \g2[21][20] , \g2[21][19] ,
         \g2[21][18] , \g2[21][17] , \g2[21][16] , \g2[21][15] , \g2[21][14] ,
         \g2[21][13] , \g2[21][12] , \g2[21][11] , \g2[21][10] , \g2[21][9] ,
         \g2[21][8] , \g2[21][7] , \g2[21][6] , \g2[21][5] , \g2[21][4] ,
         \g2[21][3] , \g2[21][2] , \g2[21][1] , \g2[20][63] , \g2[20][62] ,
         \g2[20][61] , \g2[20][60] , \g2[20][59] , \g2[20][58] , \g2[20][57] ,
         \g2[20][56] , \g2[20][55] , \g2[20][54] , \g2[20][53] , \g2[20][52] ,
         \g2[20][51] , \g2[20][50] , \g2[20][49] , \g2[20][48] , \g2[20][47] ,
         \g2[20][46] , \g2[20][45] , \g2[20][44] , \g2[20][43] , \g2[20][42] ,
         \g2[20][41] , \g2[20][40] , \g2[20][39] , \g2[20][38] , \g2[20][37] ,
         \g2[20][36] , \g2[20][35] , \g2[20][34] , \g2[20][33] , \g2[20][32] ,
         \g2[20][31] , \g2[20][30] , \g2[20][29] , \g2[20][28] , \g2[20][27] ,
         \g2[20][26] , \g2[20][25] , \g2[20][24] , \g2[20][23] , \g2[20][22] ,
         \g2[20][21] , \g2[20][20] , \g2[20][19] , \g2[20][18] , \g2[20][17] ,
         \g2[20][16] , \g2[20][15] , \g2[20][14] , \g2[20][13] , \g2[20][12] ,
         \g2[20][11] , \g2[20][10] , \g2[20][9] , \g2[20][8] , \g2[20][7] ,
         \g2[20][6] , \g2[20][5] , \g2[20][4] , \g2[20][3] , \g2[20][2] ,
         \g2[20][1] , \g2[19][63] , \g2[19][62] , \g2[19][61] , \g2[19][60] ,
         \g2[19][59] , \g2[19][58] , \g2[19][57] , \g2[19][56] , \g2[19][55] ,
         \g2[19][54] , \g2[19][53] , \g2[19][52] , \g2[19][51] , \g2[19][50] ,
         \g2[19][49] , \g2[19][48] , \g2[19][47] , \g2[19][46] , \g2[19][45] ,
         \g2[19][44] , \g2[19][43] , \g2[19][42] , \g2[19][41] , \g2[19][40] ,
         \g2[19][39] , \g2[19][38] , \g2[19][37] , \g2[19][36] , \g2[19][35] ,
         \g2[19][34] , \g2[19][33] , \g2[19][32] , \g2[19][31] , \g2[19][30] ,
         \g2[19][29] , \g2[19][28] , \g2[19][27] , \g2[19][26] , \g2[19][25] ,
         \g2[19][24] , \g2[19][23] , \g2[19][22] , \g2[19][21] , \g2[19][20] ,
         \g2[19][19] , \g2[19][18] , \g2[19][17] , \g2[19][16] , \g2[19][15] ,
         \g2[19][14] , \g2[19][13] , \g2[19][12] , \g2[19][11] , \g2[19][10] ,
         \g2[19][9] , \g2[19][8] , \g2[19][7] , \g2[19][6] , \g2[19][5] ,
         \g2[19][4] , \g2[19][3] , \g2[19][2] , \g2[19][1] , \g2[18][63] ,
         \g2[18][62] , \g2[18][61] , \g2[18][60] , \g2[18][59] , \g2[18][58] ,
         \g2[18][57] , \g2[18][56] , \g2[18][55] , \g2[18][54] , \g2[18][53] ,
         \g2[18][52] , \g2[18][51] , \g2[18][50] , \g2[18][49] , \g2[18][48] ,
         \g2[18][47] , \g2[18][46] , \g2[18][45] , \g2[18][44] , \g2[18][43] ,
         \g2[18][42] , \g2[18][41] , \g2[18][40] , \g2[18][39] , \g2[18][38] ,
         \g2[18][37] , \g2[18][36] , \g2[18][35] , \g2[18][34] , \g2[18][33] ,
         \g2[18][32] , \g2[18][31] , \g2[18][30] , \g2[18][29] , \g2[18][28] ,
         \g2[18][27] , \g2[18][26] , \g2[18][25] , \g2[18][24] , \g2[18][23] ,
         \g2[18][22] , \g2[18][21] , \g2[18][20] , \g2[18][19] , \g2[18][18] ,
         \g2[18][17] , \g2[18][16] , \g2[18][15] , \g2[18][14] , \g2[18][13] ,
         \g2[18][12] , \g2[18][11] , \g2[18][10] , \g2[18][9] , \g2[18][8] ,
         \g2[18][7] , \g2[18][6] , \g2[18][5] , \g2[18][4] , \g2[18][3] ,
         \g2[18][2] , \g2[18][1] , \g2[17][63] , \g2[17][62] , \g2[17][61] ,
         \g2[17][60] , \g2[17][59] , \g2[17][58] , \g2[17][57] , \g2[17][56] ,
         \g2[17][55] , \g2[17][54] , \g2[17][53] , \g2[17][52] , \g2[17][51] ,
         \g2[17][50] , \g2[17][49] , \g2[17][48] , \g2[17][47] , \g2[17][46] ,
         \g2[17][45] , \g2[17][44] , \g2[17][43] , \g2[17][42] , \g2[17][41] ,
         \g2[17][40] , \g2[17][39] , \g2[17][38] , \g2[17][37] , \g2[17][36] ,
         \g2[17][35] , \g2[17][34] , \g2[17][33] , \g2[17][32] , \g2[17][31] ,
         \g2[17][30] , \g2[17][29] , \g2[17][28] , \g2[17][27] , \g2[17][26] ,
         \g2[17][25] , \g2[17][24] , \g2[17][23] , \g2[17][22] , \g2[17][21] ,
         \g2[17][20] , \g2[17][19] , \g2[17][18] , \g2[17][17] , \g2[17][16] ,
         \g2[17][15] , \g2[17][14] , \g2[17][13] , \g2[17][12] , \g2[17][11] ,
         \g2[17][10] , \g2[17][9] , \g2[17][8] , \g2[17][7] , \g2[17][6] ,
         \g2[17][5] , \g2[17][4] , \g2[17][3] , \g2[17][2] , \g2[17][1] ,
         \g2[16][63] , \g2[16][62] , \g2[16][61] , \g2[16][60] , \g2[16][59] ,
         \g2[16][58] , \g2[16][57] , \g2[16][56] , \g2[16][55] , \g2[16][54] ,
         \g2[16][53] , \g2[16][52] , \g2[16][51] , \g2[16][50] , \g2[16][49] ,
         \g2[16][48] , \g2[16][47] , \g2[16][46] , \g2[16][45] , \g2[16][44] ,
         \g2[16][43] , \g2[16][42] , \g2[16][41] , \g2[16][40] , \g2[16][39] ,
         \g2[16][38] , \g2[16][37] , \g2[16][36] , \g2[16][35] , \g2[16][34] ,
         \g2[16][33] , \g2[16][32] , \g2[16][31] , \g2[16][30] , \g2[16][29] ,
         \g2[16][28] , \g2[16][27] , \g2[16][26] , \g2[16][25] , \g2[16][24] ,
         \g2[16][23] , \g2[16][22] , \g2[16][21] , \g2[16][20] , \g2[16][19] ,
         \g2[16][18] , \g2[16][17] , \g2[16][16] , \g2[16][15] , \g2[16][14] ,
         \g2[16][13] , \g2[16][12] , \g2[16][11] , \g2[16][10] , \g2[16][9] ,
         \g2[16][8] , \g2[16][7] , \g2[16][6] , \g2[16][5] , \g2[16][4] ,
         \g2[16][3] , \g2[16][2] , \g2[16][1] , \g2[15][63] , \g2[15][62] ,
         \g2[15][61] , \g2[15][60] , \g2[15][59] , \g2[15][58] , \g2[15][57] ,
         \g2[15][56] , \g2[15][55] , \g2[15][54] , \g2[15][53] , \g2[15][52] ,
         \g2[15][51] , \g2[15][50] , \g2[15][49] , \g2[15][48] , \g2[15][47] ,
         \g2[15][46] , \g2[15][45] , \g2[15][44] , \g2[15][43] , \g2[15][42] ,
         \g2[15][41] , \g2[15][40] , \g2[15][39] , \g2[15][38] , \g2[15][37] ,
         \g2[15][36] , \g2[15][35] , \g2[15][34] , \g2[15][33] , \g2[15][32] ,
         \g2[15][31] , \g2[15][30] , \g2[15][29] , \g2[15][28] , \g2[15][27] ,
         \g2[15][26] , \g2[15][25] , \g2[15][24] , \g2[15][23] , \g2[15][22] ,
         \g2[15][21] , \g2[15][20] , \g2[15][19] , \g2[15][18] , \g2[15][17] ,
         \g2[15][16] , \g2[15][15] , \g2[15][14] , \g2[15][13] , \g2[15][12] ,
         \g2[15][11] , \g2[15][10] , \g2[15][9] , \g2[15][8] , \g2[15][7] ,
         \g2[15][6] , \g2[15][5] , \g2[15][4] , \g2[15][3] , \g2[15][2] ,
         \g2[15][1] , \g2[14][63] , \g2[14][62] , \g2[14][61] , \g2[14][60] ,
         \g2[14][59] , \g2[14][58] , \g2[14][57] , \g2[14][56] , \g2[14][55] ,
         \g2[14][54] , \g2[14][53] , \g2[14][52] , \g2[14][51] , \g2[14][50] ,
         \g2[14][49] , \g2[14][48] , \g2[14][47] , \g2[14][46] , \g2[14][45] ,
         \g2[14][44] , \g2[14][43] , \g2[14][42] , \g2[14][41] , \g2[14][40] ,
         \g2[14][39] , \g2[14][38] , \g2[14][37] , \g2[14][36] , \g2[14][35] ,
         \g2[14][34] , \g2[14][33] , \g2[14][32] , \g2[14][31] , \g2[14][30] ,
         \g2[14][29] , \g2[14][28] , \g2[14][27] , \g2[14][26] , \g2[14][25] ,
         \g2[14][24] , \g2[14][23] , \g2[14][22] , \g2[14][21] , \g2[14][20] ,
         \g2[14][19] , \g2[14][18] , \g2[14][17] , \g2[14][16] , \g2[14][15] ,
         \g2[14][14] , \g2[14][13] , \g2[14][12] , \g2[14][11] , \g2[14][10] ,
         \g2[14][9] , \g2[14][8] , \g2[14][7] , \g2[14][6] , \g2[14][5] ,
         \g2[14][4] , \g2[14][3] , \g2[14][2] , \g2[14][1] , \g2[13][63] ,
         \g2[13][62] , \g2[13][61] , \g2[13][60] , \g2[13][59] , \g2[13][58] ,
         \g2[13][57] , \g2[13][56] , \g2[13][55] , \g2[13][54] , \g2[13][53] ,
         \g2[13][52] , \g2[13][51] , \g2[13][50] , \g2[13][49] , \g2[13][48] ,
         \g2[13][47] , \g2[13][46] , \g2[13][45] , \g2[13][44] , \g2[13][43] ,
         \g2[13][42] , \g2[13][41] , \g2[13][40] , \g2[13][39] , \g2[13][38] ,
         \g2[13][37] , \g2[13][36] , \g2[13][35] , \g2[13][34] , \g2[13][33] ,
         \g2[13][32] , \g2[13][31] , \g2[13][30] , \g2[13][29] , \g2[13][28] ,
         \g2[13][27] , \g2[13][26] , \g2[13][25] , \g2[13][24] , \g2[13][23] ,
         \g2[13][22] , \g2[13][21] , \g2[13][20] , \g2[13][19] , \g2[13][18] ,
         \g2[13][17] , \g2[13][16] , \g2[13][15] , \g2[13][14] , \g2[13][13] ,
         \g2[13][12] , \g2[13][11] , \g2[13][10] , \g2[13][9] , \g2[13][8] ,
         \g2[13][7] , \g2[13][6] , \g2[13][5] , \g2[13][4] , \g2[13][3] ,
         \g2[13][2] , \g2[13][1] , \g2[13][0] , \g2[12][63] , \g2[12][62] ,
         \g2[12][61] , \g2[12][60] , \g2[12][59] , \g2[12][58] , \g2[12][57] ,
         \g2[12][56] , \g2[12][55] , \g2[12][54] , \g2[12][53] , \g2[12][52] ,
         \g2[12][51] , \g2[12][50] , \g2[12][49] , \g2[12][48] , \g2[12][47] ,
         \g2[12][46] , \g2[12][45] , \g2[12][44] , \g2[12][43] , \g2[12][42] ,
         \g2[12][41] , \g2[12][40] , \g2[12][39] , \g2[12][38] , \g2[12][37] ,
         \g2[12][36] , \g2[12][35] , \g2[12][34] , \g2[12][33] , \g2[12][32] ,
         \g2[12][31] , \g2[12][30] , \g2[12][29] , \g2[12][28] , \g2[12][27] ,
         \g2[12][26] , \g2[12][25] , \g2[12][24] , \g2[12][23] , \g2[12][22] ,
         \g2[12][21] , \g2[12][20] , \g2[12][19] , \g2[12][18] , \g2[12][17] ,
         \g2[12][16] , \g2[12][15] , \g2[12][14] , \g2[12][13] , \g2[12][12] ,
         \g2[12][11] , \g2[12][10] , \g2[12][9] , \g2[12][8] , \g2[12][7] ,
         \g2[12][6] , \g2[12][5] , \g2[12][4] , \g2[12][3] , \g2[12][2] ,
         \g2[12][1] , \g2[12][0] , \g2[11][63] , \g2[11][62] , \g2[11][61] ,
         \g2[11][60] , \g2[11][59] , \g2[11][58] , \g2[11][57] , \g2[11][56] ,
         \g2[11][55] , \g2[11][54] , \g2[11][53] , \g2[11][52] , \g2[11][51] ,
         \g2[11][50] , \g2[11][49] , \g2[11][48] , \g2[11][47] , \g2[11][46] ,
         \g2[11][45] , \g2[11][44] , \g2[11][43] , \g2[11][42] , \g2[11][41] ,
         \g2[11][40] , \g2[11][39] , \g2[11][38] , \g2[11][37] , \g2[11][36] ,
         \g2[11][35] , \g2[11][34] , \g2[11][33] , \g2[11][32] , \g2[11][31] ,
         \g2[11][30] , \g2[11][29] , \g2[11][28] , \g2[11][27] , \g2[11][26] ,
         \g2[11][25] , \g2[11][24] , \g2[11][23] , \g2[11][22] , \g2[11][21] ,
         \g2[11][20] , \g2[11][19] , \g2[11][18] , \g2[11][17] , \g2[11][16] ,
         \g2[11][15] , \g2[11][14] , \g2[11][13] , \g2[11][12] , \g2[11][11] ,
         \g2[11][10] , \g2[11][9] , \g2[11][8] , \g2[11][7] , \g2[11][6] ,
         \g2[11][5] , \g2[11][4] , \g2[11][3] , \g2[11][2] , \g2[11][1] ,
         \g2[11][0] , \g2[10][63] , \g2[10][62] , \g2[10][61] , \g2[10][60] ,
         \g2[10][59] , \g2[10][58] , \g2[10][57] , \g2[10][56] , \g2[10][55] ,
         \g2[10][54] , \g2[10][53] , \g2[10][52] , \g2[10][51] , \g2[10][50] ,
         \g2[10][49] , \g2[10][48] , \g2[10][47] , \g2[10][46] , \g2[10][45] ,
         \g2[10][44] , \g2[10][43] , \g2[10][42] , \g2[10][41] , \g2[10][40] ,
         \g2[10][39] , \g2[10][38] , \g2[10][37] , \g2[10][36] , \g2[10][35] ,
         \g2[10][34] , \g2[10][33] , \g2[10][32] , \g2[10][31] , \g2[10][30] ,
         \g2[10][29] , \g2[10][28] , \g2[10][27] , \g2[10][26] , \g2[10][25] ,
         \g2[10][24] , \g2[10][23] , \g2[10][22] , \g2[10][21] , \g2[10][20] ,
         \g2[10][19] , \g2[10][18] , \g2[10][17] , \g2[10][16] , \g2[10][15] ,
         \g2[10][14] , \g2[10][13] , \g2[10][12] , \g2[10][11] , \g2[10][10] ,
         \g2[10][9] , \g2[10][8] , \g2[10][7] , \g2[10][6] , \g2[10][5] ,
         \g2[10][4] , \g2[10][3] , \g2[10][2] , \g2[10][1] , \g2[10][0] ,
         \g2[9][63] , \g2[9][62] , \g2[9][61] , \g2[9][60] , \g2[9][59] ,
         \g2[9][58] , \g2[9][57] , \g2[9][56] , \g2[9][55] , \g2[9][54] ,
         \g2[9][53] , \g2[9][52] , \g2[9][51] , \g2[9][50] , \g2[9][49] ,
         \g2[9][48] , \g2[9][47] , \g2[9][46] , \g2[9][45] , \g2[9][44] ,
         \g2[9][43] , \g2[9][42] , \g2[9][41] , \g2[9][40] , \g2[9][39] ,
         \g2[9][38] , \g2[9][37] , \g2[9][36] , \g2[9][35] , \g2[9][34] ,
         \g2[9][33] , \g2[9][32] , \g2[9][31] , \g2[9][30] , \g2[9][29] ,
         \g2[9][28] , \g2[9][27] , \g2[9][26] , \g2[9][25] , \g2[9][24] ,
         \g2[9][23] , \g2[9][22] , \g2[9][21] , \g2[9][20] , \g2[9][19] ,
         \g2[9][18] , \g2[9][17] , \g2[9][16] , \g2[9][15] , \g2[9][14] ,
         \g2[9][13] , \g2[9][12] , \g2[9][11] , \g2[9][10] , \g2[9][9] ,
         \g2[9][8] , \g2[9][7] , \g2[9][6] , \g2[9][5] , \g2[9][4] ,
         \g2[9][3] , \g2[9][2] , \g2[9][1] , \g2[9][0] , \g2[8][63] ,
         \g2[8][62] , \g2[8][61] , \g2[8][60] , \g2[8][59] , \g2[8][58] ,
         \g2[8][57] , \g2[8][56] , \g2[8][55] , \g2[8][54] , \g2[8][53] ,
         \g2[8][52] , \g2[8][51] , \g2[8][50] , \g2[8][49] , \g2[8][48] ,
         \g2[8][47] , \g2[8][46] , \g2[8][45] , \g2[8][44] , \g2[8][43] ,
         \g2[8][42] , \g2[8][41] , \g2[8][40] , \g2[8][39] , \g2[8][38] ,
         \g2[8][37] , \g2[8][36] , \g2[8][35] , \g2[8][34] , \g2[8][33] ,
         \g2[8][32] , \g2[8][31] , \g2[8][30] , \g2[8][29] , \g2[8][28] ,
         \g2[8][27] , \g2[8][26] , \g2[8][25] , \g2[8][24] , \g2[8][23] ,
         \g2[8][22] , \g2[8][21] , \g2[8][20] , \g2[8][19] , \g2[8][18] ,
         \g2[8][17] , \g2[8][16] , \g2[8][15] , \g2[8][14] , \g2[8][13] ,
         \g2[8][12] , \g2[8][11] , \g2[8][10] , \g2[8][9] , \g2[8][8] ,
         \g2[8][7] , \g2[8][6] , \g2[8][5] , \g2[8][4] , \g2[8][3] ,
         \g2[8][2] , \g2[8][1] , \g2[8][0] , \g2[7][63] , \g2[7][62] ,
         \g2[7][61] , \g2[7][60] , \g2[7][59] , \g2[7][58] , \g2[7][57] ,
         \g2[7][56] , \g2[7][55] , \g2[7][54] , \g2[7][53] , \g2[7][52] ,
         \g2[7][51] , \g2[7][50] , \g2[7][49] , \g2[7][48] , \g2[7][47] ,
         \g2[7][46] , \g2[7][45] , \g2[7][44] , \g2[7][43] , \g2[7][42] ,
         \g2[7][41] , \g2[7][40] , \g2[7][39] , \g2[7][38] , \g2[7][37] ,
         \g2[7][36] , \g2[7][35] , \g2[7][34] , \g2[7][33] , \g2[7][32] ,
         \g2[7][31] , \g2[7][30] , \g2[7][29] , \g2[7][28] , \g2[7][27] ,
         \g2[7][26] , \g2[7][25] , \g2[7][24] , \g2[7][23] , \g2[7][22] ,
         \g2[7][21] , \g2[7][20] , \g2[7][19] , \g2[7][18] , \g2[7][17] ,
         \g2[7][16] , \g2[7][15] , \g2[7][14] , \g2[7][13] , \g2[7][12] ,
         \g2[7][11] , \g2[7][10] , \g2[7][9] , \g2[7][8] , \g2[7][7] ,
         \g2[7][6] , \g2[7][5] , \g2[7][4] , \g2[7][3] , \g2[7][2] ,
         \g2[7][1] , \g2[7][0] , \g2[6][63] , \g2[6][62] , \g2[6][61] ,
         \g2[6][60] , \g2[6][59] , \g2[6][58] , \g2[6][57] , \g2[6][56] ,
         \g2[6][55] , \g2[6][54] , \g2[6][53] , \g2[6][52] , \g2[6][51] ,
         \g2[6][50] , \g2[6][49] , \g2[6][48] , \g2[6][47] , \g2[6][46] ,
         \g2[6][45] , \g2[6][44] , \g2[6][43] , \g2[6][42] , \g2[6][41] ,
         \g2[6][40] , \g2[6][39] , \g2[6][38] , \g2[6][37] , \g2[6][36] ,
         \g2[6][35] , \g2[6][34] , \g2[6][33] , \g2[6][32] , \g2[6][31] ,
         \g2[6][30] , \g2[6][29] , \g2[6][28] , \g2[6][27] , \g2[6][26] ,
         \g2[6][25] , \g2[6][24] , \g2[6][23] , \g2[6][22] , \g2[6][21] ,
         \g2[6][20] , \g2[6][19] , \g2[6][18] , \g2[6][17] , \g2[6][16] ,
         \g2[6][15] , \g2[6][14] , \g2[6][13] , \g2[6][12] , \g2[6][11] ,
         \g2[6][10] , \g2[6][9] , \g2[6][8] , \g2[6][7] , \g2[6][6] ,
         \g2[6][5] , \g2[6][4] , \g2[6][3] , \g2[6][2] , \g2[6][1] ,
         \g2[6][0] , \g2[5][63] , \g2[5][62] , \g2[5][61] , \g2[5][60] ,
         \g2[5][59] , \g2[5][58] , \g2[5][57] , \g2[5][56] , \g2[5][55] ,
         \g2[5][54] , \g2[5][53] , \g2[5][52] , \g2[5][51] , \g2[5][50] ,
         \g2[5][49] , \g2[5][48] , \g2[5][47] , \g2[5][46] , \g2[5][45] ,
         \g2[5][44] , \g2[5][43] , \g2[5][42] , \g2[5][41] , \g2[5][40] ,
         \g2[5][39] , \g2[5][38] , \g2[5][37] , \g2[5][36] , \g2[5][35] ,
         \g2[5][34] , \g2[5][33] , \g2[5][32] , \g2[5][31] , \g2[5][30] ,
         \g2[5][29] , \g2[5][28] , \g2[5][27] , \g2[5][26] , \g2[5][25] ,
         \g2[5][24] , \g2[5][23] , \g2[5][22] , \g2[5][21] , \g2[5][20] ,
         \g2[5][19] , \g2[5][18] , \g2[5][17] , \g2[5][16] , \g2[5][15] ,
         \g2[5][14] , \g2[5][13] , \g2[5][12] , \g2[5][11] , \g2[5][10] ,
         \g2[5][9] , \g2[5][8] , \g2[5][7] , \g2[5][6] , \g2[5][5] ,
         \g2[5][4] , \g2[5][3] , \g2[5][2] , \g2[5][1] , \g2[5][0] ,
         \g2[4][63] , \g2[4][62] , \g2[4][61] , \g2[4][60] , \g2[4][59] ,
         \g2[4][58] , \g2[4][57] , \g2[4][56] , \g2[4][55] , \g2[4][54] ,
         \g2[4][53] , \g2[4][52] , \g2[4][51] , \g2[4][50] , \g2[4][49] ,
         \g2[4][48] , \g2[4][47] , \g2[4][46] , \g2[4][45] , \g2[4][44] ,
         \g2[4][43] , \g2[4][42] , \g2[4][41] , \g2[4][40] , \g2[4][39] ,
         \g2[4][38] , \g2[4][37] , \g2[4][36] , \g2[4][35] , \g2[4][34] ,
         \g2[4][33] , \g2[4][32] , \g2[4][31] , \g2[4][30] , \g2[4][29] ,
         \g2[4][28] , \g2[4][27] , \g2[4][26] , \g2[4][25] , \g2[4][24] ,
         \g2[4][23] , \g2[4][22] , \g2[4][21] , \g2[4][20] , \g2[4][19] ,
         \g2[4][18] , \g2[4][17] , \g2[4][16] , \g2[4][15] , \g2[4][14] ,
         \g2[4][13] , \g2[4][12] , \g2[4][11] , \g2[4][10] , \g2[4][9] ,
         \g2[4][8] , \g2[4][7] , \g2[4][6] , \g2[4][5] , \g2[4][4] ,
         \g2[4][3] , \g2[4][2] , \g2[4][1] , \g2[4][0] , \g2[3][63] ,
         \g2[3][62] , \g2[3][61] , \g2[3][60] , \g2[3][59] , \g2[3][58] ,
         \g2[3][57] , \g2[3][56] , \g2[3][55] , \g2[3][54] , \g2[3][53] ,
         \g2[3][52] , \g2[3][51] , \g2[3][50] , \g2[3][49] , \g2[3][48] ,
         \g2[3][47] , \g2[3][46] , \g2[3][45] , \g2[3][44] , \g2[3][43] ,
         \g2[3][42] , \g2[3][41] , \g2[3][40] , \g2[3][39] , \g2[3][38] ,
         \g2[3][37] , \g2[3][36] , \g2[3][35] , \g2[3][34] , \g2[3][33] ,
         \g2[3][32] , \g2[3][31] , \g2[3][30] , \g2[3][29] , \g2[3][28] ,
         \g2[3][27] , \g2[3][26] , \g2[3][25] , \g2[3][24] , \g2[3][23] ,
         \g2[3][22] , \g2[3][21] , \g2[3][20] , \g2[3][19] , \g2[3][18] ,
         \g2[3][17] , \g2[3][16] , \g2[3][15] , \g2[3][14] , \g2[3][13] ,
         \g2[3][12] , \g2[3][11] , \g2[3][10] , \g2[3][9] , \g2[3][8] ,
         \g2[3][7] , \g2[3][6] , \g2[3][5] , \g2[3][4] , \g2[3][3] ,
         \g2[3][2] , \g2[3][1] , \g2[3][0] , \g2[2][63] , \g2[2][62] ,
         \g2[2][61] , \g2[2][60] , \g2[2][59] , \g2[2][58] , \g2[2][57] ,
         \g2[2][56] , \g2[2][55] , \g2[2][54] , \g2[2][53] , \g2[2][52] ,
         \g2[2][51] , \g2[2][50] , \g2[2][49] , \g2[2][48] , \g2[2][47] ,
         \g2[2][46] , \g2[2][45] , \g2[2][44] , \g2[2][43] , \g2[2][42] ,
         \g2[2][41] , \g2[2][40] , \g2[2][39] , \g2[2][38] , \g2[2][37] ,
         \g2[2][36] , \g2[2][35] , \g2[2][34] , \g2[2][33] , \g2[2][32] ,
         \g2[2][31] , \g2[2][30] , \g2[2][29] , \g2[2][28] , \g2[2][27] ,
         \g2[2][26] , \g2[2][25] , \g2[2][24] , \g2[2][23] , \g2[2][22] ,
         \g2[2][21] , \g2[2][20] , \g2[2][19] , \g2[2][18] , \g2[2][17] ,
         \g2[2][16] , \g2[2][15] , \g2[2][14] , \g2[2][13] , \g2[2][12] ,
         \g2[2][11] , \g2[2][10] , \g2[2][9] , \g2[2][8] , \g2[2][7] ,
         \g2[2][6] , \g2[2][5] , \g2[2][4] , \g2[2][3] , \g2[2][2] ,
         \g2[2][1] , \g2[2][0] , \g2[1][63] , \g2[1][62] , \g2[1][61] ,
         \g2[1][60] , \g2[1][59] , \g2[1][58] , \g2[1][57] , \g2[1][56] ,
         \g2[1][55] , \g2[1][54] , \g2[1][53] , \g2[1][52] , \g2[1][51] ,
         \g2[1][50] , \g2[1][49] , \g2[1][48] , \g2[1][47] , \g2[1][46] ,
         \g2[1][45] , \g2[1][44] , \g2[1][43] , \g2[1][42] , \g2[1][41] ,
         \g2[1][40] , \g2[1][39] , \g2[1][38] , \g2[1][37] , \g2[1][36] ,
         \g2[1][35] , \g2[1][34] , \g2[1][33] , \g2[1][32] , \g2[1][31] ,
         \g2[1][30] , \g2[1][29] , \g2[1][28] , \g2[1][27] , \g2[1][26] ,
         \g2[1][25] , \g2[1][24] , \g2[1][23] , \g2[1][22] , \g2[1][21] ,
         \g2[1][20] , \g2[1][19] , \g2[1][18] , \g2[1][17] , \g2[1][16] ,
         \g2[1][15] , \g2[1][14] , \g2[1][13] , \g2[1][12] , \g2[1][11] ,
         \g2[1][10] , \g2[1][9] , \g2[1][8] , \g2[1][7] , \g2[1][6] ,
         \g2[1][5] , \g2[1][4] , \g2[1][3] , \g2[1][2] , \g2[1][1] ,
         \g2[1][0] , \g2[0][63] , \g2[0][62] , \g2[0][61] , \g2[0][60] ,
         \g2[0][59] , \g2[0][58] , \g2[0][57] , \g2[0][56] , \g2[0][55] ,
         \g2[0][54] , \g2[0][53] , \g2[0][52] , \g2[0][51] , \g2[0][50] ,
         \g2[0][49] , \g2[0][48] , \g2[0][47] , \g2[0][46] , \g2[0][45] ,
         \g2[0][44] , \g2[0][43] , \g2[0][42] , \g2[0][41] , \g2[0][40] ,
         \g2[0][39] , \g2[0][38] , \g2[0][37] , \g2[0][36] , \g2[0][35] ,
         \g2[0][34] , \g2[0][33] , \g2[0][32] , \g2[0][31] , \g2[0][30] ,
         \g2[0][29] , \g2[0][28] , \g2[0][27] , \g2[0][26] , \g2[0][25] ,
         \g2[0][24] , \g2[0][23] , \g2[0][22] , \g2[0][21] , \g2[0][20] ,
         \g2[0][19] , \g2[0][18] , \g2[0][17] , \g2[0][16] , \g2[0][15] ,
         \g2[0][14] , \g2[0][13] , \g2[0][12] , \g2[0][11] , \g2[0][10] ,
         \g2[0][9] , \g2[0][8] , \g2[0][7] , \g2[0][6] , \g2[0][5] ,
         \g2[0][4] , \g2[0][3] , \g2[0][2] , \g2[0][1] , \g2[0][0] ,
         \g3[17][63] , \g3[17][62] , \g3[17][61] , \g3[17][60] , \g3[17][59] ,
         \g3[17][58] , \g3[17][57] , \g3[17][56] , \g3[17][55] , \g3[17][54] ,
         \g3[17][53] , \g3[17][52] , \g3[17][51] , \g3[17][50] , \g3[17][49] ,
         \g3[17][48] , \g3[17][47] , \g3[17][46] , \g3[17][45] , \g3[17][44] ,
         \g3[17][43] , \g3[17][42] , \g3[17][41] , \g3[17][40] , \g3[17][39] ,
         \g3[17][38] , \g3[17][37] , \g3[17][36] , \g3[17][35] , \g3[17][34] ,
         \g3[17][33] , \g3[17][32] , \g3[17][31] , \g3[17][30] , \g3[17][29] ,
         \g3[17][28] , \g3[17][27] , \g3[17][26] , \g3[17][25] , \g3[17][24] ,
         \g3[17][23] , \g3[17][22] , \g3[17][21] , \g3[17][20] , \g3[17][19] ,
         \g3[17][18] , \g3[17][17] , \g3[17][16] , \g3[17][15] , \g3[17][14] ,
         \g3[17][13] , \g3[17][12] , \g3[17][11] , \g3[17][10] , \g3[17][9] ,
         \g3[17][8] , \g3[17][7] , \g3[17][6] , \g3[17][5] , \g3[17][4] ,
         \g3[17][3] , \g3[17][2] , \g3[17][1] , \g3[16][63] , \g3[16][62] ,
         \g3[16][61] , \g3[16][60] , \g3[16][59] , \g3[16][58] , \g3[16][57] ,
         \g3[16][56] , \g3[16][55] , \g3[16][54] , \g3[16][53] , \g3[16][52] ,
         \g3[16][51] , \g3[16][50] , \g3[16][49] , \g3[16][48] , \g3[16][47] ,
         \g3[16][46] , \g3[16][45] , \g3[16][44] , \g3[16][43] , \g3[16][42] ,
         \g3[16][41] , \g3[16][40] , \g3[16][39] , \g3[16][38] , \g3[16][37] ,
         \g3[16][36] , \g3[16][35] , \g3[16][34] , \g3[16][33] , \g3[16][32] ,
         \g3[16][31] , \g3[16][30] , \g3[16][29] , \g3[16][28] , \g3[16][27] ,
         \g3[16][26] , \g3[16][25] , \g3[16][24] , \g3[16][23] , \g3[16][22] ,
         \g3[16][21] , \g3[16][20] , \g3[16][19] , \g3[16][18] , \g3[16][17] ,
         \g3[16][16] , \g3[16][15] , \g3[16][14] , \g3[16][13] , \g3[16][12] ,
         \g3[16][11] , \g3[16][10] , \g3[16][9] , \g3[16][8] , \g3[16][7] ,
         \g3[16][6] , \g3[16][5] , \g3[16][4] , \g3[16][3] , \g3[16][2] ,
         \g3[16][1] , \g3[15][63] , \g3[15][62] , \g3[15][61] , \g3[15][60] ,
         \g3[15][59] , \g3[15][58] , \g3[15][57] , \g3[15][56] , \g3[15][55] ,
         \g3[15][54] , \g3[15][53] , \g3[15][52] , \g3[15][51] , \g3[15][50] ,
         \g3[15][49] , \g3[15][48] , \g3[15][47] , \g3[15][46] , \g3[15][45] ,
         \g3[15][44] , \g3[15][43] , \g3[15][42] , \g3[15][41] , \g3[15][40] ,
         \g3[15][39] , \g3[15][38] , \g3[15][37] , \g3[15][36] , \g3[15][35] ,
         \g3[15][34] , \g3[15][33] , \g3[15][32] , \g3[15][31] , \g3[15][30] ,
         \g3[15][29] , \g3[15][28] , \g3[15][27] , \g3[15][26] , \g3[15][25] ,
         \g3[15][24] , \g3[15][23] , \g3[15][22] , \g3[15][21] , \g3[15][20] ,
         \g3[15][19] , \g3[15][18] , \g3[15][17] , \g3[15][16] , \g3[15][15] ,
         \g3[15][14] , \g3[15][13] , \g3[15][12] , \g3[15][11] , \g3[15][10] ,
         \g3[15][9] , \g3[15][8] , \g3[15][7] , \g3[15][6] , \g3[15][5] ,
         \g3[15][4] , \g3[15][3] , \g3[15][2] , \g3[15][1] , \g3[14][63] ,
         \g3[14][62] , \g3[14][61] , \g3[14][60] , \g3[14][59] , \g3[14][58] ,
         \g3[14][57] , \g3[14][56] , \g3[14][55] , \g3[14][54] , \g3[14][53] ,
         \g3[14][52] , \g3[14][51] , \g3[14][50] , \g3[14][49] , \g3[14][48] ,
         \g3[14][47] , \g3[14][46] , \g3[14][45] , \g3[14][44] , \g3[14][43] ,
         \g3[14][42] , \g3[14][41] , \g3[14][40] , \g3[14][39] , \g3[14][38] ,
         \g3[14][37] , \g3[14][36] , \g3[14][35] , \g3[14][34] , \g3[14][33] ,
         \g3[14][32] , \g3[14][31] , \g3[14][30] , \g3[14][29] , \g3[14][28] ,
         \g3[14][27] , \g3[14][26] , \g3[14][25] , \g3[14][24] , \g3[14][23] ,
         \g3[14][22] , \g3[14][21] , \g3[14][20] , \g3[14][19] , \g3[14][18] ,
         \g3[14][17] , \g3[14][16] , \g3[14][15] , \g3[14][14] , \g3[14][13] ,
         \g3[14][12] , \g3[14][11] , \g3[14][10] , \g3[14][9] , \g3[14][8] ,
         \g3[14][7] , \g3[14][6] , \g3[14][5] , \g3[14][4] , \g3[14][3] ,
         \g3[14][2] , \g3[14][1] , \g3[13][63] , \g3[13][62] , \g3[13][61] ,
         \g3[13][60] , \g3[13][59] , \g3[13][58] , \g3[13][57] , \g3[13][56] ,
         \g3[13][55] , \g3[13][54] , \g3[13][53] , \g3[13][52] , \g3[13][51] ,
         \g3[13][50] , \g3[13][49] , \g3[13][48] , \g3[13][47] , \g3[13][46] ,
         \g3[13][45] , \g3[13][44] , \g3[13][43] , \g3[13][42] , \g3[13][41] ,
         \g3[13][40] , \g3[13][39] , \g3[13][38] , \g3[13][37] , \g3[13][36] ,
         \g3[13][35] , \g3[13][34] , \g3[13][33] , \g3[13][32] , \g3[13][31] ,
         \g3[13][30] , \g3[13][29] , \g3[13][28] , \g3[13][27] , \g3[13][26] ,
         \g3[13][25] , \g3[13][24] , \g3[13][23] , \g3[13][22] , \g3[13][21] ,
         \g3[13][20] , \g3[13][19] , \g3[13][18] , \g3[13][17] , \g3[13][16] ,
         \g3[13][15] , \g3[13][14] , \g3[13][13] , \g3[13][12] , \g3[13][11] ,
         \g3[13][10] , \g3[13][9] , \g3[13][8] , \g3[13][7] , \g3[13][6] ,
         \g3[13][5] , \g3[13][4] , \g3[13][3] , \g3[13][2] , \g3[13][1] ,
         \g3[12][63] , \g3[12][62] , \g3[12][61] , \g3[12][60] , \g3[12][59] ,
         \g3[12][58] , \g3[12][57] , \g3[12][56] , \g3[12][55] , \g3[12][54] ,
         \g3[12][53] , \g3[12][52] , \g3[12][51] , \g3[12][50] , \g3[12][49] ,
         \g3[12][48] , \g3[12][47] , \g3[12][46] , \g3[12][45] , \g3[12][44] ,
         \g3[12][43] , \g3[12][42] , \g3[12][41] , \g3[12][40] , \g3[12][39] ,
         \g3[12][38] , \g3[12][37] , \g3[12][36] , \g3[12][35] , \g3[12][34] ,
         \g3[12][33] , \g3[12][32] , \g3[12][31] , \g3[12][30] , \g3[12][29] ,
         \g3[12][28] , \g3[12][27] , \g3[12][26] , \g3[12][25] , \g3[12][24] ,
         \g3[12][23] , \g3[12][22] , \g3[12][21] , \g3[12][20] , \g3[12][19] ,
         \g3[12][18] , \g3[12][17] , \g3[12][16] , \g3[12][15] , \g3[12][14] ,
         \g3[12][13] , \g3[12][12] , \g3[12][11] , \g3[12][10] , \g3[12][9] ,
         \g3[12][8] , \g3[12][7] , \g3[12][6] , \g3[12][5] , \g3[12][4] ,
         \g3[12][3] , \g3[12][2] , \g3[12][1] , \g3[11][63] , \g3[11][62] ,
         \g3[11][61] , \g3[11][60] , \g3[11][59] , \g3[11][58] , \g3[11][57] ,
         \g3[11][56] , \g3[11][55] , \g3[11][54] , \g3[11][53] , \g3[11][52] ,
         \g3[11][51] , \g3[11][50] , \g3[11][49] , \g3[11][48] , \g3[11][47] ,
         \g3[11][46] , \g3[11][45] , \g3[11][44] , \g3[11][43] , \g3[11][42] ,
         \g3[11][41] , \g3[11][40] , \g3[11][39] , \g3[11][38] , \g3[11][37] ,
         \g3[11][36] , \g3[11][35] , \g3[11][34] , \g3[11][33] , \g3[11][32] ,
         \g3[11][31] , \g3[11][30] , \g3[11][29] , \g3[11][28] , \g3[11][27] ,
         \g3[11][26] , \g3[11][25] , \g3[11][24] , \g3[11][23] , \g3[11][22] ,
         \g3[11][21] , \g3[11][20] , \g3[11][19] , \g3[11][18] , \g3[11][17] ,
         \g3[11][16] , \g3[11][15] , \g3[11][14] , \g3[11][13] , \g3[11][12] ,
         \g3[11][11] , \g3[11][10] , \g3[11][9] , \g3[11][8] , \g3[11][7] ,
         \g3[11][6] , \g3[11][5] , \g3[11][4] , \g3[11][3] , \g3[11][2] ,
         \g3[11][1] , \g3[10][63] , \g3[10][62] , \g3[10][61] , \g3[10][60] ,
         \g3[10][59] , \g3[10][58] , \g3[10][57] , \g3[10][56] , \g3[10][55] ,
         \g3[10][54] , \g3[10][53] , \g3[10][52] , \g3[10][51] , \g3[10][50] ,
         \g3[10][49] , \g3[10][48] , \g3[10][47] , \g3[10][46] , \g3[10][45] ,
         \g3[10][44] , \g3[10][43] , \g3[10][42] , \g3[10][41] , \g3[10][40] ,
         \g3[10][39] , \g3[10][38] , \g3[10][37] , \g3[10][36] , \g3[10][35] ,
         \g3[10][34] , \g3[10][33] , \g3[10][32] , \g3[10][31] , \g3[10][30] ,
         \g3[10][29] , \g3[10][28] , \g3[10][27] , \g3[10][26] , \g3[10][25] ,
         \g3[10][24] , \g3[10][23] , \g3[10][22] , \g3[10][21] , \g3[10][20] ,
         \g3[10][19] , \g3[10][18] , \g3[10][17] , \g3[10][16] , \g3[10][15] ,
         \g3[10][14] , \g3[10][13] , \g3[10][12] , \g3[10][11] , \g3[10][10] ,
         \g3[10][9] , \g3[10][8] , \g3[10][7] , \g3[10][6] , \g3[10][5] ,
         \g3[10][4] , \g3[10][3] , \g3[10][2] , \g3[10][1] , \g3[9][63] ,
         \g3[9][62] , \g3[9][61] , \g3[9][60] , \g3[9][59] , \g3[9][58] ,
         \g3[9][57] , \g3[9][56] , \g3[9][55] , \g3[9][54] , \g3[9][53] ,
         \g3[9][52] , \g3[9][51] , \g3[9][50] , \g3[9][49] , \g3[9][48] ,
         \g3[9][47] , \g3[9][46] , \g3[9][45] , \g3[9][44] , \g3[9][43] ,
         \g3[9][42] , \g3[9][41] , \g3[9][40] , \g3[9][39] , \g3[9][38] ,
         \g3[9][37] , \g3[9][36] , \g3[9][35] , \g3[9][34] , \g3[9][33] ,
         \g3[9][32] , \g3[9][31] , \g3[9][30] , \g3[9][29] , \g3[9][28] ,
         \g3[9][27] , \g3[9][26] , \g3[9][25] , \g3[9][24] , \g3[9][23] ,
         \g3[9][22] , \g3[9][21] , \g3[9][20] , \g3[9][19] , \g3[9][18] ,
         \g3[9][17] , \g3[9][16] , \g3[9][15] , \g3[9][14] , \g3[9][13] ,
         \g3[9][12] , \g3[9][11] , \g3[9][10] , \g3[9][9] , \g3[9][8] ,
         \g3[9][7] , \g3[9][6] , \g3[9][5] , \g3[9][4] , \g3[9][3] ,
         \g3[9][2] , \g3[9][1] , \g3[8][63] , \g3[8][62] , \g3[8][61] ,
         \g3[8][60] , \g3[8][59] , \g3[8][58] , \g3[8][57] , \g3[8][56] ,
         \g3[8][55] , \g3[8][54] , \g3[8][53] , \g3[8][52] , \g3[8][51] ,
         \g3[8][50] , \g3[8][49] , \g3[8][48] , \g3[8][47] , \g3[8][46] ,
         \g3[8][45] , \g3[8][44] , \g3[8][43] , \g3[8][42] , \g3[8][41] ,
         \g3[8][40] , \g3[8][39] , \g3[8][38] , \g3[8][37] , \g3[8][36] ,
         \g3[8][35] , \g3[8][34] , \g3[8][33] , \g3[8][32] , \g3[8][31] ,
         \g3[8][30] , \g3[8][29] , \g3[8][28] , \g3[8][27] , \g3[8][26] ,
         \g3[8][25] , \g3[8][24] , \g3[8][23] , \g3[8][22] , \g3[8][21] ,
         \g3[8][20] , \g3[8][19] , \g3[8][18] , \g3[8][17] , \g3[8][16] ,
         \g3[8][15] , \g3[8][14] , \g3[8][13] , \g3[8][12] , \g3[8][11] ,
         \g3[8][10] , \g3[8][9] , \g3[8][8] , \g3[8][7] , \g3[8][6] ,
         \g3[8][5] , \g3[8][4] , \g3[8][3] , \g3[8][2] , \g3[8][1] ,
         \g3[8][0] , \g3[7][63] , \g3[7][62] , \g3[7][61] , \g3[7][60] ,
         \g3[7][59] , \g3[7][58] , \g3[7][57] , \g3[7][56] , \g3[7][55] ,
         \g3[7][54] , \g3[7][53] , \g3[7][52] , \g3[7][51] , \g3[7][50] ,
         \g3[7][49] , \g3[7][48] , \g3[7][47] , \g3[7][46] , \g3[7][45] ,
         \g3[7][44] , \g3[7][43] , \g3[7][42] , \g3[7][41] , \g3[7][40] ,
         \g3[7][39] , \g3[7][38] , \g3[7][37] , \g3[7][36] , \g3[7][35] ,
         \g3[7][34] , \g3[7][33] , \g3[7][32] , \g3[7][31] , \g3[7][30] ,
         \g3[7][29] , \g3[7][28] , \g3[7][27] , \g3[7][26] , \g3[7][25] ,
         \g3[7][24] , \g3[7][23] , \g3[7][22] , \g3[7][21] , \g3[7][20] ,
         \g3[7][19] , \g3[7][18] , \g3[7][17] , \g3[7][16] , \g3[7][15] ,
         \g3[7][14] , \g3[7][13] , \g3[7][12] , \g3[7][11] , \g3[7][10] ,
         \g3[7][9] , \g3[7][8] , \g3[7][7] , \g3[7][6] , \g3[7][5] ,
         \g3[7][4] , \g3[7][3] , \g3[7][2] , \g3[7][1] , \g3[7][0] ,
         \g3[6][63] , \g3[6][62] , \g3[6][61] , \g3[6][60] , \g3[6][59] ,
         \g3[6][58] , \g3[6][57] , \g3[6][56] , \g3[6][55] , \g3[6][54] ,
         \g3[6][53] , \g3[6][52] , \g3[6][51] , \g3[6][50] , \g3[6][49] ,
         \g3[6][48] , \g3[6][47] , \g3[6][46] , \g3[6][45] , \g3[6][44] ,
         \g3[6][43] , \g3[6][42] , \g3[6][41] , \g3[6][40] , \g3[6][39] ,
         \g3[6][38] , \g3[6][37] , \g3[6][36] , \g3[6][35] , \g3[6][34] ,
         \g3[6][33] , \g3[6][32] , \g3[6][31] , \g3[6][30] , \g3[6][29] ,
         \g3[6][28] , \g3[6][27] , \g3[6][26] , \g3[6][25] , \g3[6][24] ,
         \g3[6][23] , \g3[6][22] , \g3[6][21] , \g3[6][20] , \g3[6][19] ,
         \g3[6][18] , \g3[6][17] , \g3[6][16] , \g3[6][15] , \g3[6][14] ,
         \g3[6][13] , \g3[6][12] , \g3[6][11] , \g3[6][10] , \g3[6][9] ,
         \g3[6][8] , \g3[6][7] , \g3[6][6] , \g3[6][5] , \g3[6][4] ,
         \g3[6][3] , \g3[6][2] , \g3[6][1] , \g3[6][0] , \g3[5][63] ,
         \g3[5][62] , \g3[5][61] , \g3[5][60] , \g3[5][59] , \g3[5][58] ,
         \g3[5][57] , \g3[5][56] , \g3[5][55] , \g3[5][54] , \g3[5][53] ,
         \g3[5][52] , \g3[5][51] , \g3[5][50] , \g3[5][49] , \g3[5][48] ,
         \g3[5][47] , \g3[5][46] , \g3[5][45] , \g3[5][44] , \g3[5][43] ,
         \g3[5][42] , \g3[5][41] , \g3[5][40] , \g3[5][39] , \g3[5][38] ,
         \g3[5][37] , \g3[5][36] , \g3[5][35] , \g3[5][34] , \g3[5][33] ,
         \g3[5][32] , \g3[5][31] , \g3[5][30] , \g3[5][29] , \g3[5][28] ,
         \g3[5][27] , \g3[5][26] , \g3[5][25] , \g3[5][24] , \g3[5][23] ,
         \g3[5][22] , \g3[5][21] , \g3[5][20] , \g3[5][19] , \g3[5][18] ,
         \g3[5][17] , \g3[5][16] , \g3[5][15] , \g3[5][14] , \g3[5][13] ,
         \g3[5][12] , \g3[5][11] , \g3[5][10] , \g3[5][9] , \g3[5][8] ,
         \g3[5][7] , \g3[5][6] , \g3[5][5] , \g3[5][4] , \g3[5][3] ,
         \g3[5][2] , \g3[5][1] , \g3[5][0] , \g3[4][63] , \g3[4][62] ,
         \g3[4][61] , \g3[4][60] , \g3[4][59] , \g3[4][58] , \g3[4][57] ,
         \g3[4][56] , \g3[4][55] , \g3[4][54] , \g3[4][53] , \g3[4][52] ,
         \g3[4][51] , \g3[4][50] , \g3[4][49] , \g3[4][48] , \g3[4][47] ,
         \g3[4][46] , \g3[4][45] , \g3[4][44] , \g3[4][43] , \g3[4][42] ,
         \g3[4][41] , \g3[4][40] , \g3[4][39] , \g3[4][38] , \g3[4][37] ,
         \g3[4][36] , \g3[4][35] , \g3[4][34] , \g3[4][33] , \g3[4][32] ,
         \g3[4][31] , \g3[4][30] , \g3[4][29] , \g3[4][28] , \g3[4][27] ,
         \g3[4][26] , \g3[4][25] , \g3[4][24] , \g3[4][23] , \g3[4][22] ,
         \g3[4][21] , \g3[4][20] , \g3[4][19] , \g3[4][18] , \g3[4][17] ,
         \g3[4][16] , \g3[4][15] , \g3[4][14] , \g3[4][13] , \g3[4][12] ,
         \g3[4][11] , \g3[4][10] , \g3[4][9] , \g3[4][8] , \g3[4][7] ,
         \g3[4][6] , \g3[4][5] , \g3[4][4] , \g3[4][3] , \g3[4][2] ,
         \g3[4][1] , \g3[4][0] , \g3[3][63] , \g3[3][62] , \g3[3][61] ,
         \g3[3][60] , \g3[3][59] , \g3[3][58] , \g3[3][57] , \g3[3][56] ,
         \g3[3][55] , \g3[3][54] , \g3[3][53] , \g3[3][52] , \g3[3][51] ,
         \g3[3][50] , \g3[3][49] , \g3[3][48] , \g3[3][47] , \g3[3][46] ,
         \g3[3][45] , \g3[3][44] , \g3[3][43] , \g3[3][42] , \g3[3][41] ,
         \g3[3][40] , \g3[3][39] , \g3[3][38] , \g3[3][37] , \g3[3][36] ,
         \g3[3][35] , \g3[3][34] , \g3[3][33] , \g3[3][32] , \g3[3][31] ,
         \g3[3][30] , \g3[3][29] , \g3[3][28] , \g3[3][27] , \g3[3][26] ,
         \g3[3][25] , \g3[3][24] , \g3[3][23] , \g3[3][22] , \g3[3][21] ,
         \g3[3][20] , \g3[3][19] , \g3[3][18] , \g3[3][17] , \g3[3][16] ,
         \g3[3][15] , \g3[3][14] , \g3[3][13] , \g3[3][12] , \g3[3][11] ,
         \g3[3][10] , \g3[3][9] , \g3[3][8] , \g3[3][7] , \g3[3][6] ,
         \g3[3][5] , \g3[3][4] , \g3[3][3] , \g3[3][2] , \g3[3][1] ,
         \g3[3][0] , \g3[2][63] , \g3[2][62] , \g3[2][61] , \g3[2][60] ,
         \g3[2][59] , \g3[2][58] , \g3[2][57] , \g3[2][56] , \g3[2][55] ,
         \g3[2][54] , \g3[2][53] , \g3[2][52] , \g3[2][51] , \g3[2][50] ,
         \g3[2][49] , \g3[2][48] , \g3[2][47] , \g3[2][46] , \g3[2][45] ,
         \g3[2][44] , \g3[2][43] , \g3[2][42] , \g3[2][41] , \g3[2][40] ,
         \g3[2][39] , \g3[2][38] , \g3[2][37] , \g3[2][36] , \g3[2][35] ,
         \g3[2][34] , \g3[2][33] , \g3[2][32] , \g3[2][31] , \g3[2][30] ,
         \g3[2][29] , \g3[2][28] , \g3[2][27] , \g3[2][26] , \g3[2][25] ,
         \g3[2][24] , \g3[2][23] , \g3[2][22] , \g3[2][21] , \g3[2][20] ,
         \g3[2][19] , \g3[2][18] , \g3[2][17] , \g3[2][16] , \g3[2][15] ,
         \g3[2][14] , \g3[2][13] , \g3[2][12] , \g3[2][11] , \g3[2][10] ,
         \g3[2][9] , \g3[2][8] , \g3[2][7] , \g3[2][6] , \g3[2][5] ,
         \g3[2][4] , \g3[2][3] , \g3[2][2] , \g3[2][1] , \g3[2][0] ,
         \g3[1][63] , \g3[1][62] , \g3[1][61] , \g3[1][60] , \g3[1][59] ,
         \g3[1][58] , \g3[1][57] , \g3[1][56] , \g3[1][55] , \g3[1][54] ,
         \g3[1][53] , \g3[1][52] , \g3[1][51] , \g3[1][50] , \g3[1][49] ,
         \g3[1][48] , \g3[1][47] , \g3[1][46] , \g3[1][45] , \g3[1][44] ,
         \g3[1][43] , \g3[1][42] , \g3[1][41] , \g3[1][40] , \g3[1][39] ,
         \g3[1][38] , \g3[1][37] , \g3[1][36] , \g3[1][35] , \g3[1][34] ,
         \g3[1][33] , \g3[1][32] , \g3[1][31] , \g3[1][30] , \g3[1][29] ,
         \g3[1][28] , \g3[1][27] , \g3[1][26] , \g3[1][25] , \g3[1][24] ,
         \g3[1][23] , \g3[1][22] , \g3[1][21] , \g3[1][20] , \g3[1][19] ,
         \g3[1][18] , \g3[1][17] , \g3[1][16] , \g3[1][15] , \g3[1][14] ,
         \g3[1][13] , \g3[1][12] , \g3[1][11] , \g3[1][10] , \g3[1][9] ,
         \g3[1][8] , \g3[1][7] , \g3[1][6] , \g3[1][5] , \g3[1][4] ,
         \g3[1][3] , \g3[1][2] , \g3[1][1] , \g3[1][0] , \g3[0][63] ,
         \g3[0][62] , \g3[0][61] , \g3[0][60] , \g3[0][59] , \g3[0][58] ,
         \g3[0][57] , \g3[0][56] , \g3[0][55] , \g3[0][54] , \g3[0][53] ,
         \g3[0][52] , \g3[0][51] , \g3[0][50] , \g3[0][49] , \g3[0][48] ,
         \g3[0][47] , \g3[0][46] , \g3[0][45] , \g3[0][44] , \g3[0][43] ,
         \g3[0][42] , \g3[0][41] , \g3[0][40] , \g3[0][39] , \g3[0][38] ,
         \g3[0][37] , \g3[0][36] , \g3[0][35] , \g3[0][34] , \g3[0][33] ,
         \g3[0][32] , \g3[0][31] , \g3[0][30] , \g3[0][29] , \g3[0][28] ,
         \g3[0][27] , \g3[0][26] , \g3[0][25] , \g3[0][24] , \g3[0][23] ,
         \g3[0][22] , \g3[0][21] , \g3[0][20] , \g3[0][19] , \g3[0][18] ,
         \g3[0][17] , \g3[0][16] , \g3[0][15] , \g3[0][14] , \g3[0][13] ,
         \g3[0][12] , \g3[0][11] , \g3[0][10] , \g3[0][9] , \g3[0][8] ,
         \g3[0][7] , \g3[0][6] , \g3[0][5] , \g3[0][4] , \g3[0][3] ,
         \g3[0][2] , \g3[0][1] , \g3[0][0] , \g4[11][63] , \g4[11][62] ,
         \g4[11][61] , \g4[11][60] , \g4[11][59] , \g4[11][58] , \g4[11][57] ,
         \g4[11][56] , \g4[11][55] , \g4[11][54] , \g4[11][53] , \g4[11][52] ,
         \g4[11][51] , \g4[11][50] , \g4[11][49] , \g4[11][48] , \g4[11][47] ,
         \g4[11][46] , \g4[11][45] , \g4[11][44] , \g4[11][43] , \g4[11][42] ,
         \g4[11][41] , \g4[11][40] , \g4[11][39] , \g4[11][38] , \g4[11][37] ,
         \g4[11][36] , \g4[11][35] , \g4[11][34] , \g4[11][33] , \g4[11][32] ,
         \g4[11][31] , \g4[11][30] , \g4[11][29] , \g4[11][28] , \g4[11][27] ,
         \g4[11][26] , \g4[11][25] , \g4[11][24] , \g4[11][23] , \g4[11][22] ,
         \g4[11][21] , \g4[11][20] , \g4[11][19] , \g4[11][18] , \g4[11][17] ,
         \g4[11][16] , \g4[11][15] , \g4[11][14] , \g4[11][13] , \g4[11][12] ,
         \g4[11][11] , \g4[11][10] , \g4[11][9] , \g4[11][8] , \g4[11][7] ,
         \g4[11][6] , \g4[11][5] , \g4[11][4] , \g4[11][3] , \g4[11][2] ,
         \g4[11][1] , \g4[10][63] , \g4[10][62] , \g4[10][61] , \g4[10][60] ,
         \g4[10][59] , \g4[10][58] , \g4[10][57] , \g4[10][56] , \g4[10][55] ,
         \g4[10][54] , \g4[10][53] , \g4[10][52] , \g4[10][51] , \g4[10][50] ,
         \g4[10][49] , \g4[10][48] , \g4[10][47] , \g4[10][46] , \g4[10][45] ,
         \g4[10][44] , \g4[10][43] , \g4[10][42] , \g4[10][41] , \g4[10][40] ,
         \g4[10][39] , \g4[10][38] , \g4[10][37] , \g4[10][36] , \g4[10][35] ,
         \g4[10][34] , \g4[10][33] , \g4[10][32] , \g4[10][31] , \g4[10][30] ,
         \g4[10][29] , \g4[10][28] , \g4[10][27] , \g4[10][26] , \g4[10][25] ,
         \g4[10][24] , \g4[10][23] , \g4[10][22] , \g4[10][21] , \g4[10][20] ,
         \g4[10][19] , \g4[10][18] , \g4[10][17] , \g4[10][16] , \g4[10][15] ,
         \g4[10][14] , \g4[10][13] , \g4[10][12] , \g4[10][11] , \g4[10][10] ,
         \g4[10][9] , \g4[10][8] , \g4[10][7] , \g4[10][6] , \g4[10][5] ,
         \g4[10][4] , \g4[10][3] , \g4[10][2] , \g4[10][1] , \g4[9][63] ,
         \g4[9][62] , \g4[9][61] , \g4[9][60] , \g4[9][59] , \g4[9][58] ,
         \g4[9][57] , \g4[9][56] , \g4[9][55] , \g4[9][54] , \g4[9][53] ,
         \g4[9][52] , \g4[9][51] , \g4[9][50] , \g4[9][49] , \g4[9][48] ,
         \g4[9][47] , \g4[9][46] , \g4[9][45] , \g4[9][44] , \g4[9][43] ,
         \g4[9][42] , \g4[9][41] , \g4[9][40] , \g4[9][39] , \g4[9][38] ,
         \g4[9][37] , \g4[9][36] , \g4[9][35] , \g4[9][34] , \g4[9][33] ,
         \g4[9][32] , \g4[9][31] , \g4[9][30] , \g4[9][29] , \g4[9][28] ,
         \g4[9][27] , \g4[9][26] , \g4[9][25] , \g4[9][24] , \g4[9][23] ,
         \g4[9][22] , \g4[9][21] , \g4[9][20] , \g4[9][19] , \g4[9][18] ,
         \g4[9][17] , \g4[9][16] , \g4[9][15] , \g4[9][14] , \g4[9][13] ,
         \g4[9][12] , \g4[9][11] , \g4[9][10] , \g4[9][9] , \g4[9][8] ,
         \g4[9][7] , \g4[9][6] , \g4[9][5] , \g4[9][4] , \g4[9][3] ,
         \g4[9][2] , \g4[9][1] , \g4[8][63] , \g4[8][62] , \g4[8][61] ,
         \g4[8][60] , \g4[8][59] , \g4[8][58] , \g4[8][57] , \g4[8][56] ,
         \g4[8][55] , \g4[8][54] , \g4[8][53] , \g4[8][52] , \g4[8][51] ,
         \g4[8][50] , \g4[8][49] , \g4[8][48] , \g4[8][47] , \g4[8][46] ,
         \g4[8][45] , \g4[8][44] , \g4[8][43] , \g4[8][42] , \g4[8][41] ,
         \g4[8][40] , \g4[8][39] , \g4[8][38] , \g4[8][37] , \g4[8][36] ,
         \g4[8][35] , \g4[8][34] , \g4[8][33] , \g4[8][32] , \g4[8][31] ,
         \g4[8][30] , \g4[8][29] , \g4[8][28] , \g4[8][27] , \g4[8][26] ,
         \g4[8][25] , \g4[8][24] , \g4[8][23] , \g4[8][22] , \g4[8][21] ,
         \g4[8][20] , \g4[8][19] , \g4[8][18] , \g4[8][17] , \g4[8][16] ,
         \g4[8][15] , \g4[8][14] , \g4[8][13] , \g4[8][12] , \g4[8][11] ,
         \g4[8][10] , \g4[8][9] , \g4[8][8] , \g4[8][7] , \g4[8][6] ,
         \g4[8][5] , \g4[8][4] , \g4[8][3] , \g4[8][2] , \g4[8][1] ,
         \g4[7][63] , \g4[7][62] , \g4[7][61] , \g4[7][60] , \g4[7][59] ,
         \g4[7][58] , \g4[7][57] , \g4[7][56] , \g4[7][55] , \g4[7][54] ,
         \g4[7][53] , \g4[7][52] , \g4[7][51] , \g4[7][50] , \g4[7][49] ,
         \g4[7][48] , \g4[7][47] , \g4[7][46] , \g4[7][45] , \g4[7][44] ,
         \g4[7][43] , \g4[7][42] , \g4[7][41] , \g4[7][40] , \g4[7][39] ,
         \g4[7][38] , \g4[7][37] , \g4[7][36] , \g4[7][35] , \g4[7][34] ,
         \g4[7][33] , \g4[7][32] , \g4[7][31] , \g4[7][30] , \g4[7][29] ,
         \g4[7][28] , \g4[7][27] , \g4[7][26] , \g4[7][25] , \g4[7][24] ,
         \g4[7][23] , \g4[7][22] , \g4[7][21] , \g4[7][20] , \g4[7][19] ,
         \g4[7][18] , \g4[7][17] , \g4[7][16] , \g4[7][15] , \g4[7][14] ,
         \g4[7][13] , \g4[7][12] , \g4[7][11] , \g4[7][10] , \g4[7][9] ,
         \g4[7][8] , \g4[7][7] , \g4[7][6] , \g4[7][5] , \g4[7][4] ,
         \g4[7][3] , \g4[7][2] , \g4[7][1] , \g4[6][63] , \g4[6][62] ,
         \g4[6][61] , \g4[6][60] , \g4[6][59] , \g4[6][58] , \g4[6][57] ,
         \g4[6][56] , \g4[6][55] , \g4[6][54] , \g4[6][53] , \g4[6][52] ,
         \g4[6][51] , \g4[6][50] , \g4[6][49] , \g4[6][48] , \g4[6][47] ,
         \g4[6][46] , \g4[6][45] , \g4[6][44] , \g4[6][43] , \g4[6][42] ,
         \g4[6][41] , \g4[6][40] , \g4[6][39] , \g4[6][38] , \g4[6][37] ,
         \g4[6][36] , \g4[6][35] , \g4[6][34] , \g4[6][33] , \g4[6][32] ,
         \g4[6][31] , \g4[6][30] , \g4[6][29] , \g4[6][28] , \g4[6][27] ,
         \g4[6][26] , \g4[6][25] , \g4[6][24] , \g4[6][23] , \g4[6][22] ,
         \g4[6][21] , \g4[6][20] , \g4[6][19] , \g4[6][18] , \g4[6][17] ,
         \g4[6][16] , \g4[6][15] , \g4[6][14] , \g4[6][13] , \g4[6][12] ,
         \g4[6][11] , \g4[6][10] , \g4[6][9] , \g4[6][8] , \g4[6][7] ,
         \g4[6][6] , \g4[6][5] , \g4[6][4] , \g4[6][3] , \g4[6][2] ,
         \g4[6][1] , \g4[5][63] , \g4[5][62] , \g4[5][61] , \g4[5][60] ,
         \g4[5][59] , \g4[5][58] , \g4[5][57] , \g4[5][56] , \g4[5][55] ,
         \g4[5][54] , \g4[5][53] , \g4[5][52] , \g4[5][51] , \g4[5][50] ,
         \g4[5][49] , \g4[5][48] , \g4[5][47] , \g4[5][46] , \g4[5][45] ,
         \g4[5][44] , \g4[5][43] , \g4[5][42] , \g4[5][41] , \g4[5][40] ,
         \g4[5][39] , \g4[5][38] , \g4[5][37] , \g4[5][36] , \g4[5][35] ,
         \g4[5][34] , \g4[5][33] , \g4[5][32] , \g4[5][31] , \g4[5][30] ,
         \g4[5][29] , \g4[5][28] , \g4[5][27] , \g4[5][26] , \g4[5][25] ,
         \g4[5][24] , \g4[5][23] , \g4[5][22] , \g4[5][21] , \g4[5][20] ,
         \g4[5][19] , \g4[5][18] , \g4[5][17] , \g4[5][16] , \g4[5][15] ,
         \g4[5][14] , \g4[5][13] , \g4[5][12] , \g4[5][11] , \g4[5][10] ,
         \g4[5][9] , \g4[5][8] , \g4[5][7] , \g4[5][6] , \g4[5][5] ,
         \g4[5][4] , \g4[5][3] , \g4[5][2] , \g4[5][1] , \g4[5][0] ,
         \g4[4][63] , \g4[4][62] , \g4[4][61] , \g4[4][60] , \g4[4][59] ,
         \g4[4][58] , \g4[4][57] , \g4[4][56] , \g4[4][55] , \g4[4][54] ,
         \g4[4][53] , \g4[4][52] , \g4[4][51] , \g4[4][50] , \g4[4][49] ,
         \g4[4][48] , \g4[4][47] , \g4[4][46] , \g4[4][45] , \g4[4][44] ,
         \g4[4][43] , \g4[4][42] , \g4[4][41] , \g4[4][40] , \g4[4][39] ,
         \g4[4][38] , \g4[4][37] , \g4[4][36] , \g4[4][35] , \g4[4][34] ,
         \g4[4][33] , \g4[4][32] , \g4[4][31] , \g4[4][30] , \g4[4][29] ,
         \g4[4][28] , \g4[4][27] , \g4[4][26] , \g4[4][25] , \g4[4][24] ,
         \g4[4][23] , \g4[4][22] , \g4[4][21] , \g4[4][20] , \g4[4][19] ,
         \g4[4][18] , \g4[4][17] , \g4[4][16] , \g4[4][15] , \g4[4][14] ,
         \g4[4][13] , \g4[4][12] , \g4[4][11] , \g4[4][10] , \g4[4][9] ,
         \g4[4][8] , \g4[4][7] , \g4[4][6] , \g4[4][5] , \g4[4][4] ,
         \g4[4][3] , \g4[4][2] , \g4[4][1] , \g4[4][0] , \g4[3][63] ,
         \g4[3][62] , \g4[3][61] , \g4[3][60] , \g4[3][59] , \g4[3][58] ,
         \g4[3][57] , \g4[3][56] , \g4[3][55] , \g4[3][54] , \g4[3][53] ,
         \g4[3][52] , \g4[3][51] , \g4[3][50] , \g4[3][49] , \g4[3][48] ,
         \g4[3][47] , \g4[3][46] , \g4[3][45] , \g4[3][44] , \g4[3][43] ,
         \g4[3][42] , \g4[3][41] , \g4[3][40] , \g4[3][39] , \g4[3][38] ,
         \g4[3][37] , \g4[3][36] , \g4[3][35] , \g4[3][34] , \g4[3][33] ,
         \g4[3][32] , \g4[3][31] , \g4[3][30] , \g4[3][29] , \g4[3][28] ,
         \g4[3][27] , \g4[3][26] , \g4[3][25] , \g4[3][24] , \g4[3][23] ,
         \g4[3][22] , \g4[3][21] , \g4[3][20] , \g4[3][19] , \g4[3][18] ,
         \g4[3][17] , \g4[3][16] , \g4[3][15] , \g4[3][14] , \g4[3][13] ,
         \g4[3][12] , \g4[3][11] , \g4[3][10] , \g4[3][9] , \g4[3][8] ,
         \g4[3][7] , \g4[3][6] , \g4[3][5] , \g4[3][4] , \g4[3][3] ,
         \g4[3][2] , \g4[3][1] , \g4[3][0] , \g4[2][63] , \g4[2][62] ,
         \g4[2][61] , \g4[2][60] , \g4[2][59] , \g4[2][58] , \g4[2][57] ,
         \g4[2][56] , \g4[2][55] , \g4[2][54] , \g4[2][53] , \g4[2][52] ,
         \g4[2][51] , \g4[2][50] , \g4[2][49] , \g4[2][48] , \g4[2][47] ,
         \g4[2][46] , \g4[2][45] , \g4[2][44] , \g4[2][43] , \g4[2][42] ,
         \g4[2][41] , \g4[2][40] , \g4[2][39] , \g4[2][38] , \g4[2][37] ,
         \g4[2][36] , \g4[2][35] , \g4[2][34] , \g4[2][33] , \g4[2][32] ,
         \g4[2][31] , \g4[2][30] , \g4[2][29] , \g4[2][28] , \g4[2][27] ,
         \g4[2][26] , \g4[2][25] , \g4[2][24] , \g4[2][23] , \g4[2][22] ,
         \g4[2][21] , \g4[2][20] , \g4[2][19] , \g4[2][18] , \g4[2][17] ,
         \g4[2][16] , \g4[2][15] , \g4[2][14] , \g4[2][13] , \g4[2][12] ,
         \g4[2][11] , \g4[2][10] , \g4[2][9] , \g4[2][8] , \g4[2][7] ,
         \g4[2][6] , \g4[2][5] , \g4[2][4] , \g4[2][3] , \g4[2][2] ,
         \g4[2][1] , \g4[2][0] , \g4[1][63] , \g4[1][62] , \g4[1][61] ,
         \g4[1][60] , \g4[1][59] , \g4[1][58] , \g4[1][57] , \g4[1][56] ,
         \g4[1][55] , \g4[1][54] , \g4[1][53] , \g4[1][52] , \g4[1][51] ,
         \g4[1][50] , \g4[1][49] , \g4[1][48] , \g4[1][47] , \g4[1][46] ,
         \g4[1][45] , \g4[1][44] , \g4[1][43] , \g4[1][42] , \g4[1][41] ,
         \g4[1][40] , \g4[1][39] , \g4[1][38] , \g4[1][37] , \g4[1][36] ,
         \g4[1][35] , \g4[1][34] , \g4[1][33] , \g4[1][32] , \g4[1][31] ,
         \g4[1][30] , \g4[1][29] , \g4[1][28] , \g4[1][27] , \g4[1][26] ,
         \g4[1][25] , \g4[1][24] , \g4[1][23] , \g4[1][22] , \g4[1][21] ,
         \g4[1][20] , \g4[1][19] , \g4[1][18] , \g4[1][17] , \g4[1][16] ,
         \g4[1][15] , \g4[1][14] , \g4[1][13] , \g4[1][12] , \g4[1][11] ,
         \g4[1][10] , \g4[1][9] , \g4[1][8] , \g4[1][7] , \g4[1][6] ,
         \g4[1][5] , \g4[1][4] , \g4[1][3] , \g4[1][2] , \g4[1][1] ,
         \g4[1][0] , \g4[0][63] , \g4[0][62] , \g4[0][61] , \g4[0][60] ,
         \g4[0][59] , \g4[0][58] , \g4[0][57] , \g4[0][56] , \g4[0][55] ,
         \g4[0][54] , \g4[0][53] , \g4[0][52] , \g4[0][51] , \g4[0][50] ,
         \g4[0][49] , \g4[0][48] , \g4[0][47] , \g4[0][46] , \g4[0][45] ,
         \g4[0][44] , \g4[0][43] , \g4[0][42] , \g4[0][41] , \g4[0][40] ,
         \g4[0][39] , \g4[0][38] , \g4[0][37] , \g4[0][36] , \g4[0][35] ,
         \g4[0][34] , \g4[0][33] , \g4[0][32] , \g4[0][31] , \g4[0][30] ,
         \g4[0][29] , \g4[0][28] , \g4[0][27] , \g4[0][26] , \g4[0][25] ,
         \g4[0][24] , \g4[0][23] , \g4[0][22] , \g4[0][21] , \g4[0][20] ,
         \g4[0][19] , \g4[0][18] , \g4[0][17] , \g4[0][16] , \g4[0][15] ,
         \g4[0][14] , \g4[0][13] , \g4[0][12] , \g4[0][11] , \g4[0][10] ,
         \g4[0][9] , \g4[0][8] , \g4[0][7] , \g4[0][6] , \g4[0][5] ,
         \g4[0][4] , \g4[0][3] , \g4[0][2] , \g4[0][1] , \g4[0][0] ,
         \g5[7][63] , \g5[7][62] , \g5[7][61] , \g5[7][60] , \g5[7][59] ,
         \g5[7][58] , \g5[7][57] , \g5[7][56] , \g5[7][55] , \g5[7][54] ,
         \g5[7][53] , \g5[7][52] , \g5[7][51] , \g5[7][50] , \g5[7][49] ,
         \g5[7][48] , \g5[7][47] , \g5[7][46] , \g5[7][45] , \g5[7][44] ,
         \g5[7][43] , \g5[7][42] , \g5[7][41] , \g5[7][40] , \g5[7][39] ,
         \g5[7][38] , \g5[7][37] , \g5[7][36] , \g5[7][35] , \g5[7][34] ,
         \g5[7][33] , \g5[7][32] , \g5[7][31] , \g5[7][30] , \g5[7][29] ,
         \g5[7][28] , \g5[7][27] , \g5[7][26] , \g5[7][25] , \g5[7][24] ,
         \g5[7][23] , \g5[7][22] , \g5[7][21] , \g5[7][20] , \g5[7][19] ,
         \g5[7][18] , \g5[7][17] , \g5[7][16] , \g5[7][15] , \g5[7][14] ,
         \g5[7][13] , \g5[7][12] , \g5[7][11] , \g5[7][10] , \g5[7][9] ,
         \g5[7][8] , \g5[7][7] , \g5[7][6] , \g5[7][5] , \g5[7][4] ,
         \g5[7][3] , \g5[7][2] , \g5[7][1] , \g5[6][63] , \g5[6][62] ,
         \g5[6][61] , \g5[6][60] , \g5[6][59] , \g5[6][58] , \g5[6][57] ,
         \g5[6][56] , \g5[6][55] , \g5[6][54] , \g5[6][53] , \g5[6][52] ,
         \g5[6][51] , \g5[6][50] , \g5[6][49] , \g5[6][48] , \g5[6][47] ,
         \g5[6][46] , \g5[6][45] , \g5[6][44] , \g5[6][43] , \g5[6][42] ,
         \g5[6][41] , \g5[6][40] , \g5[6][39] , \g5[6][38] , \g5[6][37] ,
         \g5[6][36] , \g5[6][35] , \g5[6][34] , \g5[6][33] , \g5[6][32] ,
         \g5[6][31] , \g5[6][30] , \g5[6][29] , \g5[6][28] , \g5[6][27] ,
         \g5[6][26] , \g5[6][25] , \g5[6][24] , \g5[6][23] , \g5[6][22] ,
         \g5[6][21] , \g5[6][20] , \g5[6][19] , \g5[6][18] , \g5[6][17] ,
         \g5[6][16] , \g5[6][15] , \g5[6][14] , \g5[6][13] , \g5[6][12] ,
         \g5[6][11] , \g5[6][10] , \g5[6][9] , \g5[6][8] , \g5[6][7] ,
         \g5[6][6] , \g5[6][5] , \g5[6][4] , \g5[6][3] , \g5[6][2] ,
         \g5[6][1] , \g5[5][63] , \g5[5][62] , \g5[5][61] , \g5[5][60] ,
         \g5[5][59] , \g5[5][58] , \g5[5][57] , \g5[5][56] , \g5[5][55] ,
         \g5[5][54] , \g5[5][53] , \g5[5][52] , \g5[5][51] , \g5[5][50] ,
         \g5[5][49] , \g5[5][48] , \g5[5][47] , \g5[5][46] , \g5[5][45] ,
         \g5[5][44] , \g5[5][43] , \g5[5][42] , \g5[5][41] , \g5[5][40] ,
         \g5[5][39] , \g5[5][38] , \g5[5][37] , \g5[5][36] , \g5[5][35] ,
         \g5[5][34] , \g5[5][33] , \g5[5][32] , \g5[5][31] , \g5[5][30] ,
         \g5[5][29] , \g5[5][28] , \g5[5][27] , \g5[5][26] , \g5[5][25] ,
         \g5[5][24] , \g5[5][23] , \g5[5][22] , \g5[5][21] , \g5[5][20] ,
         \g5[5][19] , \g5[5][18] , \g5[5][17] , \g5[5][16] , \g5[5][15] ,
         \g5[5][14] , \g5[5][13] , \g5[5][12] , \g5[5][11] , \g5[5][10] ,
         \g5[5][9] , \g5[5][8] , \g5[5][7] , \g5[5][6] , \g5[5][5] ,
         \g5[5][4] , \g5[5][3] , \g5[5][2] , \g5[5][1] , \g5[4][63] ,
         \g5[4][62] , \g5[4][61] , \g5[4][60] , \g5[4][59] , \g5[4][58] ,
         \g5[4][57] , \g5[4][56] , \g5[4][55] , \g5[4][54] , \g5[4][53] ,
         \g5[4][52] , \g5[4][51] , \g5[4][50] , \g5[4][49] , \g5[4][48] ,
         \g5[4][47] , \g5[4][46] , \g5[4][45] , \g5[4][44] , \g5[4][43] ,
         \g5[4][42] , \g5[4][41] , \g5[4][40] , \g5[4][39] , \g5[4][38] ,
         \g5[4][37] , \g5[4][36] , \g5[4][35] , \g5[4][34] , \g5[4][33] ,
         \g5[4][32] , \g5[4][31] , \g5[4][30] , \g5[4][29] , \g5[4][28] ,
         \g5[4][27] , \g5[4][26] , \g5[4][25] , \g5[4][24] , \g5[4][23] ,
         \g5[4][22] , \g5[4][21] , \g5[4][20] , \g5[4][19] , \g5[4][18] ,
         \g5[4][17] , \g5[4][16] , \g5[4][15] , \g5[4][14] , \g5[4][13] ,
         \g5[4][12] , \g5[4][11] , \g5[4][10] , \g5[4][9] , \g5[4][8] ,
         \g5[4][7] , \g5[4][6] , \g5[4][5] , \g5[4][4] , \g5[4][3] ,
         \g5[4][2] , \g5[4][1] , \g5[3][63] , \g5[3][62] , \g5[3][61] ,
         \g5[3][60] , \g5[3][59] , \g5[3][58] , \g5[3][57] , \g5[3][56] ,
         \g5[3][55] , \g5[3][54] , \g5[3][53] , \g5[3][52] , \g5[3][51] ,
         \g5[3][50] , \g5[3][49] , \g5[3][48] , \g5[3][47] , \g5[3][46] ,
         \g5[3][45] , \g5[3][44] , \g5[3][43] , \g5[3][42] , \g5[3][41] ,
         \g5[3][40] , \g5[3][39] , \g5[3][38] , \g5[3][37] , \g5[3][36] ,
         \g5[3][35] , \g5[3][34] , \g5[3][33] , \g5[3][32] , \g5[3][31] ,
         \g5[3][30] , \g5[3][29] , \g5[3][28] , \g5[3][27] , \g5[3][26] ,
         \g5[3][25] , \g5[3][24] , \g5[3][23] , \g5[3][22] , \g5[3][21] ,
         \g5[3][20] , \g5[3][19] , \g5[3][18] , \g5[3][17] , \g5[3][16] ,
         \g5[3][15] , \g5[3][14] , \g5[3][13] , \g5[3][12] , \g5[3][11] ,
         \g5[3][10] , \g5[3][9] , \g5[3][8] , \g5[3][7] , \g5[3][6] ,
         \g5[3][5] , \g5[3][4] , \g5[3][3] , \g5[3][2] , \g5[3][1] ,
         \g5[3][0] , \g5[2][63] , \g5[2][62] , \g5[2][61] , \g5[2][60] ,
         \g5[2][59] , \g5[2][58] , \g5[2][57] , \g5[2][56] , \g5[2][55] ,
         \g5[2][54] , \g5[2][53] , \g5[2][52] , \g5[2][51] , \g5[2][50] ,
         \g5[2][49] , \g5[2][48] , \g5[2][47] , \g5[2][46] , \g5[2][45] ,
         \g5[2][44] , \g5[2][43] , \g5[2][42] , \g5[2][41] , \g5[2][40] ,
         \g5[2][39] , \g5[2][38] , \g5[2][37] , \g5[2][36] , \g5[2][35] ,
         \g5[2][34] , \g5[2][33] , \g5[2][32] , \g5[2][31] , \g5[2][30] ,
         \g5[2][29] , \g5[2][28] , \g5[2][27] , \g5[2][26] , \g5[2][25] ,
         \g5[2][24] , \g5[2][23] , \g5[2][22] , \g5[2][21] , \g5[2][20] ,
         \g5[2][19] , \g5[2][18] , \g5[2][17] , \g5[2][16] , \g5[2][15] ,
         \g5[2][14] , \g5[2][13] , \g5[2][12] , \g5[2][11] , \g5[2][10] ,
         \g5[2][9] , \g5[2][8] , \g5[2][7] , \g5[2][6] , \g5[2][5] ,
         \g5[2][4] , \g5[2][3] , \g5[2][2] , \g5[2][1] , \g5[2][0] ,
         \g5[1][63] , \g5[1][62] , \g5[1][61] , \g5[1][60] , \g5[1][59] ,
         \g5[1][58] , \g5[1][57] , \g5[1][56] , \g5[1][55] , \g5[1][54] ,
         \g5[1][53] , \g5[1][52] , \g5[1][51] , \g5[1][50] , \g5[1][49] ,
         \g5[1][48] , \g5[1][47] , \g5[1][46] , \g5[1][45] , \g5[1][44] ,
         \g5[1][43] , \g5[1][42] , \g5[1][41] , \g5[1][40] , \g5[1][39] ,
         \g5[1][38] , \g5[1][37] , \g5[1][36] , \g5[1][35] , \g5[1][34] ,
         \g5[1][33] , \g5[1][32] , \g5[1][31] , \g5[1][30] , \g5[1][29] ,
         \g5[1][28] , \g5[1][27] , \g5[1][26] , \g5[1][25] , \g5[1][24] ,
         \g5[1][23] , \g5[1][22] , \g5[1][21] , \g5[1][20] , \g5[1][19] ,
         \g5[1][18] , \g5[1][17] , \g5[1][16] , \g5[1][15] , \g5[1][14] ,
         \g5[1][13] , \g5[1][12] , \g5[1][11] , \g5[1][10] , \g5[1][9] ,
         \g5[1][8] , \g5[1][7] , \g5[1][6] , \g5[1][5] , \g5[1][4] ,
         \g5[1][3] , \g5[1][2] , \g5[1][1] , \g5[1][0] , \g5[0][63] ,
         \g5[0][62] , \g5[0][61] , \g5[0][60] , \g5[0][59] , \g5[0][58] ,
         \g5[0][57] , \g5[0][56] , \g5[0][55] , \g5[0][54] , \g5[0][53] ,
         \g5[0][52] , \g5[0][51] , \g5[0][50] , \g5[0][49] , \g5[0][48] ,
         \g5[0][47] , \g5[0][46] , \g5[0][45] , \g5[0][44] , \g5[0][43] ,
         \g5[0][42] , \g5[0][41] , \g5[0][40] , \g5[0][39] , \g5[0][38] ,
         \g5[0][37] , \g5[0][36] , \g5[0][35] , \g5[0][34] , \g5[0][33] ,
         \g5[0][32] , \g5[0][31] , \g5[0][30] , \g5[0][29] , \g5[0][28] ,
         \g5[0][27] , \g5[0][26] , \g5[0][25] , \g5[0][24] , \g5[0][23] ,
         \g5[0][22] , \g5[0][21] , \g5[0][20] , \g5[0][19] , \g5[0][18] ,
         \g5[0][17] , \g5[0][16] , \g5[0][15] , \g5[0][14] , \g5[0][13] ,
         \g5[0][12] , \g5[0][11] , \g5[0][10] , \g5[0][9] , \g5[0][8] ,
         \g5[0][7] , \g5[0][6] , \g5[0][5] , \g5[0][4] , \g5[0][3] ,
         \g5[0][2] , \g5[0][1] , \g5[0][0] , \g6[5][63] , \g6[5][62] ,
         \g6[5][61] , \g6[5][60] , \g6[5][59] , \g6[5][58] , \g6[5][57] ,
         \g6[5][56] , \g6[5][55] , \g6[5][54] , \g6[5][53] , \g6[5][52] ,
         \g6[5][51] , \g6[5][50] , \g6[5][49] , \g6[5][48] , \g6[5][47] ,
         \g6[5][46] , \g6[5][45] , \g6[5][44] , \g6[5][43] , \g6[5][42] ,
         \g6[5][41] , \g6[5][40] , \g6[5][39] , \g6[5][38] , \g6[5][37] ,
         \g6[5][36] , \g6[5][35] , \g6[5][34] , \g6[5][33] , \g6[5][32] ,
         \g6[5][31] , \g6[5][30] , \g6[5][29] , \g6[5][28] , \g6[5][27] ,
         \g6[5][26] , \g6[5][25] , \g6[5][24] , \g6[5][23] , \g6[5][22] ,
         \g6[5][21] , \g6[5][20] , \g6[5][19] , \g6[5][18] , \g6[5][17] ,
         \g6[5][16] , \g6[5][15] , \g6[5][14] , \g6[5][13] , \g6[5][12] ,
         \g6[5][11] , \g6[5][10] , \g6[5][9] , \g6[5][8] , \g6[5][7] ,
         \g6[5][6] , \g6[5][5] , \g6[5][4] , \g6[5][3] , \g6[5][2] ,
         \g6[5][1] , \g6[4][63] , \g6[4][62] , \g6[4][61] , \g6[4][60] ,
         \g6[4][59] , \g6[4][58] , \g6[4][57] , \g6[4][56] , \g6[4][55] ,
         \g6[4][54] , \g6[4][53] , \g6[4][52] , \g6[4][51] , \g6[4][50] ,
         \g6[4][49] , \g6[4][48] , \g6[4][47] , \g6[4][46] , \g6[4][45] ,
         \g6[4][44] , \g6[4][43] , \g6[4][42] , \g6[4][41] , \g6[4][40] ,
         \g6[4][39] , \g6[4][38] , \g6[4][37] , \g6[4][36] , \g6[4][35] ,
         \g6[4][34] , \g6[4][33] , \g6[4][32] , \g6[4][31] , \g6[4][30] ,
         \g6[4][29] , \g6[4][28] , \g6[4][27] , \g6[4][26] , \g6[4][25] ,
         \g6[4][24] , \g6[4][23] , \g6[4][22] , \g6[4][21] , \g6[4][20] ,
         \g6[4][19] , \g6[4][18] , \g6[4][17] , \g6[4][16] , \g6[4][15] ,
         \g6[4][14] , \g6[4][13] , \g6[4][12] , \g6[4][11] , \g6[4][10] ,
         \g6[4][9] , \g6[4][8] , \g6[4][7] , \g6[4][6] , \g6[4][5] ,
         \g6[4][4] , \g6[4][3] , \g6[4][2] , \g6[4][1] , \g6[4][0] ,
         \g6[3][63] , \g6[3][62] , \g6[3][61] , \g6[3][60] , \g6[3][59] ,
         \g6[3][58] , \g6[3][57] , \g6[3][56] , \g6[3][55] , \g6[3][54] ,
         \g6[3][53] , \g6[3][52] , \g6[3][51] , \g6[3][50] , \g6[3][49] ,
         \g6[3][48] , \g6[3][47] , \g6[3][46] , \g6[3][45] , \g6[3][44] ,
         \g6[3][43] , \g6[3][42] , \g6[3][41] , \g6[3][40] , \g6[3][39] ,
         \g6[3][38] , \g6[3][37] , \g6[3][36] , \g6[3][35] , \g6[3][34] ,
         \g6[3][33] , \g6[3][32] , \g6[3][31] , \g6[3][30] , \g6[3][29] ,
         \g6[3][28] , \g6[3][27] , \g6[3][26] , \g6[3][25] , \g6[3][24] ,
         \g6[3][23] , \g6[3][22] , \g6[3][21] , \g6[3][20] , \g6[3][19] ,
         \g6[3][18] , \g6[3][17] , \g6[3][16] , \g6[3][15] , \g6[3][14] ,
         \g6[3][13] , \g6[3][12] , \g6[3][11] , \g6[3][10] , \g6[3][9] ,
         \g6[3][8] , \g6[3][7] , \g6[3][6] , \g6[3][5] , \g6[3][4] ,
         \g6[3][3] , \g6[3][2] , \g6[3][1] , \g6[2][63] , \g6[2][62] ,
         \g6[2][61] , \g6[2][60] , \g6[2][59] , \g6[2][58] , \g6[2][57] ,
         \g6[2][56] , \g6[2][55] , \g6[2][54] , \g6[2][53] , \g6[2][52] ,
         \g6[2][51] , \g6[2][50] , \g6[2][49] , \g6[2][48] , \g6[2][47] ,
         \g6[2][46] , \g6[2][45] , \g6[2][44] , \g6[2][43] , \g6[2][42] ,
         \g6[2][41] , \g6[2][40] , \g6[2][39] , \g6[2][38] , \g6[2][37] ,
         \g6[2][36] , \g6[2][35] , \g6[2][34] , \g6[2][33] , \g6[2][32] ,
         \g6[2][31] , \g6[2][30] , \g6[2][29] , \g6[2][28] , \g6[2][27] ,
         \g6[2][26] , \g6[2][25] , \g6[2][24] , \g6[2][23] , \g6[2][22] ,
         \g6[2][21] , \g6[2][20] , \g6[2][19] , \g6[2][18] , \g6[2][17] ,
         \g6[2][16] , \g6[2][15] , \g6[2][14] , \g6[2][13] , \g6[2][12] ,
         \g6[2][11] , \g6[2][10] , \g6[2][9] , \g6[2][8] , \g6[2][7] ,
         \g6[2][6] , \g6[2][5] , \g6[2][4] , \g6[2][3] , \g6[2][2] ,
         \g6[2][1] , \g6[2][0] , \g6[1][63] , \g6[1][62] , \g6[1][61] ,
         \g6[1][60] , \g6[1][59] , \g6[1][58] , \g6[1][57] , \g6[1][56] ,
         \g6[1][55] , \g6[1][54] , \g6[1][53] , \g6[1][52] , \g6[1][51] ,
         \g6[1][50] , \g6[1][49] , \g6[1][48] , \g6[1][47] , \g6[1][46] ,
         \g6[1][45] , \g6[1][44] , \g6[1][43] , \g6[1][42] , \g6[1][41] ,
         \g6[1][40] , \g6[1][39] , \g6[1][38] , \g6[1][37] , \g6[1][36] ,
         \g6[1][35] , \g6[1][34] , \g6[1][33] , \g6[1][32] , \g6[1][31] ,
         \g6[1][30] , \g6[1][29] , \g6[1][28] , \g6[1][27] , \g6[1][26] ,
         \g6[1][25] , \g6[1][24] , \g6[1][23] , \g6[1][22] , \g6[1][21] ,
         \g6[1][20] , \g6[1][19] , \g6[1][18] , \g6[1][17] , \g6[1][16] ,
         \g6[1][15] , \g6[1][14] , \g6[1][13] , \g6[1][12] , \g6[1][11] ,
         \g6[1][10] , \g6[1][9] , \g6[1][8] , \g6[1][7] , \g6[1][6] ,
         \g6[1][5] , \g6[1][4] , \g6[1][3] , \g6[1][2] , \g6[1][1] ,
         \g6[0][63] , \g6[0][62] , \g6[0][61] , \g6[0][60] , \g6[0][59] ,
         \g6[0][58] , \g6[0][57] , \g6[0][56] , \g6[0][55] , \g6[0][54] ,
         \g6[0][53] , \g6[0][52] , \g6[0][51] , \g6[0][50] , \g6[0][49] ,
         \g6[0][48] , \g6[0][47] , \g6[0][46] , \g6[0][45] , \g6[0][44] ,
         \g6[0][43] , \g6[0][42] , \g6[0][41] , \g6[0][40] , \g6[0][39] ,
         \g6[0][38] , \g6[0][37] , \g6[0][36] , \g6[0][35] , \g6[0][34] ,
         \g6[0][33] , \g6[0][32] , \g6[0][31] , \g6[0][30] , \g6[0][29] ,
         \g6[0][28] , \g6[0][27] , \g6[0][26] , \g6[0][25] , \g6[0][24] ,
         \g6[0][23] , \g6[0][22] , \g6[0][21] , \g6[0][20] , \g6[0][19] ,
         \g6[0][18] , \g6[0][17] , \g6[0][16] , \g6[0][15] , \g6[0][14] ,
         \g6[0][13] , \g6[0][12] , \g6[0][11] , \g6[0][10] , \g6[0][9] ,
         \g6[0][8] , \g6[0][7] , \g6[0][6] , \g6[0][5] , \g6[0][4] ,
         \g6[0][3] , \g6[0][2] , \g6[0][1] , \g6[0][0] , \g7[3][63] ,
         \g7[3][62] , \g7[3][61] , \g7[3][60] , \g7[3][59] , \g7[3][58] ,
         \g7[3][57] , \g7[3][56] , \g7[3][55] , \g7[3][54] , \g7[3][53] ,
         \g7[3][52] , \g7[3][51] , \g7[3][50] , \g7[3][49] , \g7[3][48] ,
         \g7[3][47] , \g7[3][46] , \g7[3][45] , \g7[3][44] , \g7[3][43] ,
         \g7[3][42] , \g7[3][41] , \g7[3][40] , \g7[3][39] , \g7[3][38] ,
         \g7[3][37] , \g7[3][36] , \g7[3][35] , \g7[3][34] , \g7[3][33] ,
         \g7[3][32] , \g7[3][31] , \g7[3][30] , \g7[3][29] , \g7[3][28] ,
         \g7[3][27] , \g7[3][26] , \g7[3][25] , \g7[3][24] , \g7[3][23] ,
         \g7[3][22] , \g7[3][21] , \g7[3][20] , \g7[3][19] , \g7[3][18] ,
         \g7[3][17] , \g7[3][16] , \g7[3][15] , \g7[3][14] , \g7[3][13] ,
         \g7[3][12] , \g7[3][11] , \g7[3][10] , \g7[3][9] , \g7[3][8] ,
         \g7[3][7] , \g7[3][6] , \g7[3][5] , \g7[3][4] , \g7[3][3] ,
         \g7[3][2] , \g7[3][1] , \g7[2][63] , \g7[2][62] , \g7[2][61] ,
         \g7[2][60] , \g7[2][59] , \g7[2][58] , \g7[2][57] , \g7[2][56] ,
         \g7[2][55] , \g7[2][54] , \g7[2][53] , \g7[2][52] , \g7[2][51] ,
         \g7[2][50] , \g7[2][49] , \g7[2][48] , \g7[2][47] , \g7[2][46] ,
         \g7[2][45] , \g7[2][44] , \g7[2][43] , \g7[2][42] , \g7[2][41] ,
         \g7[2][40] , \g7[2][39] , \g7[2][38] , \g7[2][37] , \g7[2][36] ,
         \g7[2][35] , \g7[2][34] , \g7[2][33] , \g7[2][32] , \g7[2][31] ,
         \g7[2][30] , \g7[2][29] , \g7[2][28] , \g7[2][27] , \g7[2][26] ,
         \g7[2][25] , \g7[2][24] , \g7[2][23] , \g7[2][22] , \g7[2][21] ,
         \g7[2][20] , \g7[2][19] , \g7[2][18] , \g7[2][17] , \g7[2][16] ,
         \g7[2][15] , \g7[2][14] , \g7[2][13] , \g7[2][12] , \g7[2][11] ,
         \g7[2][10] , \g7[2][9] , \g7[2][8] , \g7[2][7] , \g7[2][6] ,
         \g7[2][5] , \g7[2][4] , \g7[2][3] , \g7[2][2] , \g7[2][1] ,
         \g7[2][0] , \g7[1][63] , \g7[1][62] , \g7[1][61] , \g7[1][60] ,
         \g7[1][59] , \g7[1][58] , \g7[1][57] , \g7[1][56] , \g7[1][55] ,
         \g7[1][54] , \g7[1][53] , \g7[1][52] , \g7[1][51] , \g7[1][50] ,
         \g7[1][49] , \g7[1][48] , \g7[1][47] , \g7[1][46] , \g7[1][45] ,
         \g7[1][44] , \g7[1][43] , \g7[1][42] , \g7[1][41] , \g7[1][40] ,
         \g7[1][39] , \g7[1][38] , \g7[1][37] , \g7[1][36] , \g7[1][35] ,
         \g7[1][34] , \g7[1][33] , \g7[1][32] , \g7[1][31] , \g7[1][30] ,
         \g7[1][29] , \g7[1][28] , \g7[1][27] , \g7[1][26] , \g7[1][25] ,
         \g7[1][24] , \g7[1][23] , \g7[1][22] , \g7[1][21] , \g7[1][20] ,
         \g7[1][19] , \g7[1][18] , \g7[1][17] , \g7[1][16] , \g7[1][15] ,
         \g7[1][14] , \g7[1][13] , \g7[1][12] , \g7[1][11] , \g7[1][10] ,
         \g7[1][9] , \g7[1][8] , \g7[1][7] , \g7[1][6] , \g7[1][5] ,
         \g7[1][4] , \g7[1][3] , \g7[1][2] , \g7[1][1] , \g7[0][63] ,
         \g7[0][62] , \g7[0][61] , \g7[0][60] , \g7[0][59] , \g7[0][58] ,
         \g7[0][57] , \g7[0][56] , \g7[0][55] , \g7[0][54] , \g7[0][53] ,
         \g7[0][52] , \g7[0][51] , \g7[0][50] , \g7[0][49] , \g7[0][48] ,
         \g7[0][47] , \g7[0][46] , \g7[0][45] , \g7[0][44] , \g7[0][43] ,
         \g7[0][42] , \g7[0][41] , \g7[0][40] , \g7[0][39] , \g7[0][38] ,
         \g7[0][37] , \g7[0][36] , \g7[0][35] , \g7[0][34] , \g7[0][33] ,
         \g7[0][32] , \g7[0][31] , \g7[0][30] , \g7[0][29] , \g7[0][28] ,
         \g7[0][27] , \g7[0][26] , \g7[0][25] , \g7[0][24] , \g7[0][23] ,
         \g7[0][22] , \g7[0][21] , \g7[0][20] , \g7[0][19] , \g7[0][18] ,
         \g7[0][17] , \g7[0][16] , \g7[0][15] , \g7[0][14] , \g7[0][13] ,
         \g7[0][12] , \g7[0][11] , \g7[0][10] , \g7[0][9] , \g7[0][8] ,
         \g7[0][7] , \g7[0][6] , \g7[0][5] , \g7[0][4] , \g7[0][3] ,
         \g7[0][2] , \g7[0][1] , \g7[0][0] , \g8[1][63] , \g8[1][62] ,
         \g8[1][61] , \g8[1][60] , \g8[1][59] , \g8[1][58] , \g8[1][57] ,
         \g8[1][56] , \g8[1][55] , \g8[1][54] , \g8[1][53] , \g8[1][52] ,
         \g8[1][51] , \g8[1][50] , \g8[1][49] , \g8[1][48] , \g8[1][47] ,
         \g8[1][46] , \g8[1][45] , \g8[1][44] , \g8[1][43] , \g8[1][42] ,
         \g8[1][41] , \g8[1][40] , \g8[1][39] , \g8[1][38] , \g8[1][37] ,
         \g8[1][36] , \g8[1][35] , \g8[1][34] , \g8[1][33] , \g8[1][32] ,
         \g8[1][31] , \g8[1][30] , \g8[1][29] , \g8[1][28] , \g8[1][27] ,
         \g8[1][26] , \g8[1][25] , \g8[1][24] , \g8[1][23] , \g8[1][22] ,
         \g8[1][21] , \g8[1][20] , \g8[1][19] , \g8[1][18] , \g8[1][17] ,
         \g8[1][16] , \g8[1][15] , \g8[1][14] , \g8[1][13] , \g8[1][12] ,
         \g8[1][11] , \g8[1][10] , \g8[1][9] , \g8[1][8] , \g8[1][7] ,
         \g8[1][6] , \g8[1][5] , \g8[1][4] , \g8[1][3] , \g8[1][2] ,
         \g8[1][1] , \g8[0][63] , \g8[0][62] , \g8[0][61] , \g8[0][60] ,
         \g8[0][59] , \g8[0][58] , \g8[0][57] , \g8[0][56] , \g8[0][55] ,
         \g8[0][54] , \g8[0][53] , \g8[0][52] , \g8[0][51] , \g8[0][50] ,
         \g8[0][49] , \g8[0][48] , \g8[0][47] , \g8[0][46] , \g8[0][45] ,
         \g8[0][44] , \g8[0][43] , \g8[0][42] , \g8[0][41] , \g8[0][40] ,
         \g8[0][39] , \g8[0][38] , \g8[0][37] , \g8[0][36] , \g8[0][35] ,
         \g8[0][34] , \g8[0][33] , \g8[0][32] , \g8[0][31] , \g8[0][30] ,
         \g8[0][29] , \g8[0][28] , \g8[0][27] , \g8[0][26] , \g8[0][25] ,
         \g8[0][24] , \g8[0][23] , \g8[0][22] , \g8[0][21] , \g8[0][20] ,
         \g8[0][19] , \g8[0][18] , \g8[0][17] , \g8[0][16] , \g8[0][15] ,
         \g8[0][14] , \g8[0][13] , \g8[0][12] , \g8[0][11] , \g8[0][10] ,
         \g8[0][9] , \g8[0][8] , \g8[0][7] , \g8[0][6] , \g8[0][5] ,
         \g8[0][4] , \g8[0][3] , \g8[0][2] , \g8[0][1] , \g8[0][0] ,
         \g9[1][63] , \g9[1][62] , \g9[1][61] , \g9[1][60] , \g9[1][59] ,
         \g9[1][58] , \g9[1][57] , \g9[1][56] , \g9[1][55] , \g9[1][54] ,
         \g9[1][53] , \g9[1][52] , \g9[1][51] , \g9[1][50] , \g9[1][49] ,
         \g9[1][48] , \g9[1][47] , \g9[1][46] , \g9[1][45] , \g9[1][44] ,
         \g9[1][43] , \g9[1][42] , \g9[1][41] , \g9[1][40] , \g9[1][39] ,
         \g9[1][38] , \g9[1][37] , \g9[1][36] , \g9[1][35] , \g9[1][34] ,
         \g9[1][33] , \g9[1][32] , \g9[1][31] , \g9[1][30] , \g9[1][29] ,
         \g9[1][28] , \g9[1][27] , \g9[1][26] , \g9[1][25] , \g9[1][24] ,
         \g9[1][23] , \g9[1][22] , \g9[1][21] , \g9[1][20] , \g9[1][19] ,
         \g9[1][18] , \g9[1][17] , \g9[1][16] , \g9[1][15] , \g9[1][14] ,
         \g9[1][13] , \g9[1][12] , \g9[1][11] , \g9[1][10] , \g9[1][9] ,
         \g9[1][8] , \g9[1][7] , \g9[1][6] , \g9[1][5] , \g9[1][4] ,
         \g9[1][3] , \g9[1][2] , \g9[1][1] , \g9[0][63] , \g9[0][62] ,
         \g9[0][61] , \g9[0][60] , \g9[0][59] , \g9[0][58] , \g9[0][57] ,
         \g9[0][56] , \g9[0][55] , \g9[0][54] , \g9[0][53] , \g9[0][52] ,
         \g9[0][51] , \g9[0][50] , \g9[0][49] , \g9[0][48] , \g9[0][47] ,
         \g9[0][46] , \g9[0][45] , \g9[0][44] , \g9[0][43] , \g9[0][42] ,
         \g9[0][41] , \g9[0][40] , \g9[0][39] , \g9[0][38] , \g9[0][37] ,
         \g9[0][36] , \g9[0][35] , \g9[0][34] , \g9[0][33] , \g9[0][32] ,
         \g9[0][31] , \g9[0][30] , \g9[0][29] , \g9[0][28] , \g9[0][27] ,
         \g9[0][26] , \g9[0][25] , \g9[0][24] , \g9[0][23] , \g9[0][22] ,
         \g9[0][21] , \g9[0][20] , \g9[0][19] , \g9[0][18] , \g9[0][17] ,
         \g9[0][16] , \g9[0][15] , \g9[0][14] , \g9[0][13] , \g9[0][12] ,
         \g9[0][11] , \g9[0][10] , \g9[0][9] , \g9[0][8] , \g9[0][7] ,
         \g9[0][6] , \g9[0][5] , \g9[0][4] , \g9[0][3] , \g9[0][2] ,
         \g9[0][1] , \g9[0][0] , \g10[1][63] , \g10[1][62] , \g10[1][61] ,
         \g10[1][60] , \g10[1][59] , \g10[1][58] , \g10[1][57] , \g10[1][56] ,
         \g10[1][55] , \g10[1][54] , \g10[1][53] , \g10[1][52] , \g10[1][51] ,
         \g10[1][50] , \g10[1][49] , \g10[1][48] , \g10[1][47] , \g10[1][46] ,
         \g10[1][45] , \g10[1][44] , \g10[1][43] , \g10[1][42] , \g10[1][41] ,
         \g10[1][40] , \g10[1][39] , \g10[1][38] , \g10[1][37] , \g10[1][36] ,
         \g10[1][35] , \g10[1][34] , \g10[1][33] , \g10[1][32] , \g10[1][31] ,
         \g10[1][30] , \g10[1][29] , \g10[1][28] , \g10[1][27] , \g10[1][26] ,
         \g10[1][25] , \g10[1][24] , \g10[1][23] , \g10[1][22] , \g10[1][21] ,
         \g10[1][20] , \g10[1][19] , \g10[1][18] , \g10[1][17] , \g10[1][16] ,
         \g10[1][15] , \g10[1][14] , \g10[1][13] , \g10[1][12] , \g10[1][11] ,
         \g10[1][10] , \g10[1][9] , \g10[1][8] , \g10[1][7] , \g10[1][6] ,
         \g10[1][5] , \g10[1][4] , \g10[1][3] , \g10[1][2] , \g10[1][1] ,
         \g10[0][63] , \g10[0][62] , \g10[0][61] , \g10[0][60] , \g10[0][59] ,
         \g10[0][58] , \g10[0][57] , \g10[0][56] , \g10[0][55] , \g10[0][54] ,
         \g10[0][53] , \g10[0][52] , \g10[0][51] , \g10[0][50] , \g10[0][49] ,
         \g10[0][48] , \g10[0][47] , \g10[0][46] , \g10[0][45] , \g10[0][44] ,
         \g10[0][43] , \g10[0][42] , \g10[0][41] , \g10[0][40] , \g10[0][39] ,
         \g10[0][38] , \g10[0][37] , \g10[0][36] , \g10[0][35] , \g10[0][34] ,
         \g10[0][33] , \g10[0][32] , \g10[0][31] , \g10[0][30] , \g10[0][29] ,
         \g10[0][28] , \g10[0][27] , \g10[0][26] , \g10[0][25] , \g10[0][24] ,
         \g10[0][23] , \g10[0][22] , \g10[0][21] , \g10[0][20] , \g10[0][19] ,
         \g10[0][18] , \g10[0][17] , \g10[0][16] , \g10[0][15] , \g10[0][14] ,
         \g10[0][13] , \g10[0][12] , \g10[0][11] , \g10[0][10] , \g10[0][9] ,
         \g10[0][8] , \g10[0][7] , \g10[0][6] , \g10[0][5] , \g10[0][4] ,
         \g10[0][3] , \g10[0][2] , \g10[0][1] , \g10[0][0] , N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445;
  wire   [31:0] A_reg;
  wire   [31:0] B_reg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61;

  DFF_X1 \A_reg_reg[31]  ( .D(N66), .CK(clk), .Q(A_reg[31]) );
  DFF_X1 \A_reg_reg[30]  ( .D(N65), .CK(clk), .Q(A_reg[30]), .QN(n95) );
  DFF_X1 \A_reg_reg[29]  ( .D(N64), .CK(clk), .Q(A_reg[29]), .QN(n96) );
  DFF_X1 \A_reg_reg[28]  ( .D(N63), .CK(clk), .Q(A_reg[28]), .QN(n97) );
  DFF_X1 \A_reg_reg[27]  ( .D(N62), .CK(clk), .Q(A_reg[27]), .QN(n98) );
  DFF_X1 \A_reg_reg[26]  ( .D(N61), .CK(clk), .Q(A_reg[26]), .QN(n99) );
  DFF_X1 \A_reg_reg[25]  ( .D(N60), .CK(clk), .Q(A_reg[25]), .QN(n100) );
  DFF_X1 \A_reg_reg[24]  ( .D(N59), .CK(clk), .Q(A_reg[24]), .QN(n94) );
  DFF_X1 \A_reg_reg[23]  ( .D(N58), .CK(clk), .Q(A_reg[23]), .QN(n78) );
  DFF_X1 \A_reg_reg[22]  ( .D(N57), .CK(clk), .Q(A_reg[22]), .QN(n79) );
  DFF_X1 \A_reg_reg[21]  ( .D(N56), .CK(clk), .Q(A_reg[21]), .QN(n77) );
  DFF_X1 \A_reg_reg[20]  ( .D(N55), .CK(clk), .Q(A_reg[20]), .QN(n71) );
  DFF_X1 \A_reg_reg[19]  ( .D(N54), .CK(clk), .Q(A_reg[19]), .QN(n74) );
  DFF_X1 \A_reg_reg[18]  ( .D(N53), .CK(clk), .Q(A_reg[18]), .QN(n70) );
  DFF_X1 \A_reg_reg[17]  ( .D(N52), .CK(clk), .Q(A_reg[17]), .QN(n76) );
  DFF_X1 \A_reg_reg[16]  ( .D(N51), .CK(clk), .Q(A_reg[16]), .QN(n75) );
  DFF_X1 \A_reg_reg[15]  ( .D(N50), .CK(clk), .Q(A_reg[15]), .QN(n73) );
  DFF_X1 \A_reg_reg[14]  ( .D(N49), .CK(clk), .Q(A_reg[14]), .QN(n72) );
  DFF_X1 \A_reg_reg[13]  ( .D(N48), .CK(clk), .Q(A_reg[13]), .QN(n69) );
  DFF_X1 \A_reg_reg[12]  ( .D(N47), .CK(clk), .Q(A_reg[12]), .QN(n90) );
  DFF_X1 \A_reg_reg[11]  ( .D(N46), .CK(clk), .Q(A_reg[11]), .QN(n91) );
  DFF_X1 \A_reg_reg[10]  ( .D(N45), .CK(clk), .Q(A_reg[10]), .QN(n66) );
  DFF_X1 \A_reg_reg[9]  ( .D(N44), .CK(clk), .Q(A_reg[9]), .QN(n67) );
  DFF_X1 \A_reg_reg[8]  ( .D(N43), .CK(clk), .Q(A_reg[8]), .QN(n117) );
  DFF_X1 \A_reg_reg[7]  ( .D(N42), .CK(clk), .Q(A_reg[7]), .QN(n141) );
  DFF_X1 \A_reg_reg[6]  ( .D(N41), .CK(clk), .Q(A_reg[6]), .QN(n139) );
  DFF_X1 \A_reg_reg[5]  ( .D(N40), .CK(clk), .Q(A_reg[5]), .QN(n128) );
  DFF_X1 \A_reg_reg[4]  ( .D(N39), .CK(clk), .Q(A_reg[4]), .QN(n138) );
  DFF_X1 \A_reg_reg[3]  ( .D(N38), .CK(clk), .Q(A_reg[3]), .QN(n140) );
  DFF_X1 \A_reg_reg[2]  ( .D(N37), .CK(clk), .Q(A_reg[2]), .QN(n121) );
  DFF_X1 \A_reg_reg[1]  ( .D(N36), .CK(clk), .Q(A_reg[1]), .QN(n124) );
  DFF_X1 \A_reg_reg[0]  ( .D(N35), .CK(clk), .Q(A_reg[0]), .QN(n120) );
  DFF_X1 \B_reg_reg[31]  ( .D(N98), .CK(clk), .Q(B_reg[31]) );
  DFF_X1 \B_reg_reg[30]  ( .D(N97), .CK(clk), .Q(B_reg[30]), .QN(n106) );
  DFF_X1 \B_reg_reg[29]  ( .D(N96), .CK(clk), .Q(B_reg[29]), .QN(n105) );
  DFF_X1 \B_reg_reg[28]  ( .D(N95), .CK(clk), .Q(B_reg[28]), .QN(n107) );
  DFF_X1 \B_reg_reg[27]  ( .D(N94), .CK(clk), .Q(B_reg[27]), .QN(n108) );
  DFF_X1 \B_reg_reg[26]  ( .D(N93), .CK(clk), .Q(B_reg[26]), .QN(n101) );
  DFF_X1 \B_reg_reg[25]  ( .D(N92), .CK(clk), .Q(B_reg[25]), .QN(n102) );
  DFF_X1 \B_reg_reg[24]  ( .D(N91), .CK(clk), .Q(B_reg[24]), .QN(n103) );
  DFF_X1 \B_reg_reg[23]  ( .D(N90), .CK(clk), .Q(B_reg[23]), .QN(n104) );
  DFF_X1 \B_reg_reg[22]  ( .D(N89), .CK(clk), .Q(B_reg[22]), .QN(n80) );
  DFF_X1 \B_reg_reg[21]  ( .D(N88), .CK(clk), .Q(B_reg[21]), .QN(n82) );
  DFF_X1 \B_reg_reg[20]  ( .D(N87), .CK(clk), .Q(B_reg[20]), .QN(n81) );
  DFF_X1 \B_reg_reg[19]  ( .D(N86), .CK(clk), .Q(B_reg[19]), .QN(n83) );
  DFF_X1 \B_reg_reg[18]  ( .D(N85), .CK(clk), .Q(B_reg[18]), .QN(n85) );
  DFF_X1 \B_reg_reg[17]  ( .D(N84), .CK(clk), .Q(B_reg[17]), .QN(n84) );
  DFF_X1 \B_reg_reg[16]  ( .D(N83), .CK(clk), .Q(B_reg[16]), .QN(n86) );
  DFF_X1 \B_reg_reg[15]  ( .D(N82), .CK(clk), .Q(B_reg[15]), .QN(n87) );
  DFF_X1 \B_reg_reg[14]  ( .D(N81), .CK(clk), .Q(B_reg[14]), .QN(n88) );
  DFF_X1 \B_reg_reg[13]  ( .D(N80), .CK(clk), .Q(B_reg[13]), .QN(n89) );
  DFF_X1 \B_reg_reg[12]  ( .D(N79), .CK(clk), .Q(B_reg[12]), .QN(n93) );
  DFF_X1 \B_reg_reg[11]  ( .D(N78), .CK(clk), .Q(B_reg[11]), .QN(n92) );
  DFF_X1 \B_reg_reg[10]  ( .D(N77), .CK(clk), .Q(B_reg[10]), .QN(n112) );
  DFF_X1 \B_reg_reg[9]  ( .D(N76), .CK(clk), .Q(B_reg[9]), .QN(n115) );
  DFF_X1 \B_reg_reg[8]  ( .D(N75), .CK(clk), .Q(B_reg[8]), .QN(n68) );
  DFF_X1 \B_reg_reg[7]  ( .D(N74), .CK(clk), .Q(B_reg[7]), .QN(n119) );
  DFF_X1 \B_reg_reg[6]  ( .D(N73), .CK(clk), .Q(B_reg[6]), .QN(n125) );
  DFF_X1 \B_reg_reg[5]  ( .D(N72), .CK(clk), .Q(B_reg[5]), .QN(n122) );
  DFF_X1 \B_reg_reg[4]  ( .D(N71), .CK(clk), .Q(B_reg[4]), .QN(n130) );
  DFF_X1 \B_reg_reg[3]  ( .D(N70), .CK(clk), .Q(B_reg[3]), .QN(n133) );
  DFF_X1 \B_reg_reg[2]  ( .D(N69), .CK(clk), .Q(B_reg[2]), .QN(n118) );
  DFF_X1 \B_reg_reg[1]  ( .D(N68), .CK(clk), .Q(B_reg[1]), .QN(n131) );
  DFF_X1 \B_reg_reg[0]  ( .D(N67), .CK(clk), .Q(B_reg[0]), .QN(n132) );
  DFF_X1 \out_reg[62]  ( .D(N257), .CK(clk), .Q(out[62]) );
  DFF_X1 \out_reg[61]  ( .D(N256), .CK(clk), .Q(out[61]) );
  DFF_X1 \out_reg[60]  ( .D(N255), .CK(clk), .Q(out[60]) );
  DFF_X1 \out_reg[59]  ( .D(N254), .CK(clk), .Q(out[59]) );
  DFF_X1 \out_reg[58]  ( .D(N253), .CK(clk), .Q(out[58]) );
  DFF_X1 \out_reg[57]  ( .D(N252), .CK(clk), .Q(out[57]) );
  DFF_X1 \out_reg[56]  ( .D(N251), .CK(clk), .Q(out[56]) );
  DFF_X1 \out_reg[55]  ( .D(N250), .CK(clk), .Q(out[55]) );
  DFF_X1 \out_reg[54]  ( .D(N249), .CK(clk), .Q(out[54]) );
  DFF_X1 \out_reg[53]  ( .D(N248), .CK(clk), .Q(out[53]) );
  DFF_X1 \out_reg[52]  ( .D(N247), .CK(clk), .Q(out[52]) );
  DFF_X1 \out_reg[51]  ( .D(N246), .CK(clk), .Q(out[51]) );
  DFF_X1 \out_reg[50]  ( .D(N245), .CK(clk), .Q(out[50]) );
  DFF_X1 \out_reg[49]  ( .D(N244), .CK(clk), .Q(out[49]) );
  DFF_X1 \out_reg[48]  ( .D(N243), .CK(clk), .Q(out[48]) );
  DFF_X1 \out_reg[47]  ( .D(N242), .CK(clk), .Q(out[47]) );
  DFF_X1 \out_reg[46]  ( .D(N241), .CK(clk), .Q(out[46]) );
  DFF_X1 \out_reg[45]  ( .D(N240), .CK(clk), .Q(out[45]) );
  DFF_X1 \out_reg[44]  ( .D(N239), .CK(clk), .Q(out[44]) );
  DFF_X1 \out_reg[43]  ( .D(N238), .CK(clk), .Q(out[43]) );
  DFF_X1 \out_reg[42]  ( .D(N237), .CK(clk), .Q(out[42]) );
  DFF_X1 \out_reg[41]  ( .D(N236), .CK(clk), .Q(out[41]) );
  DFF_X1 \out_reg[40]  ( .D(N235), .CK(clk), .Q(out[40]) );
  DFF_X1 \out_reg[39]  ( .D(N234), .CK(clk), .Q(out[39]) );
  DFF_X1 \out_reg[38]  ( .D(N233), .CK(clk), .Q(out[38]) );
  DFF_X1 \out_reg[37]  ( .D(N232), .CK(clk), .Q(out[37]) );
  DFF_X1 \out_reg[36]  ( .D(N231), .CK(clk), .Q(out[36]) );
  DFF_X1 \out_reg[35]  ( .D(N230), .CK(clk), .Q(out[35]) );
  DFF_X1 \out_reg[34]  ( .D(N229), .CK(clk), .Q(out[34]) );
  DFF_X1 \out_reg[33]  ( .D(N228), .CK(clk), .Q(out[33]) );
  DFF_X1 \out_reg[32]  ( .D(N227), .CK(clk), .Q(out[32]) );
  DFF_X1 \out_reg[31]  ( .D(N226), .CK(clk), .Q(out[31]) );
  DFF_X1 \out_reg[30]  ( .D(N225), .CK(clk), .Q(out[30]) );
  DFF_X1 \out_reg[29]  ( .D(N224), .CK(clk), .Q(out[29]) );
  DFF_X1 \out_reg[28]  ( .D(N223), .CK(clk), .Q(out[28]) );
  DFF_X1 \out_reg[27]  ( .D(N222), .CK(clk), .Q(out[27]) );
  DFF_X1 \out_reg[26]  ( .D(N221), .CK(clk), .Q(out[26]) );
  DFF_X1 \out_reg[25]  ( .D(N220), .CK(clk), .Q(out[25]) );
  DFF_X1 \out_reg[24]  ( .D(N219), .CK(clk), .Q(out[24]) );
  DFF_X1 \out_reg[23]  ( .D(N218), .CK(clk), .Q(out[23]) );
  DFF_X1 \out_reg[22]  ( .D(N217), .CK(clk), .Q(out[22]) );
  DFF_X1 \out_reg[21]  ( .D(N216), .CK(clk), .Q(out[21]) );
  DFF_X1 \out_reg[20]  ( .D(N215), .CK(clk), .Q(out[20]) );
  DFF_X1 \out_reg[19]  ( .D(N214), .CK(clk), .Q(out[19]) );
  DFF_X1 \out_reg[18]  ( .D(N213), .CK(clk), .Q(out[18]) );
  DFF_X1 \out_reg[17]  ( .D(N212), .CK(clk), .Q(out[17]) );
  DFF_X1 \out_reg[16]  ( .D(N211), .CK(clk), .Q(out[16]) );
  DFF_X1 \out_reg[15]  ( .D(N210), .CK(clk), .Q(out[15]) );
  DFF_X1 \out_reg[14]  ( .D(N209), .CK(clk), .Q(out[14]) );
  DFF_X1 \out_reg[13]  ( .D(N208), .CK(clk), .Q(out[13]) );
  DFF_X1 \out_reg[12]  ( .D(N207), .CK(clk), .Q(out[12]) );
  DFF_X1 \out_reg[11]  ( .D(N206), .CK(clk), .Q(out[11]) );
  DFF_X1 \out_reg[10]  ( .D(N205), .CK(clk), .Q(out[10]) );
  DFF_X1 \out_reg[9]  ( .D(N204), .CK(clk), .Q(out[9]) );
  DFF_X1 \out_reg[8]  ( .D(N203), .CK(clk), .Q(out[8]) );
  DFF_X1 \out_reg[7]  ( .D(N202), .CK(clk), .Q(out[7]) );
  DFF_X1 \out_reg[6]  ( .D(N201), .CK(clk), .Q(out[6]) );
  DFF_X1 \out_reg[5]  ( .D(N200), .CK(clk), .Q(out[5]) );
  DFF_X1 \out_reg[4]  ( .D(N199), .CK(clk), .Q(out[4]) );
  DFF_X1 \out_reg[3]  ( .D(N198), .CK(clk), .Q(out[3]) );
  DFF_X1 \out_reg[2]  ( .D(N197), .CK(clk), .Q(out[2]) );
  DFF_X1 \out_reg[1]  ( .D(N196), .CK(clk), .Q(out[1]) );
  DFF_X1 \out_reg[0]  ( .D(N195), .CK(clk), .Q(out[0]) );
  FullAdder \level1[0].x6  ( .a({n410, n410, n410, n410, n410, n410, n410, 
        n410, n410, n409, n409, n409, n409, n409, n409, n409, n409, n409, n409, 
        n409, n409, n408, n408, n408, n408, n408, n408, n408, n408, n408, n408, 
        n408, n408, \p[0][30] , \p[0][29] , \p[0][28] , \p[0][27] , \p[0][26] , 
        \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] , \p[0][21] , \p[0][20] , 
        \p[0][19] , \p[0][18] , \p[0][17] , \p[0][16] , \p[0][15] , \p[0][14] , 
        \p[0][13] , \p[0][12] , \p[0][11] , \p[0][10] , \p[0][9] , \p[0][8] , 
        \p[0][7] , \p[0][6] , \p[0][5] , \p[0][4] , \p[0][3] , \p[0][2] , 
        \p[0][1] , \p[0][0] }), .b({n413, n413, n413, n413, n413, n413, n413, 
        n413, n412, n412, n412, n412, n412, n412, n412, n412, n412, n412, n412, 
        n412, n411, n411, n411, n411, n411, n411, n411, n411, n411, n411, n411, 
        n411, \p[1][31] , \p[1][30] , \p[1][29] , \p[1][28] , \p[1][27] , 
        \p[1][26] , \p[1][25] , \p[1][24] , \p[1][23] , \p[1][22] , \p[1][21] , 
        \p[1][20] , \p[1][19] , \p[1][18] , \p[1][17] , \p[1][16] , \p[1][15] , 
        \p[1][14] , \p[1][13] , \p[1][12] , \p[1][11] , \p[1][10] , \p[1][9] , 
        \p[1][8] , \p[1][7] , \p[1][6] , \p[1][5] , \p[1][4] , \p[1][3] , 
        \p[1][2] , \p[1][1] , 1'b0}), .cin({n416, n416, n416, n416, n416, n416, 
        n416, n415, n415, n415, n415, n415, n415, n415, n415, n415, n415, n415, 
        n415, n414, n414, n414, n414, n414, n414, n414, n414, n414, n414, n414, 
        n414, \p[2][32] , \p[2][31] , \p[2][30] , \p[2][29] , \p[2][28] , 
        \p[2][27] , \p[2][26] , \p[2][25] , \p[2][24] , \p[2][23] , \p[2][22] , 
        \p[2][21] , \p[2][20] , \p[2][19] , \p[2][18] , \p[2][17] , \p[2][16] , 
        \p[2][15] , \p[2][14] , \p[2][13] , \p[2][12] , \p[2][11] , \p[2][10] , 
        \p[2][9] , \p[2][8] , \p[2][7] , \p[2][6] , \p[2][5] , \p[2][4] , 
        \p[2][3] , \p[2][2] , 1'b0, 1'b0}), .sum({\g[0][63] , \g[0][62] , 
        \g[0][61] , \g[0][60] , \g[0][59] , \g[0][58] , \g[0][57] , \g[0][56] , 
        \g[0][55] , \g[0][54] , \g[0][53] , \g[0][52] , \g[0][51] , \g[0][50] , 
        \g[0][49] , \g[0][48] , \g[0][47] , \g[0][46] , \g[0][45] , \g[0][44] , 
        \g[0][43] , \g[0][42] , \g[0][41] , \g[0][40] , \g[0][39] , \g[0][38] , 
        \g[0][37] , \g[0][36] , \g[0][35] , \g[0][34] , \g[0][33] , \g[0][32] , 
        \g[0][31] , \g[0][30] , \g[0][29] , \g[0][28] , \g[0][27] , \g[0][26] , 
        \g[0][25] , \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , 
        \g[0][19] , \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] , 
        \g[0][13] , \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] , 
        \g[0][7] , \g[0][6] , \g[0][5] , \g[0][4] , \g[0][3] , \g[0][2] , 
        \g[0][1] , \g[0][0] }), .cout({\g[21][63] , \g[21][62] , \g[21][61] , 
        \g[21][60] , \g[21][59] , \g[21][58] , \g[21][57] , \g[21][56] , 
        \g[21][55] , \g[21][54] , \g[21][53] , \g[21][52] , \g[21][51] , 
        \g[21][50] , \g[21][49] , \g[21][48] , \g[21][47] , \g[21][46] , 
        \g[21][45] , \g[21][44] , \g[21][43] , \g[21][42] , \g[21][41] , 
        \g[21][40] , \g[21][39] , \g[21][38] , \g[21][37] , \g[21][36] , 
        \g[21][35] , \g[21][34] , \g[21][33] , \g[21][32] , \g[21][31] , 
        \g[21][30] , \g[21][29] , \g[21][28] , \g[21][27] , \g[21][26] , 
        \g[21][25] , \g[21][24] , \g[21][23] , \g[21][22] , \g[21][21] , 
        \g[21][20] , \g[21][19] , \g[21][18] , \g[21][17] , \g[21][16] , 
        \g[21][15] , \g[21][14] , \g[21][13] , \g[21][12] , \g[21][11] , 
        \g[21][10] , \g[21][9] , \g[21][8] , \g[21][7] , \g[21][6] , 
        \g[21][5] , \g[21][4] , \g[21][3] , \g[21][2] , \g[21][1] , 
        SYNOPSYS_UNCONNECTED__0}) );
  FullAdder \level1[1].x6  ( .a({n419, n419, n419, n419, n419, n419, n418, 
        n418, n418, n418, n418, n418, n418, n418, n418, n418, n418, n418, n417, 
        n417, n417, n417, n417, n417, n417, n417, n417, n417, n417, n417, 
        \p[3][33] , \p[3][32] , \p[3][31] , \p[3][30] , \p[3][29] , \p[3][28] , 
        \p[3][27] , \p[3][26] , \p[3][25] , \p[3][24] , \p[3][23] , \p[3][22] , 
        \p[3][21] , \p[3][20] , \p[3][19] , \p[3][18] , \p[3][17] , \p[3][16] , 
        \p[3][15] , \p[3][14] , \p[3][13] , \p[3][12] , \p[3][11] , \p[3][10] , 
        \p[3][9] , \p[3][8] , \p[3][7] , \p[3][6] , \p[3][5] , \p[3][4] , 
        \p[3][3] , 1'b0, 1'b0, 1'b0}), .b({n422, n422, n422, n422, n422, n421, 
        n421, n421, n421, n421, n421, n421, n421, n421, n421, n421, n421, n420, 
        n420, n420, n420, n420, n420, n420, n420, n420, n420, n420, n420, 
        \p[4][34] , \p[4][33] , \p[4][32] , \p[4][31] , \p[4][30] , \p[4][29] , 
        \p[4][28] , \p[4][27] , \p[4][26] , \p[4][25] , \p[4][24] , \p[4][23] , 
        \p[4][22] , \p[4][21] , \p[4][20] , \p[4][19] , \p[4][18] , \p[4][17] , 
        \p[4][16] , \p[4][15] , \p[4][14] , \p[4][13] , \p[4][12] , \p[4][11] , 
        \p[4][10] , \p[4][9] , \p[4][8] , \p[4][7] , \p[4][6] , \p[4][5] , 
        \p[4][4] , 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n425, n425, n425, n425, 
        n424, n424, n424, n424, n424, n424, n424, n424, n424, n424, n424, n424, 
        n423, n423, n423, n423, n423, n423, n423, n423, n423, n423, n423, n423, 
        \p[5][35] , \p[5][34] , \p[5][33] , \p[5][32] , \p[5][31] , \p[5][30] , 
        \p[5][29] , \p[5][28] , \p[5][27] , \p[5][26] , \p[5][25] , \p[5][24] , 
        \p[5][23] , \p[5][22] , \p[5][21] , \p[5][20] , \p[5][19] , \p[5][18] , 
        \p[5][17] , \p[5][16] , \p[5][15] , \p[5][14] , \p[5][13] , \p[5][12] , 
        \p[5][11] , \p[5][10] , \p[5][9] , \p[5][8] , \p[5][7] , \p[5][6] , 
        \p[5][5] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[1][63] , 
        \g[1][62] , \g[1][61] , \g[1][60] , \g[1][59] , \g[1][58] , \g[1][57] , 
        \g[1][56] , \g[1][55] , \g[1][54] , \g[1][53] , \g[1][52] , \g[1][51] , 
        \g[1][50] , \g[1][49] , \g[1][48] , \g[1][47] , \g[1][46] , \g[1][45] , 
        \g[1][44] , \g[1][43] , \g[1][42] , \g[1][41] , \g[1][40] , \g[1][39] , 
        \g[1][38] , \g[1][37] , \g[1][36] , \g[1][35] , \g[1][34] , \g[1][33] , 
        \g[1][32] , \g[1][31] , \g[1][30] , \g[1][29] , \g[1][28] , \g[1][27] , 
        \g[1][26] , \g[1][25] , \g[1][24] , \g[1][23] , \g[1][22] , \g[1][21] , 
        \g[1][20] , \g[1][19] , \g[1][18] , \g[1][17] , \g[1][16] , \g[1][15] , 
        \g[1][14] , \g[1][13] , \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , 
        \g[1][8] , \g[1][7] , \g[1][6] , \g[1][5] , \g[1][4] , \g[1][3] , 
        \g[1][2] , \g[1][1] , \g[1][0] }), .cout({\g[22][63] , \g[22][62] , 
        \g[22][61] , \g[22][60] , \g[22][59] , \g[22][58] , \g[22][57] , 
        \g[22][56] , \g[22][55] , \g[22][54] , \g[22][53] , \g[22][52] , 
        \g[22][51] , \g[22][50] , \g[22][49] , \g[22][48] , \g[22][47] , 
        \g[22][46] , \g[22][45] , \g[22][44] , \g[22][43] , \g[22][42] , 
        \g[22][41] , \g[22][40] , \g[22][39] , \g[22][38] , \g[22][37] , 
        \g[22][36] , \g[22][35] , \g[22][34] , \g[22][33] , \g[22][32] , 
        \g[22][31] , \g[22][30] , \g[22][29] , \g[22][28] , \g[22][27] , 
        \g[22][26] , \g[22][25] , \g[22][24] , \g[22][23] , \g[22][22] , 
        \g[22][21] , \g[22][20] , \g[22][19] , \g[22][18] , \g[22][17] , 
        \g[22][16] , \g[22][15] , \g[22][14] , \g[22][13] , \g[22][12] , 
        \g[22][11] , \g[22][10] , \g[22][9] , \g[22][8] , \g[22][7] , 
        \g[22][6] , \g[22][5] , \g[22][4] , \g[22][3] , \g[22][2] , \g[22][1] , 
        SYNOPSYS_UNCONNECTED__1}) );
  FullAdder \level1[2].x6  ( .a({n428, n428, n428, n427, n427, n427, n427, 
        n427, n427, n427, n427, n427, n427, n427, n427, n426, n426, n426, n426, 
        n426, n426, n426, n426, n426, n426, n426, n426, \p[6][36] , \p[6][35] , 
        \p[6][34] , \p[6][33] , \p[6][32] , \p[6][31] , \p[6][30] , \p[6][29] , 
        \p[6][28] , \p[6][27] , \p[6][26] , \p[6][25] , \p[6][24] , \p[6][23] , 
        \p[6][22] , \p[6][21] , \p[6][20] , \p[6][19] , \p[6][18] , \p[6][17] , 
        \p[6][16] , \p[6][15] , \p[6][14] , \p[6][13] , \p[6][12] , \p[6][11] , 
        \p[6][10] , \p[6][9] , \p[6][8] , \p[6][7] , \p[6][6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .b({n431, n431, n430, n430, n430, n430, n430, 
        n430, n430, n430, n430, n430, n430, n430, n429, n429, n429, n429, n429, 
        n429, n429, n429, n429, n429, n429, n429, \p[7][37] , \p[7][36] , 
        \p[7][35] , \p[7][34] , \p[7][33] , \p[7][32] , \p[7][31] , \p[7][30] , 
        \p[7][29] , \p[7][28] , \p[7][27] , \p[7][26] , \p[7][25] , \p[7][24] , 
        \p[7][23] , \p[7][22] , \p[7][21] , \p[7][20] , \p[7][19] , \p[7][18] , 
        \p[7][17] , \p[7][16] , \p[7][15] , \p[7][14] , \p[7][13] , \p[7][12] , 
        \p[7][11] , \p[7][10] , \p[7][9] , \p[7][8] , \p[7][7] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n321, n321, n321, n321, n321, 
        n321, n321, n320, n320, n320, n320, n320, n320, n319, n319, n319, n319, 
        n319, n319, n318, n318, n318, n318, n318, n318, \p[8][38] , \p[8][37] , 
        \p[8][36] , \p[8][35] , \p[8][34] , \p[8][33] , \p[8][32] , \p[8][31] , 
        \p[8][30] , \p[8][29] , \p[8][28] , \p[8][27] , \p[8][26] , \p[8][25] , 
        \p[8][24] , \p[8][23] , \p[8][22] , \p[8][21] , \p[8][20] , \p[8][19] , 
        \p[8][18] , \p[8][17] , \p[8][16] , \p[8][15] , \p[8][14] , \p[8][13] , 
        \p[8][12] , \p[8][11] , \p[8][10] , \p[8][9] , \p[8][8] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[2][63] , \g[2][62] , 
        \g[2][61] , \g[2][60] , \g[2][59] , \g[2][58] , \g[2][57] , \g[2][56] , 
        \g[2][55] , \g[2][54] , \g[2][53] , \g[2][52] , \g[2][51] , \g[2][50] , 
        \g[2][49] , \g[2][48] , \g[2][47] , \g[2][46] , \g[2][45] , \g[2][44] , 
        \g[2][43] , \g[2][42] , \g[2][41] , \g[2][40] , \g[2][39] , \g[2][38] , 
        \g[2][37] , \g[2][36] , \g[2][35] , \g[2][34] , \g[2][33] , \g[2][32] , 
        \g[2][31] , \g[2][30] , \g[2][29] , \g[2][28] , \g[2][27] , \g[2][26] , 
        \g[2][25] , \g[2][24] , \g[2][23] , \g[2][22] , \g[2][21] , \g[2][20] , 
        \g[2][19] , \g[2][18] , \g[2][17] , \g[2][16] , \g[2][15] , \g[2][14] , 
        \g[2][13] , \g[2][12] , \g[2][11] , \g[2][10] , \g[2][9] , \g[2][8] , 
        \g[2][7] , \g[2][6] , \g[2][5] , \g[2][4] , \g[2][3] , \g[2][2] , 
        \g[2][1] , \g[2][0] }), .cout({\g[23][63] , \g[23][62] , \g[23][61] , 
        \g[23][60] , \g[23][59] , \g[23][58] , \g[23][57] , \g[23][56] , 
        \g[23][55] , \g[23][54] , \g[23][53] , \g[23][52] , \g[23][51] , 
        \g[23][50] , \g[23][49] , \g[23][48] , \g[23][47] , \g[23][46] , 
        \g[23][45] , \g[23][44] , \g[23][43] , \g[23][42] , \g[23][41] , 
        \g[23][40] , \g[23][39] , \g[23][38] , \g[23][37] , \g[23][36] , 
        \g[23][35] , \g[23][34] , \g[23][33] , \g[23][32] , \g[23][31] , 
        \g[23][30] , \g[23][29] , \g[23][28] , \g[23][27] , \g[23][26] , 
        \g[23][25] , \g[23][24] , \g[23][23] , \g[23][22] , \g[23][21] , 
        \g[23][20] , \g[23][19] , \g[23][18] , \g[23][17] , \g[23][16] , 
        \g[23][15] , \g[23][14] , \g[23][13] , \g[23][12] , \g[23][11] , 
        \g[23][10] , \g[23][9] , \g[23][8] , \g[23][7] , \g[23][6] , 
        \g[23][5] , \g[23][4] , \g[23][3] , \g[23][2] , \g[23][1] , 
        SYNOPSYS_UNCONNECTED__2}) );
  FullAdder \level1[3].x6  ( .a({n323, n323, n323, n323, n323, n323, n323, 
        n323, n323, n323, n323, n323, n322, n322, n322, n322, n322, n322, n322, 
        n322, n322, n322, n322, n322, \p[9][39] , \p[9][38] , \p[9][37] , 
        \p[9][36] , \p[9][35] , \p[9][34] , \p[9][33] , \p[9][32] , \p[9][31] , 
        \p[9][30] , \p[9][29] , \p[9][28] , \p[9][27] , \p[9][26] , \p[9][25] , 
        \p[9][24] , \p[9][23] , \p[9][22] , \p[9][21] , \p[9][20] , \p[9][19] , 
        \p[9][18] , \p[9][17] , \p[9][16] , \p[9][15] , \p[9][14] , \p[9][13] , 
        \p[9][12] , \p[9][11] , \p[9][10] , \p[9][9] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n325, n325, n325, n325, n325, n325, 
        n325, n325, n325, n325, n325, n324, n324, n324, n324, n324, n324, n324, 
        n324, n324, n324, n324, n324, \p[10][40] , \p[10][39] , \p[10][38] , 
        \p[10][37] , \p[10][36] , \p[10][35] , \p[10][34] , \p[10][33] , 
        \p[10][32] , \p[10][31] , \p[10][30] , \p[10][29] , \p[10][28] , 
        \p[10][27] , \p[10][26] , \p[10][25] , \p[10][24] , \p[10][23] , 
        \p[10][22] , \p[10][21] , \p[10][20] , \p[10][19] , \p[10][18] , 
        \p[10][17] , \p[10][16] , \p[10][15] , \p[10][14] , \p[10][13] , 
        \p[10][12] , \p[10][11] , \p[10][10] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n327, n327, n327, n327, n327, 
        n327, n327, n327, n327, n327, n326, n326, n326, n326, n326, n326, n326, 
        n326, n326, n326, n326, n326, \p[11][41] , \p[11][40] , \p[11][39] , 
        \p[11][38] , \p[11][37] , \p[11][36] , \p[11][35] , \p[11][34] , 
        \p[11][33] , \p[11][32] , \p[11][31] , \p[11][30] , \p[11][29] , 
        \p[11][28] , \p[11][27] , \p[11][26] , \p[11][25] , \p[11][24] , 
        \p[11][23] , \p[11][22] , \p[11][21] , \p[11][20] , \p[11][19] , 
        \p[11][18] , \p[11][17] , \p[11][16] , \p[11][15] , \p[11][14] , 
        \p[11][13] , \p[11][12] , \p[11][11] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[3][63] , \g[3][62] , 
        \g[3][61] , \g[3][60] , \g[3][59] , \g[3][58] , \g[3][57] , \g[3][56] , 
        \g[3][55] , \g[3][54] , \g[3][53] , \g[3][52] , \g[3][51] , \g[3][50] , 
        \g[3][49] , \g[3][48] , \g[3][47] , \g[3][46] , \g[3][45] , \g[3][44] , 
        \g[3][43] , \g[3][42] , \g[3][41] , \g[3][40] , \g[3][39] , \g[3][38] , 
        \g[3][37] , \g[3][36] , \g[3][35] , \g[3][34] , \g[3][33] , \g[3][32] , 
        \g[3][31] , \g[3][30] , \g[3][29] , \g[3][28] , \g[3][27] , \g[3][26] , 
        \g[3][25] , \g[3][24] , \g[3][23] , \g[3][22] , \g[3][21] , \g[3][20] , 
        \g[3][19] , \g[3][18] , \g[3][17] , \g[3][16] , \g[3][15] , \g[3][14] , 
        \g[3][13] , \g[3][12] , \g[3][11] , \g[3][10] , \g[3][9] , \g[3][8] , 
        \g[3][7] , \g[3][6] , \g[3][5] , \g[3][4] , \g[3][3] , \g[3][2] , 
        \g[3][1] , \g[3][0] }), .cout({\g[24][63] , \g[24][62] , \g[24][61] , 
        \g[24][60] , \g[24][59] , \g[24][58] , \g[24][57] , \g[24][56] , 
        \g[24][55] , \g[24][54] , \g[24][53] , \g[24][52] , \g[24][51] , 
        \g[24][50] , \g[24][49] , \g[24][48] , \g[24][47] , \g[24][46] , 
        \g[24][45] , \g[24][44] , \g[24][43] , \g[24][42] , \g[24][41] , 
        \g[24][40] , \g[24][39] , \g[24][38] , \g[24][37] , \g[24][36] , 
        \g[24][35] , \g[24][34] , \g[24][33] , \g[24][32] , \g[24][31] , 
        \g[24][30] , \g[24][29] , \g[24][28] , \g[24][27] , \g[24][26] , 
        \g[24][25] , \g[24][24] , \g[24][23] , \g[24][22] , \g[24][21] , 
        \g[24][20] , \g[24][19] , \g[24][18] , \g[24][17] , \g[24][16] , 
        \g[24][15] , \g[24][14] , \g[24][13] , \g[24][12] , \g[24][11] , 
        \g[24][10] , \g[24][9] , \g[24][8] , \g[24][7] , \g[24][6] , 
        \g[24][5] , \g[24][4] , \g[24][3] , \g[24][2] , \g[24][1] , 
        SYNOPSYS_UNCONNECTED__3}) );
  FullAdder \level1[4].x6  ( .a({n329, n329, n329, n329, n329, n329, n329, 
        n329, n329, n328, n328, n328, n328, n328, n328, n328, n328, n328, n328, 
        n328, n328, \p[12][42] , \p[12][41] , \p[12][40] , \p[12][39] , 
        \p[12][38] , \p[12][37] , \p[12][36] , \p[12][35] , \p[12][34] , 
        \p[12][33] , \p[12][32] , \p[12][31] , \p[12][30] , \p[12][29] , 
        \p[12][28] , \p[12][27] , \p[12][26] , \p[12][25] , \p[12][24] , 
        \p[12][23] , \p[12][22] , \p[12][21] , \p[12][20] , \p[12][19] , 
        \p[12][18] , \p[12][17] , \p[12][16] , \p[12][15] , \p[12][14] , 
        \p[12][13] , \p[12][12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n331, n331, n331, n331, n331, n331, 
        n331, n331, n330, n330, n330, n330, n330, n330, n330, n330, n330, n330, 
        n330, n330, \p[13][43] , \p[13][42] , \p[13][41] , \p[13][40] , 
        \p[13][39] , \p[13][38] , \p[13][37] , \p[13][36] , \p[13][35] , 
        \p[13][34] , \p[13][33] , \p[13][32] , \p[13][31] , \p[13][30] , 
        \p[13][29] , \p[13][28] , \p[13][27] , \p[13][26] , \p[13][25] , 
        \p[13][24] , \p[13][23] , \p[13][22] , \p[13][21] , \p[13][20] , 
        \p[13][19] , \p[13][18] , \p[13][17] , \p[13][16] , \p[13][15] , 
        \p[13][14] , \p[13][13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n333, n333, n333, n333, 
        n333, n333, n333, n332, n332, n332, n332, n332, n332, n332, n332, n332, 
        n332, n332, n332, \p[14][44] , \p[14][43] , \p[14][42] , \p[14][41] , 
        \p[14][40] , \p[14][39] , \p[14][38] , \p[14][37] , \p[14][36] , 
        \p[14][35] , \p[14][34] , \p[14][33] , \p[14][32] , \p[14][31] , 
        \p[14][30] , \p[14][29] , \p[14][28] , \p[14][27] , \p[14][26] , 
        \p[14][25] , \p[14][24] , \p[14][23] , \p[14][22] , \p[14][21] , 
        \p[14][20] , \p[14][19] , \p[14][18] , \p[14][17] , \p[14][16] , 
        \p[14][15] , \p[14][14] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[4][63] , 
        \g[4][62] , \g[4][61] , \g[4][60] , \g[4][59] , \g[4][58] , \g[4][57] , 
        \g[4][56] , \g[4][55] , \g[4][54] , \g[4][53] , \g[4][52] , \g[4][51] , 
        \g[4][50] , \g[4][49] , \g[4][48] , \g[4][47] , \g[4][46] , \g[4][45] , 
        \g[4][44] , \g[4][43] , \g[4][42] , \g[4][41] , \g[4][40] , \g[4][39] , 
        \g[4][38] , \g[4][37] , \g[4][36] , \g[4][35] , \g[4][34] , \g[4][33] , 
        \g[4][32] , \g[4][31] , \g[4][30] , \g[4][29] , \g[4][28] , \g[4][27] , 
        \g[4][26] , \g[4][25] , \g[4][24] , \g[4][23] , \g[4][22] , \g[4][21] , 
        \g[4][20] , \g[4][19] , \g[4][18] , \g[4][17] , \g[4][16] , \g[4][15] , 
        \g[4][14] , \g[4][13] , \g[4][12] , \g[4][11] , \g[4][10] , \g[4][9] , 
        \g[4][8] , \g[4][7] , \g[4][6] , \g[4][5] , \g[4][4] , \g[4][3] , 
        \g[4][2] , \g[4][1] , \g[4][0] }), .cout({\g[25][63] , \g[25][62] , 
        \g[25][61] , \g[25][60] , \g[25][59] , \g[25][58] , \g[25][57] , 
        \g[25][56] , \g[25][55] , \g[25][54] , \g[25][53] , \g[25][52] , 
        \g[25][51] , \g[25][50] , \g[25][49] , \g[25][48] , \g[25][47] , 
        \g[25][46] , \g[25][45] , \g[25][44] , \g[25][43] , \g[25][42] , 
        \g[25][41] , \g[25][40] , \g[25][39] , \g[25][38] , \g[25][37] , 
        \g[25][36] , \g[25][35] , \g[25][34] , \g[25][33] , \g[25][32] , 
        \g[25][31] , \g[25][30] , \g[25][29] , \g[25][28] , \g[25][27] , 
        \g[25][26] , \g[25][25] , \g[25][24] , \g[25][23] , \g[25][22] , 
        \g[25][21] , \g[25][20] , \g[25][19] , \g[25][18] , \g[25][17] , 
        \g[25][16] , \g[25][15] , \g[25][14] , \g[25][13] , \g[25][12] , 
        \g[25][11] , \g[25][10] , \g[25][9] , \g[25][8] , \g[25][7] , 
        \g[25][6] , \g[25][5] , \g[25][4] , \g[25][3] , \g[25][2] , \g[25][1] , 
        SYNOPSYS_UNCONNECTED__4}) );
  FullAdder \level1[5].x6  ( .a({n336, n336, n336, n336, n336, n336, n335, 
        n335, n335, n335, n335, n335, n334, n334, n334, n334, n334, n334, 
        \p[15][45] , \p[15][44] , \p[15][43] , \p[15][42] , \p[15][41] , 
        \p[15][40] , \p[15][39] , \p[15][38] , \p[15][37] , \p[15][36] , 
        \p[15][35] , \p[15][34] , \p[15][33] , \p[15][32] , \p[15][31] , 
        \p[15][30] , \p[15][29] , \p[15][28] , \p[15][27] , \p[15][26] , 
        \p[15][25] , \p[15][24] , \p[15][23] , \p[15][22] , \p[15][21] , 
        \p[15][20] , \p[15][19] , \p[15][18] , \p[15][17] , \p[15][16] , 
        \p[15][15] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n339, n339, n339, n339, n339, 
        n338, n338, n338, n338, n338, n338, n337, n337, n337, n337, n337, n337, 
        \p[16][46] , \p[16][45] , \p[16][44] , \p[16][43] , \p[16][42] , 
        \p[16][41] , \p[16][40] , \p[16][39] , \p[16][38] , \p[16][37] , 
        \p[16][36] , \p[16][35] , \p[16][34] , \p[16][33] , \p[16][32] , 
        \p[16][31] , \p[16][30] , \p[16][29] , \p[16][28] , \p[16][27] , 
        \p[16][26] , \p[16][25] , \p[16][24] , \p[16][23] , \p[16][22] , 
        \p[16][21] , \p[16][20] , \p[16][19] , \p[16][18] , \p[16][17] , 
        \p[16][16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n342, n342, n342, 
        n342, n341, n341, n341, n341, n341, n341, n340, n340, n340, n340, n340, 
        n340, \p[17][47] , \p[17][46] , \p[17][45] , \p[17][44] , \p[17][43] , 
        \p[17][42] , \p[17][41] , \p[17][40] , \p[17][39] , \p[17][38] , 
        \p[17][37] , \p[17][36] , \p[17][35] , \p[17][34] , \p[17][33] , 
        \p[17][32] , \p[17][31] , \p[17][30] , \p[17][29] , \p[17][28] , 
        \p[17][27] , \p[17][26] , \p[17][25] , \p[17][24] , \p[17][23] , 
        \p[17][22] , \p[17][21] , \p[17][20] , \p[17][19] , \p[17][18] , 
        \p[17][17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[5][63] , 
        \g[5][62] , \g[5][61] , \g[5][60] , \g[5][59] , \g[5][58] , \g[5][57] , 
        \g[5][56] , \g[5][55] , \g[5][54] , \g[5][53] , \g[5][52] , \g[5][51] , 
        \g[5][50] , \g[5][49] , \g[5][48] , \g[5][47] , \g[5][46] , \g[5][45] , 
        \g[5][44] , \g[5][43] , \g[5][42] , \g[5][41] , \g[5][40] , \g[5][39] , 
        \g[5][38] , \g[5][37] , \g[5][36] , \g[5][35] , \g[5][34] , \g[5][33] , 
        \g[5][32] , \g[5][31] , \g[5][30] , \g[5][29] , \g[5][28] , \g[5][27] , 
        \g[5][26] , \g[5][25] , \g[5][24] , \g[5][23] , \g[5][22] , \g[5][21] , 
        \g[5][20] , \g[5][19] , \g[5][18] , \g[5][17] , \g[5][16] , \g[5][15] , 
        \g[5][14] , \g[5][13] , \g[5][12] , \g[5][11] , \g[5][10] , \g[5][9] , 
        \g[5][8] , \g[5][7] , \g[5][6] , \g[5][5] , \g[5][4] , \g[5][3] , 
        \g[5][2] , \g[5][1] , \g[5][0] }), .cout({\g[26][63] , \g[26][62] , 
        \g[26][61] , \g[26][60] , \g[26][59] , \g[26][58] , \g[26][57] , 
        \g[26][56] , \g[26][55] , \g[26][54] , \g[26][53] , \g[26][52] , 
        \g[26][51] , \g[26][50] , \g[26][49] , \g[26][48] , \g[26][47] , 
        \g[26][46] , \g[26][45] , \g[26][44] , \g[26][43] , \g[26][42] , 
        \g[26][41] , \g[26][40] , \g[26][39] , \g[26][38] , \g[26][37] , 
        \g[26][36] , \g[26][35] , \g[26][34] , \g[26][33] , \g[26][32] , 
        \g[26][31] , \g[26][30] , \g[26][29] , \g[26][28] , \g[26][27] , 
        \g[26][26] , \g[26][25] , \g[26][24] , \g[26][23] , \g[26][22] , 
        \g[26][21] , \g[26][20] , \g[26][19] , \g[26][18] , \g[26][17] , 
        \g[26][16] , \g[26][15] , \g[26][14] , \g[26][13] , \g[26][12] , 
        \g[26][11] , \g[26][10] , \g[26][9] , \g[26][8] , \g[26][7] , 
        \g[26][6] , \g[26][5] , \g[26][4] , \g[26][3] , \g[26][2] , \g[26][1] , 
        SYNOPSYS_UNCONNECTED__5}) );
  FullAdder \level1[6].x6  ( .a({n345, n345, n345, n344, n344, n344, n344, 
        n344, n344, n343, n343, n343, n343, n343, n343, \p[18][48] , 
        \p[18][47] , \p[18][46] , \p[18][45] , \p[18][44] , \p[18][43] , 
        \p[18][42] , \p[18][41] , \p[18][40] , \p[18][39] , \p[18][38] , 
        \p[18][37] , \p[18][36] , \p[18][35] , \p[18][34] , \p[18][33] , 
        \p[18][32] , \p[18][31] , \p[18][30] , \p[18][29] , \p[18][28] , 
        \p[18][27] , \p[18][26] , \p[18][25] , \p[18][24] , \p[18][23] , 
        \p[18][22] , \p[18][21] , \p[18][20] , \p[18][19] , \p[18][18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n348, n348, n347, n347, n347, n347, 
        n347, n347, n346, n346, n346, n346, n346, n346, \p[19][49] , 
        \p[19][48] , \p[19][47] , \p[19][46] , \p[19][45] , \p[19][44] , 
        \p[19][43] , \p[19][42] , \p[19][41] , \p[19][40] , \p[19][39] , 
        \p[19][38] , \p[19][37] , \p[19][36] , \p[19][35] , \p[19][34] , 
        \p[19][33] , \p[19][32] , \p[19][31] , \p[19][30] , \p[19][29] , 
        \p[19][28] , \p[19][27] , \p[19][26] , \p[19][25] , \p[19][24] , 
        \p[19][23] , \p[19][22] , \p[19][21] , \p[19][20] , \p[19][19] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n350, n350, n350, n350, 
        n350, n350, n350, n349, n349, n349, n349, n349, n349, \p[20][50] , 
        \p[20][49] , \p[20][48] , \p[20][47] , \p[20][46] , \p[20][45] , 
        \p[20][44] , \p[20][43] , \p[20][42] , \p[20][41] , \p[20][40] , 
        \p[20][39] , \p[20][38] , \p[20][37] , \p[20][36] , \p[20][35] , 
        \p[20][34] , \p[20][33] , \p[20][32] , \p[20][31] , \p[20][30] , 
        \p[20][29] , \p[20][28] , \p[20][27] , \p[20][26] , \p[20][25] , 
        \p[20][24] , \p[20][23] , \p[20][22] , \p[20][21] , \p[20][20] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[6][63] , 
        \g[6][62] , \g[6][61] , \g[6][60] , \g[6][59] , \g[6][58] , \g[6][57] , 
        \g[6][56] , \g[6][55] , \g[6][54] , \g[6][53] , \g[6][52] , \g[6][51] , 
        \g[6][50] , \g[6][49] , \g[6][48] , \g[6][47] , \g[6][46] , \g[6][45] , 
        \g[6][44] , \g[6][43] , \g[6][42] , \g[6][41] , \g[6][40] , \g[6][39] , 
        \g[6][38] , \g[6][37] , \g[6][36] , \g[6][35] , \g[6][34] , \g[6][33] , 
        \g[6][32] , \g[6][31] , \g[6][30] , \g[6][29] , \g[6][28] , \g[6][27] , 
        \g[6][26] , \g[6][25] , \g[6][24] , \g[6][23] , \g[6][22] , \g[6][21] , 
        \g[6][20] , \g[6][19] , \g[6][18] , \g[6][17] , \g[6][16] , \g[6][15] , 
        \g[6][14] , \g[6][13] , \g[6][12] , \g[6][11] , \g[6][10] , \g[6][9] , 
        \g[6][8] , \g[6][7] , \g[6][6] , \g[6][5] , \g[6][4] , \g[6][3] , 
        \g[6][2] , \g[6][1] , \g[6][0] }), .cout({\g[27][63] , \g[27][62] , 
        \g[27][61] , \g[27][60] , \g[27][59] , \g[27][58] , \g[27][57] , 
        \g[27][56] , \g[27][55] , \g[27][54] , \g[27][53] , \g[27][52] , 
        \g[27][51] , \g[27][50] , \g[27][49] , \g[27][48] , \g[27][47] , 
        \g[27][46] , \g[27][45] , \g[27][44] , \g[27][43] , \g[27][42] , 
        \g[27][41] , \g[27][40] , \g[27][39] , \g[27][38] , \g[27][37] , 
        \g[27][36] , \g[27][35] , \g[27][34] , \g[27][33] , \g[27][32] , 
        \g[27][31] , \g[27][30] , \g[27][29] , \g[27][28] , \g[27][27] , 
        \g[27][26] , \g[27][25] , \g[27][24] , \g[27][23] , \g[27][22] , 
        \g[27][21] , \g[27][20] , \g[27][19] , \g[27][18] , \g[27][17] , 
        \g[27][16] , \g[27][15] , \g[27][14] , \g[27][13] , \g[27][12] , 
        \g[27][11] , \g[27][10] , \g[27][9] , \g[27][8] , \g[27][7] , 
        \g[27][6] , \g[27][5] , \g[27][4] , \g[27][3] , \g[27][2] , \g[27][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  FullAdder \level1[7].x6  ( .a({\p[21][63] , \p[21][63] , \p[21][63] , 
        \p[21][63] , \p[21][63] , \p[21][63] , \p[21][63] , \p[21][63] , 
        \p[21][63] , \p[21][63] , \p[21][63] , \p[21][63] , \p[21][51] , 
        \p[21][50] , \p[21][49] , \p[21][48] , \p[21][47] , \p[21][46] , 
        \p[21][45] , \p[21][44] , \p[21][43] , \p[21][42] , \p[21][41] , 
        \p[21][40] , \p[21][39] , \p[21][38] , \p[21][37] , \p[21][36] , 
        \p[21][35] , \p[21][34] , \p[21][33] , \p[21][32] , \p[21][31] , 
        \p[21][30] , \p[21][29] , \p[21][28] , \p[21][27] , \p[21][26] , 
        \p[21][25] , \p[21][24] , \p[21][23] , \p[21][22] , \p[21][21] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({\p[22][63] , 
        \p[22][63] , \p[22][63] , \p[22][63] , \p[22][63] , \p[22][63] , 
        \p[22][63] , \p[22][63] , \p[22][63] , \p[22][63] , \p[22][63] , 
        \p[22][52] , \p[22][51] , \p[22][50] , \p[22][49] , \p[22][48] , 
        \p[22][47] , \p[22][46] , \p[22][45] , \p[22][44] , \p[22][43] , 
        \p[22][42] , \p[22][41] , \p[22][40] , \p[22][39] , \p[22][38] , 
        \p[22][37] , \p[22][36] , \p[22][35] , \p[22][34] , \p[22][33] , 
        \p[22][32] , \p[22][31] , \p[22][30] , \p[22][29] , \p[22][28] , 
        \p[22][27] , \p[22][26] , \p[22][25] , \p[22][24] , \p[22][23] , 
        \p[22][22] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .cin({\p[23][63] , \p[23][63] , \p[23][63] , \p[23][63] , 
        \p[23][63] , \p[23][63] , \p[23][63] , \p[23][63] , \p[23][63] , 
        \p[23][63] , \p[23][53] , \p[23][52] , \p[23][51] , \p[23][50] , 
        \p[23][49] , \p[23][48] , \p[23][47] , \p[23][46] , \p[23][45] , 
        \p[23][44] , \p[23][43] , \p[23][42] , \p[23][41] , \p[23][40] , 
        \p[23][39] , \p[23][38] , \p[23][37] , \p[23][36] , \p[23][35] , 
        \p[23][34] , \p[23][33] , \p[23][32] , \p[23][31] , \p[23][30] , 
        \p[23][29] , \p[23][28] , \p[23][27] , \p[23][26] , \p[23][25] , 
        \p[23][24] , \p[23][23] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[7][63] , \g[7][62] , \g[7][61] , 
        \g[7][60] , \g[7][59] , \g[7][58] , \g[7][57] , \g[7][56] , \g[7][55] , 
        \g[7][54] , \g[7][53] , \g[7][52] , \g[7][51] , \g[7][50] , \g[7][49] , 
        \g[7][48] , \g[7][47] , \g[7][46] , \g[7][45] , \g[7][44] , \g[7][43] , 
        \g[7][42] , \g[7][41] , \g[7][40] , \g[7][39] , \g[7][38] , \g[7][37] , 
        \g[7][36] , \g[7][35] , \g[7][34] , \g[7][33] , \g[7][32] , \g[7][31] , 
        \g[7][30] , \g[7][29] , \g[7][28] , \g[7][27] , \g[7][26] , \g[7][25] , 
        \g[7][24] , \g[7][23] , \g[7][22] , \g[7][21] , \g[7][20] , \g[7][19] , 
        \g[7][18] , \g[7][17] , \g[7][16] , \g[7][15] , \g[7][14] , \g[7][13] , 
        \g[7][12] , \g[7][11] , \g[7][10] , \g[7][9] , \g[7][8] , \g[7][7] , 
        \g[7][6] , \g[7][5] , \g[7][4] , \g[7][3] , \g[7][2] , \g[7][1] , 
        \g[7][0] }), .cout({\g[28][63] , \g[28][62] , \g[28][61] , \g[28][60] , 
        \g[28][59] , \g[28][58] , \g[28][57] , \g[28][56] , \g[28][55] , 
        \g[28][54] , \g[28][53] , \g[28][52] , \g[28][51] , \g[28][50] , 
        \g[28][49] , \g[28][48] , \g[28][47] , \g[28][46] , \g[28][45] , 
        \g[28][44] , \g[28][43] , \g[28][42] , \g[28][41] , \g[28][40] , 
        \g[28][39] , \g[28][38] , \g[28][37] , \g[28][36] , \g[28][35] , 
        \g[28][34] , \g[28][33] , \g[28][32] , \g[28][31] , \g[28][30] , 
        \g[28][29] , \g[28][28] , \g[28][27] , \g[28][26] , \g[28][25] , 
        \g[28][24] , \g[28][23] , \g[28][22] , \g[28][21] , \g[28][20] , 
        \g[28][19] , \g[28][18] , \g[28][17] , \g[28][16] , \g[28][15] , 
        \g[28][14] , \g[28][13] , \g[28][12] , \g[28][11] , \g[28][10] , 
        \g[28][9] , \g[28][8] , \g[28][7] , \g[28][6] , \g[28][5] , \g[28][4] , 
        \g[28][3] , \g[28][2] , \g[28][1] , SYNOPSYS_UNCONNECTED__7}) );
  FullAdder \level1[8].x6  ( .a({\p[24][63] , \p[24][63] , \p[24][63] , 
        \p[24][63] , \p[24][63] , \p[24][63] , \p[24][63] , \p[24][63] , 
        \p[24][63] , \p[24][54] , \p[24][53] , \p[24][52] , \p[24][51] , 
        \p[24][50] , \p[24][49] , \p[24][48] , \p[24][47] , \p[24][46] , 
        \p[24][45] , \p[24][44] , \p[24][43] , \p[24][42] , \p[24][41] , 
        \p[24][40] , \p[24][39] , \p[24][38] , \p[24][37] , \p[24][36] , 
        \p[24][35] , \p[24][34] , \p[24][33] , \p[24][32] , \p[24][31] , 
        \p[24][30] , \p[24][29] , \p[24][28] , \p[24][27] , \p[24][26] , 
        \p[24][25] , \p[24][24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({\p[25][63] , \p[25][63] , 
        \p[25][63] , \p[25][63] , \p[25][63] , \p[25][63] , \p[25][63] , 
        \p[25][63] , \p[25][55] , \p[25][54] , \p[25][53] , \p[25][52] , 
        \p[25][51] , \p[25][50] , \p[25][49] , \p[25][48] , \p[25][47] , 
        \p[25][46] , \p[25][45] , \p[25][44] , \p[25][43] , \p[25][42] , 
        \p[25][41] , \p[25][40] , \p[25][39] , \p[25][38] , \p[25][37] , 
        \p[25][36] , \p[25][35] , \p[25][34] , \p[25][33] , \p[25][32] , 
        \p[25][31] , \p[25][30] , \p[25][29] , \p[25][28] , \p[25][27] , 
        \p[25][26] , \p[25][25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[26][63] , \p[26][63] , 
        \p[26][63] , \p[26][63] , \p[26][63] , \p[26][63] , \p[26][63] , 
        \p[26][56] , \p[26][55] , \p[26][54] , \p[26][53] , \p[26][52] , 
        \p[26][51] , \p[26][50] , \p[26][49] , \p[26][48] , \p[26][47] , 
        \p[26][46] , \p[26][45] , \p[26][44] , \p[26][43] , \p[26][42] , 
        \p[26][41] , \p[26][40] , \p[26][39] , \p[26][38] , \p[26][37] , 
        \p[26][36] , \p[26][35] , \p[26][34] , \p[26][33] , \p[26][32] , 
        \p[26][31] , \p[26][30] , \p[26][29] , \p[26][28] , \p[26][27] , 
        \p[26][26] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[8][63] , \g[8][62] , 
        \g[8][61] , \g[8][60] , \g[8][59] , \g[8][58] , \g[8][57] , \g[8][56] , 
        \g[8][55] , \g[8][54] , \g[8][53] , \g[8][52] , \g[8][51] , \g[8][50] , 
        \g[8][49] , \g[8][48] , \g[8][47] , \g[8][46] , \g[8][45] , \g[8][44] , 
        \g[8][43] , \g[8][42] , \g[8][41] , \g[8][40] , \g[8][39] , \g[8][38] , 
        \g[8][37] , \g[8][36] , \g[8][35] , \g[8][34] , \g[8][33] , \g[8][32] , 
        \g[8][31] , \g[8][30] , \g[8][29] , \g[8][28] , \g[8][27] , \g[8][26] , 
        \g[8][25] , \g[8][24] , \g[8][23] , \g[8][22] , \g[8][21] , \g[8][20] , 
        \g[8][19] , \g[8][18] , \g[8][17] , \g[8][16] , \g[8][15] , \g[8][14] , 
        \g[8][13] , \g[8][12] , \g[8][11] , \g[8][10] , \g[8][9] , \g[8][8] , 
        \g[8][7] , \g[8][6] , \g[8][5] , \g[8][4] , \g[8][3] , \g[8][2] , 
        \g[8][1] , \g[8][0] }), .cout({\g[29][63] , \g[29][62] , \g[29][61] , 
        \g[29][60] , \g[29][59] , \g[29][58] , \g[29][57] , \g[29][56] , 
        \g[29][55] , \g[29][54] , \g[29][53] , \g[29][52] , \g[29][51] , 
        \g[29][50] , \g[29][49] , \g[29][48] , \g[29][47] , \g[29][46] , 
        \g[29][45] , \g[29][44] , \g[29][43] , \g[29][42] , \g[29][41] , 
        \g[29][40] , \g[29][39] , \g[29][38] , \g[29][37] , \g[29][36] , 
        \g[29][35] , \g[29][34] , \g[29][33] , \g[29][32] , \g[29][31] , 
        \g[29][30] , \g[29][29] , \g[29][28] , \g[29][27] , \g[29][26] , 
        \g[29][25] , \g[29][24] , \g[29][23] , \g[29][22] , \g[29][21] , 
        \g[29][20] , \g[29][19] , \g[29][18] , \g[29][17] , \g[29][16] , 
        \g[29][15] , \g[29][14] , \g[29][13] , \g[29][12] , \g[29][11] , 
        \g[29][10] , \g[29][9] , \g[29][8] , \g[29][7] , \g[29][6] , 
        \g[29][5] , \g[29][4] , \g[29][3] , \g[29][2] , \g[29][1] , 
        SYNOPSYS_UNCONNECTED__8}) );
  FullAdder \level1[9].x6  ( .a({\p[27][63] , \p[27][63] , \p[27][63] , 
        \p[27][63] , \p[27][63] , \p[27][63] , \p[27][57] , \p[27][56] , 
        \p[27][55] , \p[27][54] , \p[27][53] , \p[27][52] , \p[27][51] , 
        \p[27][50] , \p[27][49] , \p[27][48] , \p[27][47] , \p[27][46] , 
        \p[27][45] , \p[27][44] , \p[27][43] , \p[27][42] , \p[27][41] , 
        \p[27][40] , \p[27][39] , \p[27][38] , \p[27][37] , \p[27][36] , 
        \p[27][35] , \p[27][34] , \p[27][33] , \p[27][32] , \p[27][31] , 
        \p[27][30] , \p[27][29] , \p[27][28] , \p[27][27] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({\p[28][63] , \p[28][63] , \p[28][63] , \p[28][63] , \p[28][63] , 
        \p[28][58] , \p[28][57] , \p[28][56] , \p[28][55] , \p[28][54] , 
        \p[28][53] , \p[28][52] , \p[28][51] , \p[28][50] , \p[28][49] , 
        \p[28][48] , \p[28][47] , \p[28][46] , \p[28][45] , \p[28][44] , 
        \p[28][43] , \p[28][42] , \p[28][41] , \p[28][40] , \p[28][39] , 
        \p[28][38] , \p[28][37] , \p[28][36] , \p[28][35] , \p[28][34] , 
        \p[28][33] , \p[28][32] , \p[28][31] , \p[28][30] , \p[28][29] , 
        \p[28][28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[29][63] , 
        \p[29][63] , \p[29][63] , \p[29][63] , \p[29][59] , \p[29][58] , 
        \p[29][57] , \p[29][56] , \p[29][55] , \p[29][54] , \p[29][53] , 
        \p[29][52] , \p[29][51] , \p[29][50] , \p[29][49] , \p[29][48] , 
        \p[29][47] , \p[29][46] , \p[29][45] , \p[29][44] , \p[29][43] , 
        \p[29][42] , \p[29][41] , \p[29][40] , \p[29][39] , \p[29][38] , 
        \p[29][37] , \p[29][36] , \p[29][35] , \p[29][34] , \p[29][33] , 
        \p[29][32] , \p[29][31] , \p[29][30] , \p[29][29] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .sum({\g[9][63] , \g[9][62] , \g[9][61] , \g[9][60] , 
        \g[9][59] , \g[9][58] , \g[9][57] , \g[9][56] , \g[9][55] , \g[9][54] , 
        \g[9][53] , \g[9][52] , \g[9][51] , \g[9][50] , \g[9][49] , \g[9][48] , 
        \g[9][47] , \g[9][46] , \g[9][45] , \g[9][44] , \g[9][43] , \g[9][42] , 
        \g[9][41] , \g[9][40] , \g[9][39] , \g[9][38] , \g[9][37] , \g[9][36] , 
        \g[9][35] , \g[9][34] , \g[9][33] , \g[9][32] , \g[9][31] , \g[9][30] , 
        \g[9][29] , \g[9][28] , \g[9][27] , \g[9][26] , \g[9][25] , \g[9][24] , 
        \g[9][23] , \g[9][22] , \g[9][21] , \g[9][20] , \g[9][19] , \g[9][18] , 
        \g[9][17] , \g[9][16] , \g[9][15] , \g[9][14] , \g[9][13] , \g[9][12] , 
        \g[9][11] , \g[9][10] , \g[9][9] , \g[9][8] , \g[9][7] , \g[9][6] , 
        \g[9][5] , \g[9][4] , \g[9][3] , \g[9][2] , \g[9][1] , \g[9][0] }), 
        .cout({\g[30][63] , \g[30][62] , \g[30][61] , \g[30][60] , \g[30][59] , 
        \g[30][58] , \g[30][57] , \g[30][56] , \g[30][55] , \g[30][54] , 
        \g[30][53] , \g[30][52] , \g[30][51] , \g[30][50] , \g[30][49] , 
        \g[30][48] , \g[30][47] , \g[30][46] , \g[30][45] , \g[30][44] , 
        \g[30][43] , \g[30][42] , \g[30][41] , \g[30][40] , \g[30][39] , 
        \g[30][38] , \g[30][37] , \g[30][36] , \g[30][35] , \g[30][34] , 
        \g[30][33] , \g[30][32] , \g[30][31] , \g[30][30] , \g[30][29] , 
        \g[30][28] , \g[30][27] , \g[30][26] , \g[30][25] , \g[30][24] , 
        \g[30][23] , \g[30][22] , \g[30][21] , \g[30][20] , \g[30][19] , 
        \g[30][18] , \g[30][17] , \g[30][16] , \g[30][15] , \g[30][14] , 
        \g[30][13] , \g[30][12] , \g[30][11] , \g[30][10] , \g[30][9] , 
        \g[30][8] , \g[30][7] , \g[30][6] , \g[30][5] , \g[30][4] , \g[30][3] , 
        \g[30][2] , \g[30][1] , SYNOPSYS_UNCONNECTED__9}) );
  FullAdder \level1[10].x6  ( .a({\p[30][63] , \p[30][63] , \p[30][63] , 
        \p[30][60] , \p[30][59] , \p[30][58] , \p[30][57] , \p[30][56] , 
        \p[30][55] , \p[30][54] , \p[30][53] , \p[30][52] , \p[30][51] , 
        \p[30][50] , \p[30][49] , \p[30][48] , \p[30][47] , \p[30][46] , 
        \p[30][45] , \p[30][44] , \p[30][43] , \p[30][42] , \p[30][41] , 
        \p[30][40] , \p[30][39] , \p[30][38] , \p[30][37] , \p[30][36] , 
        \p[30][35] , \p[30][34] , \p[30][33] , \p[30][32] , \p[30][31] , 
        \p[30][30] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({
        \p[32][63] , \p[32][63] , \p[33][63] , \p[34][63] , \p[35][63] , 
        \p[36][63] , \p[37][63] , \p[38][63] , \p[39][63] , \p[40][63] , 
        \p[41][63] , \p[42][63] , n352, n354, n358, n361, n364, n367, n369, 
        n371, n373, n375, n377, n379, n382, n385, n389, n391, n395, n398, n400, 
        n404, n407, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({
        \p[32][63] , \p[33][63] , \p[34][63] , \p[35][63] , \p[36][63] , 
        \p[37][63] , \p[38][63] , \p[39][63] , \p[40][63] , \p[41][63] , 
        \p[42][63] , n351, n353, n356, n359, n362, n365, n368, n370, n372, 
        n374, n376, n378, n380, n384, n387, n390, n393, n396, n399, n402, n405, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[10][63] , 
        \g[10][62] , \g[10][61] , \g[10][60] , \g[10][59] , \g[10][58] , 
        \g[10][57] , \g[10][56] , \g[10][55] , \g[10][54] , \g[10][53] , 
        \g[10][52] , \g[10][51] , \g[10][50] , \g[10][49] , \g[10][48] , 
        \g[10][47] , \g[10][46] , \g[10][45] , \g[10][44] , \g[10][43] , 
        \g[10][42] , \g[10][41] , \g[10][40] , \g[10][39] , \g[10][38] , 
        \g[10][37] , \g[10][36] , \g[10][35] , \g[10][34] , \g[10][33] , 
        \g[10][32] , \g[10][31] , \g[10][30] , \g[10][29] , \g[10][28] , 
        \g[10][27] , \g[10][26] , \g[10][25] , \g[10][24] , \g[10][23] , 
        \g[10][22] , \g[10][21] , \g[10][20] , \g[10][19] , \g[10][18] , 
        \g[10][17] , \g[10][16] , \g[10][15] , \g[10][14] , \g[10][13] , 
        \g[10][12] , \g[10][11] , \g[10][10] , \g[10][9] , \g[10][8] , 
        \g[10][7] , \g[10][6] , \g[10][5] , \g[10][4] , \g[10][3] , \g[10][2] , 
        \g[10][1] , \g[10][0] }), .cout({\g[31][63] , \g[31][62] , \g[31][61] , 
        \g[31][60] , \g[31][59] , \g[31][58] , \g[31][57] , \g[31][56] , 
        \g[31][55] , \g[31][54] , \g[31][53] , \g[31][52] , \g[31][51] , 
        \g[31][50] , \g[31][49] , \g[31][48] , \g[31][47] , \g[31][46] , 
        \g[31][45] , \g[31][44] , \g[31][43] , \g[31][42] , \g[31][41] , 
        \g[31][40] , \g[31][39] , \g[31][38] , \g[31][37] , \g[31][36] , 
        \g[31][35] , \g[31][34] , \g[31][33] , \g[31][32] , \g[31][31] , 
        \g[31][30] , \g[31][29] , \g[31][28] , \g[31][27] , \g[31][26] , 
        \g[31][25] , \g[31][24] , \g[31][23] , \g[31][22] , \g[31][21] , 
        \g[31][20] , \g[31][19] , \g[31][18] , \g[31][17] , \g[31][16] , 
        \g[31][15] , \g[31][14] , \g[31][13] , \g[31][12] , \g[31][11] , 
        \g[31][10] , \g[31][9] , \g[31][8] , \g[31][7] , \g[31][6] , 
        \g[31][5] , \g[31][4] , \g[31][3] , \g[31][2] , \g[31][1] , 
        SYNOPSYS_UNCONNECTED__10}) );
  FullAdder \level1[11].x6  ( .a({\p[33][63] , \p[34][63] , \p[35][63] , 
        \p[36][63] , \p[37][63] , \p[38][63] , \p[39][63] , \p[40][63] , 
        \p[41][63] , \p[42][63] , n351, n353, n356, n360, n363, n366, n368, 
        n370, n373, n375, n377, n378, n381, n384, n388, n390, n394, n397, n399, 
        n403, n406, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b({\p[34][63] , \p[35][63] , \p[36][63] , \p[37][63] , \p[38][63] , 
        \p[39][63] , \p[40][63] , \p[41][63] , \p[42][63] , n352, n354, n358, 
        n361, n364, n367, n369, n371, n373, n375, n377, n379, n383, n385, n389, 
        n392, n395, n398, n401, n404, n407, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[35][63] , \p[36][63] , \p[37][63] , 
        \p[38][63] , \p[39][63] , \p[40][63] , \p[41][63] , \p[42][63] , n351, 
        n353, n356, n359, n362, n365, n368, n370, n372, n374, n376, n378, n380, 
        n384, n387, n390, n393, n396, n399, n402, n405, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[11][63] , 
        \g[11][62] , \g[11][61] , \g[11][60] , \g[11][59] , \g[11][58] , 
        \g[11][57] , \g[11][56] , \g[11][55] , \g[11][54] , \g[11][53] , 
        \g[11][52] , \g[11][51] , \g[11][50] , \g[11][49] , \g[11][48] , 
        \g[11][47] , \g[11][46] , \g[11][45] , \g[11][44] , \g[11][43] , 
        \g[11][42] , \g[11][41] , \g[11][40] , \g[11][39] , \g[11][38] , 
        \g[11][37] , \g[11][36] , \g[11][35] , \g[11][34] , \g[11][33] , 
        \g[11][32] , \g[11][31] , \g[11][30] , \g[11][29] , \g[11][28] , 
        \g[11][27] , \g[11][26] , \g[11][25] , \g[11][24] , \g[11][23] , 
        \g[11][22] , \g[11][21] , \g[11][20] , \g[11][19] , \g[11][18] , 
        \g[11][17] , \g[11][16] , \g[11][15] , \g[11][14] , \g[11][13] , 
        \g[11][12] , \g[11][11] , \g[11][10] , \g[11][9] , \g[11][8] , 
        \g[11][7] , \g[11][6] , \g[11][5] , \g[11][4] , \g[11][3] , \g[11][2] , 
        \g[11][1] , \g[11][0] }), .cout({\g[32][63] , \g[32][62] , \g[32][61] , 
        \g[32][60] , \g[32][59] , \g[32][58] , \g[32][57] , \g[32][56] , 
        \g[32][55] , \g[32][54] , \g[32][53] , \g[32][52] , \g[32][51] , 
        \g[32][50] , \g[32][49] , \g[32][48] , \g[32][47] , \g[32][46] , 
        \g[32][45] , \g[32][44] , \g[32][43] , \g[32][42] , \g[32][41] , 
        \g[32][40] , \g[32][39] , \g[32][38] , \g[32][37] , \g[32][36] , 
        \g[32][35] , \g[32][34] , \g[32][33] , \g[32][32] , \g[32][31] , 
        \g[32][30] , \g[32][29] , \g[32][28] , \g[32][27] , \g[32][26] , 
        \g[32][25] , \g[32][24] , \g[32][23] , \g[32][22] , \g[32][21] , 
        \g[32][20] , \g[32][19] , \g[32][18] , \g[32][17] , \g[32][16] , 
        \g[32][15] , \g[32][14] , \g[32][13] , \g[32][12] , \g[32][11] , 
        \g[32][10] , \g[32][9] , \g[32][8] , \g[32][7] , \g[32][6] , 
        \g[32][5] , \g[32][4] , \g[32][3] , \g[32][2] , \g[32][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  FullAdder \level1[12].x6  ( .a({\p[36][63] , \p[37][63] , \p[38][63] , 
        \p[39][63] , \p[40][63] , \p[41][63] , \p[42][63] , n352, n354, n357, 
        n359, n363, n366, n368, n370, n372, n375, n377, n378, n381, n384, n388, 
        n390, n394, n396, n400, n403, n406, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({\p[37][63] , \p[38][63] , 
        \p[39][63] , \p[40][63] , \p[41][63] , \p[42][63] , n352, n354, n357, 
        n360, n363, n367, n369, n371, n373, n375, n377, n379, n383, n385, n388, 
        n392, n394, n397, n401, n404, n407, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[38][63] , 
        \p[39][63] , \p[40][63] , \p[41][63] , \p[42][63] , n351, n353, n356, 
        n359, n362, n365, n368, n370, n372, n374, n376, n378, n380, n384, n387, 
        n390, n393, n396, n399, n402, n405, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[12][63] , 
        \g[12][62] , \g[12][61] , \g[12][60] , \g[12][59] , \g[12][58] , 
        \g[12][57] , \g[12][56] , \g[12][55] , \g[12][54] , \g[12][53] , 
        \g[12][52] , \g[12][51] , \g[12][50] , \g[12][49] , \g[12][48] , 
        \g[12][47] , \g[12][46] , \g[12][45] , \g[12][44] , \g[12][43] , 
        \g[12][42] , \g[12][41] , \g[12][40] , \g[12][39] , \g[12][38] , 
        \g[12][37] , \g[12][36] , \g[12][35] , \g[12][34] , \g[12][33] , 
        \g[12][32] , \g[12][31] , \g[12][30] , \g[12][29] , \g[12][28] , 
        \g[12][27] , \g[12][26] , \g[12][25] , \g[12][24] , \g[12][23] , 
        \g[12][22] , \g[12][21] , \g[12][20] , \g[12][19] , \g[12][18] , 
        \g[12][17] , \g[12][16] , \g[12][15] , \g[12][14] , \g[12][13] , 
        \g[12][12] , \g[12][11] , \g[12][10] , \g[12][9] , \g[12][8] , 
        \g[12][7] , \g[12][6] , \g[12][5] , \g[12][4] , \g[12][3] , \g[12][2] , 
        \g[12][1] , \g[12][0] }), .cout({\g[33][63] , \g[33][62] , \g[33][61] , 
        \g[33][60] , \g[33][59] , \g[33][58] , \g[33][57] , \g[33][56] , 
        \g[33][55] , \g[33][54] , \g[33][53] , \g[33][52] , \g[33][51] , 
        \g[33][50] , \g[33][49] , \g[33][48] , \g[33][47] , \g[33][46] , 
        \g[33][45] , \g[33][44] , \g[33][43] , \g[33][42] , \g[33][41] , 
        \g[33][40] , \g[33][39] , \g[33][38] , \g[33][37] , \g[33][36] , 
        \g[33][35] , \g[33][34] , \g[33][33] , \g[33][32] , \g[33][31] , 
        \g[33][30] , \g[33][29] , \g[33][28] , \g[33][27] , \g[33][26] , 
        \g[33][25] , \g[33][24] , \g[33][23] , \g[33][22] , \g[33][21] , 
        \g[33][20] , \g[33][19] , \g[33][18] , \g[33][17] , \g[33][16] , 
        \g[33][15] , \g[33][14] , \g[33][13] , \g[33][12] , \g[33][11] , 
        \g[33][10] , \g[33][9] , \g[33][8] , \g[33][7] , \g[33][6] , 
        \g[33][5] , \g[33][4] , \g[33][3] , \g[33][2] , \g[33][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  FullAdder \level1[13].x6  ( .a({\p[39][63] , \p[40][63] , \p[41][63] , 
        \p[42][63] , n352, n354, n357, n360, n363, n366, n368, n370, n372, 
        n374, n376, n378, n382, n385, n388, n390, n394, n396, n400, n403, n406, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .b({\p[40][63] , \p[41][63] , \p[42][63] , n352, 
        n354, n357, n360, n363, n366, n369, n371, n373, n375, n377, n379, n383, 
        n386, n388, n392, n394, n397, n401, n404, n407, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[41][63] , \p[42][63] , n351, n353, n356, n359, n362, n365, n368, 
        n370, n372, n374, n376, n378, n380, n384, n387, n390, n393, n396, n399, 
        n402, n405, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[13][63] , 
        \g[13][62] , \g[13][61] , \g[13][60] , \g[13][59] , \g[13][58] , 
        \g[13][57] , \g[13][56] , \g[13][55] , \g[13][54] , \g[13][53] , 
        \g[13][52] , \g[13][51] , \g[13][50] , \g[13][49] , \g[13][48] , 
        \g[13][47] , \g[13][46] , \g[13][45] , \g[13][44] , \g[13][43] , 
        \g[13][42] , \g[13][41] , \g[13][40] , \g[13][39] , \g[13][38] , 
        \g[13][37] , \g[13][36] , \g[13][35] , \g[13][34] , \g[13][33] , 
        \g[13][32] , \g[13][31] , \g[13][30] , \g[13][29] , \g[13][28] , 
        \g[13][27] , \g[13][26] , \g[13][25] , \g[13][24] , \g[13][23] , 
        \g[13][22] , \g[13][21] , \g[13][20] , \g[13][19] , \g[13][18] , 
        \g[13][17] , \g[13][16] , \g[13][15] , \g[13][14] , \g[13][13] , 
        \g[13][12] , \g[13][11] , \g[13][10] , \g[13][9] , \g[13][8] , 
        \g[13][7] , \g[13][6] , \g[13][5] , \g[13][4] , \g[13][3] , \g[13][2] , 
        \g[13][1] , \g[13][0] }), .cout({\g[34][63] , \g[34][62] , \g[34][61] , 
        \g[34][60] , \g[34][59] , \g[34][58] , \g[34][57] , \g[34][56] , 
        \g[34][55] , \g[34][54] , \g[34][53] , \g[34][52] , \g[34][51] , 
        \g[34][50] , \g[34][49] , \g[34][48] , \g[34][47] , \g[34][46] , 
        \g[34][45] , \g[34][44] , \g[34][43] , \g[34][42] , \g[34][41] , 
        \g[34][40] , \g[34][39] , \g[34][38] , \g[34][37] , \g[34][36] , 
        \g[34][35] , \g[34][34] , \g[34][33] , \g[34][32] , \g[34][31] , 
        \g[34][30] , \g[34][29] , \g[34][28] , \g[34][27] , \g[34][26] , 
        \g[34][25] , \g[34][24] , \g[34][23] , \g[34][22] , \g[34][21] , 
        \g[34][20] , \g[34][19] , \g[34][18] , \g[34][17] , \g[34][16] , 
        \g[34][15] , \g[34][14] , \g[34][13] , \g[34][12] , \g[34][11] , 
        \g[34][10] , \g[34][9] , \g[34][8] , \g[34][7] , \g[34][6] , 
        \g[34][5] , \g[34][4] , \g[34][3] , \g[34][2] , \g[34][1] , 
        SYNOPSYS_UNCONNECTED__13}) );
  FullAdder \level1[14].x6  ( .a({\p[42][63] , n351, n353, n357, n360, n363, 
        n366, n368, n370, n372, n374, n376, n378, n382, n385, n388, n391, n394, 
        n397, n400, n403, n406, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n351, 
        n355, n357, n361, n364, n367, n369, n371, n373, n375, n377, n379, n383, 
        n385, n388, n391, n394, n397, n401, n403, n407, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .cin({n355, n356, n359, n362, n365, n368, n370, 
        n372, n374, n376, n378, n381, n384, n387, n390, n393, n396, n399, n402, 
        n405, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({
        \g[14][63] , \g[14][62] , \g[14][61] , \g[14][60] , \g[14][59] , 
        \g[14][58] , \g[14][57] , \g[14][56] , \g[14][55] , \g[14][54] , 
        \g[14][53] , \g[14][52] , \g[14][51] , \g[14][50] , \g[14][49] , 
        \g[14][48] , \g[14][47] , \g[14][46] , \g[14][45] , \g[14][44] , 
        \g[14][43] , \g[14][42] , \g[14][41] , \g[14][40] , \g[14][39] , 
        \g[14][38] , \g[14][37] , \g[14][36] , \g[14][35] , \g[14][34] , 
        \g[14][33] , \g[14][32] , \g[14][31] , \g[14][30] , \g[14][29] , 
        \g[14][28] , \g[14][27] , \g[14][26] , \g[14][25] , \g[14][24] , 
        \g[14][23] , \g[14][22] , \g[14][21] , \g[14][20] , \g[14][19] , 
        \g[14][18] , \g[14][17] , \g[14][16] , \g[14][15] , \g[14][14] , 
        \g[14][13] , \g[14][12] , \g[14][11] , \g[14][10] , \g[14][9] , 
        \g[14][8] , \g[14][7] , \g[14][6] , \g[14][5] , \g[14][4] , \g[14][3] , 
        \g[14][2] , \g[14][1] , \g[14][0] }), .cout({\g[35][63] , \g[35][62] , 
        \g[35][61] , \g[35][60] , \g[35][59] , \g[35][58] , \g[35][57] , 
        \g[35][56] , \g[35][55] , \g[35][54] , \g[35][53] , \g[35][52] , 
        \g[35][51] , \g[35][50] , \g[35][49] , \g[35][48] , \g[35][47] , 
        \g[35][46] , \g[35][45] , \g[35][44] , \g[35][43] , \g[35][42] , 
        \g[35][41] , \g[35][40] , \g[35][39] , \g[35][38] , \g[35][37] , 
        \g[35][36] , \g[35][35] , \g[35][34] , \g[35][33] , \g[35][32] , 
        \g[35][31] , \g[35][30] , \g[35][29] , \g[35][28] , \g[35][27] , 
        \g[35][26] , \g[35][25] , \g[35][24] , \g[35][23] , \g[35][22] , 
        \g[35][21] , \g[35][20] , \g[35][19] , \g[35][18] , \g[35][17] , 
        \g[35][16] , \g[35][15] , \g[35][14] , \g[35][13] , \g[35][12] , 
        \g[35][11] , \g[35][10] , \g[35][9] , \g[35][8] , \g[35][7] , 
        \g[35][6] , \g[35][5] , \g[35][4] , \g[35][3] , \g[35][2] , \g[35][1] , 
        SYNOPSYS_UNCONNECTED__14}) );
  FullAdder \level1[15].x6  ( .a({n358, n360, n362, n366, n368, n370, n372, 
        n374, n376, n379, n382, n385, n387, n391, n393, n397, n400, n403, n406, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n361, n364, 
        n367, n369, n371, n373, n375, n377, n379, n383, n385, n388, n391, n394, 
        n397, n401, n403, n406, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n364, n365, n368, n370, n372, n374, n376, n378, 
        n381, n384, n387, n390, n393, n396, n399, n402, n405, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[15][63] , 
        \g[15][62] , \g[15][61] , \g[15][60] , \g[15][59] , \g[15][58] , 
        \g[15][57] , \g[15][56] , \g[15][55] , \g[15][54] , \g[15][53] , 
        \g[15][52] , \g[15][51] , \g[15][50] , \g[15][49] , \g[15][48] , 
        \g[15][47] , \g[15][46] , \g[15][45] , \g[15][44] , \g[15][43] , 
        \g[15][42] , \g[15][41] , \g[15][40] , \g[15][39] , \g[15][38] , 
        \g[15][37] , \g[15][36] , \g[15][35] , \g[15][34] , \g[15][33] , 
        \g[15][32] , \g[15][31] , \g[15][30] , \g[15][29] , \g[15][28] , 
        \g[15][27] , \g[15][26] , \g[15][25] , \g[15][24] , \g[15][23] , 
        \g[15][22] , \g[15][21] , \g[15][20] , \g[15][19] , \g[15][18] , 
        \g[15][17] , \g[15][16] , \g[15][15] , \g[15][14] , \g[15][13] , 
        \g[15][12] , \g[15][11] , \g[15][10] , \g[15][9] , \g[15][8] , 
        \g[15][7] , \g[15][6] , \g[15][5] , \g[15][4] , \g[15][3] , \g[15][2] , 
        \g[15][1] , \g[15][0] }), .cout({\g[36][63] , \g[36][62] , \g[36][61] , 
        \g[36][60] , \g[36][59] , \g[36][58] , \g[36][57] , \g[36][56] , 
        \g[36][55] , \g[36][54] , \g[36][53] , \g[36][52] , \g[36][51] , 
        \g[36][50] , \g[36][49] , \g[36][48] , \g[36][47] , \g[36][46] , 
        \g[36][45] , \g[36][44] , \g[36][43] , \g[36][42] , \g[36][41] , 
        \g[36][40] , \g[36][39] , \g[36][38] , \g[36][37] , \g[36][36] , 
        \g[36][35] , \g[36][34] , \g[36][33] , \g[36][32] , \g[36][31] , 
        \g[36][30] , \g[36][29] , \g[36][28] , \g[36][27] , \g[36][26] , 
        \g[36][25] , \g[36][24] , \g[36][23] , \g[36][22] , \g[36][21] , 
        \g[36][20] , \g[36][19] , \g[36][18] , \g[36][17] , \g[36][16] , 
        \g[36][15] , \g[36][14] , \g[36][13] , \g[36][12] , \g[36][11] , 
        \g[36][10] , \g[36][9] , \g[36][8] , \g[36][7] , \g[36][6] , 
        \g[36][5] , \g[36][4] , \g[36][3] , \g[36][2] , \g[36][1] , 
        SYNOPSYS_UNCONNECTED__15}) );
  FullAdder \level1[16].x6  ( .a({n367, n368, n370, n372, n374, n376, n379, 
        n381, n385, n388, n391, n394, n397, n400, n403, n406, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n369, n371, 
        n373, n375, n377, n379, n383, n385, n388, n391, n394, n397, n401, n403, 
        n406, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n371, n372, n374, n376, n378, n380, n384, n387, 
        n390, n393, n396, n399, n402, n405, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[16][63] , 
        \g[16][62] , \g[16][61] , \g[16][60] , \g[16][59] , \g[16][58] , 
        \g[16][57] , \g[16][56] , \g[16][55] , \g[16][54] , \g[16][53] , 
        \g[16][52] , \g[16][51] , \g[16][50] , \g[16][49] , \g[16][48] , 
        \g[16][47] , \g[16][46] , \g[16][45] , \g[16][44] , \g[16][43] , 
        \g[16][42] , \g[16][41] , \g[16][40] , \g[16][39] , \g[16][38] , 
        \g[16][37] , \g[16][36] , \g[16][35] , \g[16][34] , \g[16][33] , 
        \g[16][32] , \g[16][31] , \g[16][30] , \g[16][29] , \g[16][28] , 
        \g[16][27] , \g[16][26] , \g[16][25] , \g[16][24] , \g[16][23] , 
        \g[16][22] , \g[16][21] , \g[16][20] , \g[16][19] , \g[16][18] , 
        \g[16][17] , \g[16][16] , \g[16][15] , \g[16][14] , \g[16][13] , 
        \g[16][12] , \g[16][11] , \g[16][10] , \g[16][9] , \g[16][8] , 
        \g[16][7] , \g[16][6] , \g[16][5] , \g[16][4] , \g[16][3] , \g[16][2] , 
        \g[16][1] , \g[16][0] }), .cout({\g[37][63] , \g[37][62] , \g[37][61] , 
        \g[37][60] , \g[37][59] , \g[37][58] , \g[37][57] , \g[37][56] , 
        \g[37][55] , \g[37][54] , \g[37][53] , \g[37][52] , \g[37][51] , 
        \g[37][50] , \g[37][49] , \g[37][48] , \g[37][47] , \g[37][46] , 
        \g[37][45] , \g[37][44] , \g[37][43] , \g[37][42] , \g[37][41] , 
        \g[37][40] , \g[37][39] , \g[37][38] , \g[37][37] , \g[37][36] , 
        \g[37][35] , \g[37][34] , \g[37][33] , \g[37][32] , \g[37][31] , 
        \g[37][30] , \g[37][29] , \g[37][28] , \g[37][27] , \g[37][26] , 
        \g[37][25] , \g[37][24] , \g[37][23] , \g[37][22] , \g[37][21] , 
        \g[37][20] , \g[37][19] , \g[37][18] , \g[37][17] , \g[37][16] , 
        \g[37][15] , \g[37][14] , \g[37][13] , \g[37][12] , \g[37][11] , 
        \g[37][10] , \g[37][9] , \g[37][8] , \g[37][7] , \g[37][6] , 
        \g[37][5] , \g[37][4] , \g[37][3] , \g[37][2] , \g[37][1] , 
        SYNOPSYS_UNCONNECTED__16}) );
  FullAdder \level1[17].x6  ( .a({n373, n374, n376, n379, n381, n384, n387, 
        n391, n393, n397, n400, n402, n406, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n375, n377, 
        n379, n382, n385, n388, n391, n394, n398, n400, n403, n406, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n377, n378, n380, n384, n387, n390, n393, n396, 
        n399, n402, n405, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[17][63] , 
        \g[17][62] , \g[17][61] , \g[17][60] , \g[17][59] , \g[17][58] , 
        \g[17][57] , \g[17][56] , \g[17][55] , \g[17][54] , \g[17][53] , 
        \g[17][52] , \g[17][51] , \g[17][50] , \g[17][49] , \g[17][48] , 
        \g[17][47] , \g[17][46] , \g[17][45] , \g[17][44] , \g[17][43] , 
        \g[17][42] , \g[17][41] , \g[17][40] , \g[17][39] , \g[17][38] , 
        \g[17][37] , \g[17][36] , \g[17][35] , \g[17][34] , \g[17][33] , 
        \g[17][32] , \g[17][31] , \g[17][30] , \g[17][29] , \g[17][28] , 
        \g[17][27] , \g[17][26] , \g[17][25] , \g[17][24] , \g[17][23] , 
        \g[17][22] , \g[17][21] , \g[17][20] , \g[17][19] , \g[17][18] , 
        \g[17][17] , \g[17][16] , \g[17][15] , \g[17][14] , \g[17][13] , 
        \g[17][12] , \g[17][11] , \g[17][10] , \g[17][9] , \g[17][8] , 
        \g[17][7] , \g[17][6] , \g[17][5] , \g[17][4] , \g[17][3] , \g[17][2] , 
        \g[17][1] , \g[17][0] }), .cout({\g[38][63] , \g[38][62] , \g[38][61] , 
        \g[38][60] , \g[38][59] , \g[38][58] , \g[38][57] , \g[38][56] , 
        \g[38][55] , \g[38][54] , \g[38][53] , \g[38][52] , \g[38][51] , 
        \g[38][50] , \g[38][49] , \g[38][48] , \g[38][47] , \g[38][46] , 
        \g[38][45] , \g[38][44] , \g[38][43] , \g[38][42] , \g[38][41] , 
        \g[38][40] , \g[38][39] , \g[38][38] , \g[38][37] , \g[38][36] , 
        \g[38][35] , \g[38][34] , \g[38][33] , \g[38][32] , \g[38][31] , 
        \g[38][30] , \g[38][29] , \g[38][28] , \g[38][27] , \g[38][26] , 
        \g[38][25] , \g[38][24] , \g[38][23] , \g[38][22] , \g[38][21] , 
        \g[38][20] , \g[38][19] , \g[38][18] , \g[38][17] , \g[38][16] , 
        \g[38][15] , \g[38][14] , \g[38][13] , \g[38][12] , \g[38][11] , 
        \g[38][10] , \g[38][9] , \g[38][8] , \g[38][7] , \g[38][6] , 
        \g[38][5] , \g[38][4] , \g[38][3] , \g[38][2] , \g[38][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  FullAdder \level1[18].x6  ( .a({n379, n382, n384, n387, n391, n393, n397, 
        n400, n403, n406, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n383, n385, 
        n388, n391, n395, n398, n400, n404, n407, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n386, n387, n390, n393, n396, n399, n402, n405, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[18][63] , 
        \g[18][62] , \g[18][61] , \g[18][60] , \g[18][59] , \g[18][58] , 
        \g[18][57] , \g[18][56] , \g[18][55] , \g[18][54] , \g[18][53] , 
        \g[18][52] , \g[18][51] , \g[18][50] , \g[18][49] , \g[18][48] , 
        \g[18][47] , \g[18][46] , \g[18][45] , \g[18][44] , \g[18][43] , 
        \g[18][42] , \g[18][41] , \g[18][40] , \g[18][39] , \g[18][38] , 
        \g[18][37] , \g[18][36] , \g[18][35] , \g[18][34] , \g[18][33] , 
        \g[18][32] , \g[18][31] , \g[18][30] , \g[18][29] , \g[18][28] , 
        \g[18][27] , \g[18][26] , \g[18][25] , \g[18][24] , \g[18][23] , 
        \g[18][22] , \g[18][21] , \g[18][20] , \g[18][19] , \g[18][18] , 
        \g[18][17] , \g[18][16] , \g[18][15] , \g[18][14] , \g[18][13] , 
        \g[18][12] , \g[18][11] , \g[18][10] , \g[18][9] , \g[18][8] , 
        \g[18][7] , \g[18][6] , \g[18][5] , \g[18][4] , \g[18][3] , \g[18][2] , 
        \g[18][1] , \g[18][0] }), .cout({\g[39][63] , \g[39][62] , \g[39][61] , 
        \g[39][60] , \g[39][59] , \g[39][58] , \g[39][57] , \g[39][56] , 
        \g[39][55] , \g[39][54] , \g[39][53] , \g[39][52] , \g[39][51] , 
        \g[39][50] , \g[39][49] , \g[39][48] , \g[39][47] , \g[39][46] , 
        \g[39][45] , \g[39][44] , \g[39][43] , \g[39][42] , \g[39][41] , 
        \g[39][40] , \g[39][39] , \g[39][38] , \g[39][37] , \g[39][36] , 
        \g[39][35] , \g[39][34] , \g[39][33] , \g[39][32] , \g[39][31] , 
        \g[39][30] , \g[39][29] , \g[39][28] , \g[39][27] , \g[39][26] , 
        \g[39][25] , \g[39][24] , \g[39][23] , \g[39][22] , \g[39][21] , 
        \g[39][20] , \g[39][19] , \g[39][18] , \g[39][17] , \g[39][16] , 
        \g[39][15] , \g[39][14] , \g[39][13] , \g[39][12] , \g[39][11] , 
        \g[39][10] , \g[39][9] , \g[39][8] , \g[39][7] , \g[39][6] , 
        \g[39][5] , \g[39][4] , \g[39][3] , \g[39][2] , \g[39][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  FullAdder \level1[19].x6  ( .a({n389, n391, n394, n397, n399, n402, n405, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n392, n395, 
        n398, n400, n404, n407, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n395, n396, n399, n402, n405, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[19][63] , 
        \g[19][62] , \g[19][61] , \g[19][60] , \g[19][59] , \g[19][58] , 
        \g[19][57] , \g[19][56] , \g[19][55] , \g[19][54] , \g[19][53] , 
        \g[19][52] , \g[19][51] , \g[19][50] , \g[19][49] , \g[19][48] , 
        \g[19][47] , \g[19][46] , \g[19][45] , \g[19][44] , \g[19][43] , 
        \g[19][42] , \g[19][41] , \g[19][40] , \g[19][39] , \g[19][38] , 
        \g[19][37] , \g[19][36] , \g[19][35] , \g[19][34] , \g[19][33] , 
        \g[19][32] , \g[19][31] , \g[19][30] , \g[19][29] , \g[19][28] , 
        \g[19][27] , \g[19][26] , \g[19][25] , \g[19][24] , \g[19][23] , 
        \g[19][22] , \g[19][21] , \g[19][20] , \g[19][19] , \g[19][18] , 
        \g[19][17] , \g[19][16] , \g[19][15] , \g[19][14] , \g[19][13] , 
        \g[19][12] , \g[19][11] , \g[19][10] , \g[19][9] , \g[19][8] , 
        \g[19][7] , \g[19][6] , \g[19][5] , \g[19][4] , \g[19][3] , \g[19][2] , 
        \g[19][1] , \g[19][0] }), .cout({\g[40][63] , \g[40][62] , \g[40][61] , 
        \g[40][60] , \g[40][59] , \g[40][58] , \g[40][57] , \g[40][56] , 
        \g[40][55] , \g[40][54] , \g[40][53] , \g[40][52] , \g[40][51] , 
        \g[40][50] , \g[40][49] , \g[40][48] , \g[40][47] , \g[40][46] , 
        \g[40][45] , \g[40][44] , \g[40][43] , \g[40][42] , \g[40][41] , 
        \g[40][40] , \g[40][39] , \g[40][38] , \g[40][37] , \g[40][36] , 
        \g[40][35] , \g[40][34] , \g[40][33] , \g[40][32] , \g[40][31] , 
        \g[40][30] , \g[40][29] , \g[40][28] , \g[40][27] , \g[40][26] , 
        \g[40][25] , \g[40][24] , \g[40][23] , \g[40][22] , \g[40][21] , 
        \g[40][20] , \g[40][19] , \g[40][18] , \g[40][17] , \g[40][16] , 
        \g[40][15] , \g[40][14] , \g[40][13] , \g[40][12] , \g[40][11] , 
        \g[40][10] , \g[40][9] , \g[40][8] , \g[40][7] , \g[40][6] , 
        \g[40][5] , \g[40][4] , \g[40][3] , \g[40][2] , \g[40][1] , 
        SYNOPSYS_UNCONNECTED__19}) );
  FullAdder \level1[20].x6  ( .a({n398, n400, n403, n406, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n401, n404, 
        n407, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n404, n405, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[20][63] , 
        \g[20][62] , \g[20][61] , \g[20][60] , \g[20][59] , \g[20][58] , 
        \g[20][57] , \g[20][56] , \g[20][55] , \g[20][54] , \g[20][53] , 
        \g[20][52] , \g[20][51] , \g[20][50] , \g[20][49] , \g[20][48] , 
        \g[20][47] , \g[20][46] , \g[20][45] , \g[20][44] , \g[20][43] , 
        \g[20][42] , \g[20][41] , \g[20][40] , \g[20][39] , \g[20][38] , 
        \g[20][37] , \g[20][36] , \g[20][35] , \g[20][34] , \g[20][33] , 
        \g[20][32] , \g[20][31] , \g[20][30] , \g[20][29] , \g[20][28] , 
        \g[20][27] , \g[20][26] , \g[20][25] , \g[20][24] , \g[20][23] , 
        \g[20][22] , \g[20][21] , \g[20][20] , \g[20][19] , \g[20][18] , 
        \g[20][17] , \g[20][16] , \g[20][15] , \g[20][14] , \g[20][13] , 
        \g[20][12] , \g[20][11] , \g[20][10] , \g[20][9] , \g[20][8] , 
        \g[20][7] , \g[20][6] , \g[20][5] , \g[20][4] , \g[20][3] , \g[20][2] , 
        \g[20][1] , \g[20][0] }), .cout({\g[41][63] , \g[41][62] , \g[41][61] , 
        \g[41][60] , \g[41][59] , \g[41][58] , \g[41][57] , \g[41][56] , 
        \g[41][55] , \g[41][54] , \g[41][53] , \g[41][52] , \g[41][51] , 
        \g[41][50] , \g[41][49] , \g[41][48] , \g[41][47] , \g[41][46] , 
        \g[41][45] , \g[41][44] , \g[41][43] , \g[41][42] , \g[41][41] , 
        \g[41][40] , \g[41][39] , \g[41][38] , \g[41][37] , \g[41][36] , 
        \g[41][35] , \g[41][34] , \g[41][33] , \g[41][32] , \g[41][31] , 
        \g[41][30] , \g[41][29] , \g[41][28] , \g[41][27] , \g[41][26] , 
        \g[41][25] , \g[41][24] , \g[41][23] , \g[41][22] , \g[41][21] , 
        \g[41][20] , \g[41][19] , \g[41][18] , \g[41][17] , \g[41][16] , 
        \g[41][15] , \g[41][14] , \g[41][13] , \g[41][12] , \g[41][11] , 
        \g[41][10] , \g[41][9] , \g[41][8] , \g[41][7] , \g[41][6] , 
        \g[41][5] , \g[41][4] , \g[41][3] , \g[41][2] , \g[41][1] , 
        SYNOPSYS_UNCONNECTED__20}) );
  FullAdder \level2[0].x5  ( .a({\g[0][63] , \g[0][62] , \g[0][61] , 
        \g[0][60] , \g[0][59] , \g[0][58] , \g[0][57] , \g[0][56] , \g[0][55] , 
        \g[0][54] , \g[0][53] , \g[0][52] , \g[0][51] , \g[0][50] , \g[0][49] , 
        \g[0][48] , \g[0][47] , \g[0][46] , \g[0][45] , \g[0][44] , \g[0][43] , 
        \g[0][42] , \g[0][41] , \g[0][40] , \g[0][39] , \g[0][38] , \g[0][37] , 
        \g[0][36] , \g[0][35] , \g[0][34] , \g[0][33] , \g[0][32] , \g[0][31] , 
        \g[0][30] , \g[0][29] , \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] , 
        \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , \g[0][19] , 
        \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] , \g[0][13] , 
        \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] , \g[0][7] , 
        \g[0][6] , \g[0][5] , \g[0][4] , \g[0][3] , \g[0][2] , \g[0][1] , 
        \g[0][0] }), .b({\g[1][63] , \g[1][62] , \g[1][61] , \g[1][60] , 
        \g[1][59] , \g[1][58] , \g[1][57] , \g[1][56] , \g[1][55] , \g[1][54] , 
        \g[1][53] , \g[1][52] , \g[1][51] , \g[1][50] , \g[1][49] , \g[1][48] , 
        \g[1][47] , \g[1][46] , \g[1][45] , \g[1][44] , \g[1][43] , \g[1][42] , 
        \g[1][41] , \g[1][40] , \g[1][39] , \g[1][38] , \g[1][37] , \g[1][36] , 
        \g[1][35] , \g[1][34] , \g[1][33] , \g[1][32] , \g[1][31] , \g[1][30] , 
        \g[1][29] , \g[1][28] , \g[1][27] , \g[1][26] , \g[1][25] , \g[1][24] , 
        \g[1][23] , \g[1][22] , \g[1][21] , \g[1][20] , \g[1][19] , \g[1][18] , 
        \g[1][17] , \g[1][16] , \g[1][15] , \g[1][14] , \g[1][13] , \g[1][12] , 
        \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] , \g[1][6] , 
        \g[1][5] , \g[1][4] , \g[1][3] , \g[1][2] , \g[1][1] , \g[1][0] }), 
        .cin({\g[2][63] , \g[2][62] , \g[2][61] , \g[2][60] , \g[2][59] , 
        \g[2][58] , \g[2][57] , \g[2][56] , \g[2][55] , \g[2][54] , \g[2][53] , 
        \g[2][52] , \g[2][51] , \g[2][50] , \g[2][49] , \g[2][48] , \g[2][47] , 
        \g[2][46] , \g[2][45] , \g[2][44] , \g[2][43] , \g[2][42] , \g[2][41] , 
        \g[2][40] , \g[2][39] , \g[2][38] , \g[2][37] , \g[2][36] , \g[2][35] , 
        \g[2][34] , \g[2][33] , \g[2][32] , \g[2][31] , \g[2][30] , \g[2][29] , 
        \g[2][28] , \g[2][27] , \g[2][26] , \g[2][25] , \g[2][24] , \g[2][23] , 
        \g[2][22] , \g[2][21] , \g[2][20] , \g[2][19] , \g[2][18] , \g[2][17] , 
        \g[2][16] , \g[2][15] , \g[2][14] , \g[2][13] , \g[2][12] , \g[2][11] , 
        \g[2][10] , \g[2][9] , \g[2][8] , \g[2][7] , \g[2][6] , \g[2][5] , 
        \g[2][4] , \g[2][3] , \g[2][2] , \g[2][1] , \g[2][0] }), .sum({
        \g2[0][63] , \g2[0][62] , \g2[0][61] , \g2[0][60] , \g2[0][59] , 
        \g2[0][58] , \g2[0][57] , \g2[0][56] , \g2[0][55] , \g2[0][54] , 
        \g2[0][53] , \g2[0][52] , \g2[0][51] , \g2[0][50] , \g2[0][49] , 
        \g2[0][48] , \g2[0][47] , \g2[0][46] , \g2[0][45] , \g2[0][44] , 
        \g2[0][43] , \g2[0][42] , \g2[0][41] , \g2[0][40] , \g2[0][39] , 
        \g2[0][38] , \g2[0][37] , \g2[0][36] , \g2[0][35] , \g2[0][34] , 
        \g2[0][33] , \g2[0][32] , \g2[0][31] , \g2[0][30] , \g2[0][29] , 
        \g2[0][28] , \g2[0][27] , \g2[0][26] , \g2[0][25] , \g2[0][24] , 
        \g2[0][23] , \g2[0][22] , \g2[0][21] , \g2[0][20] , \g2[0][19] , 
        \g2[0][18] , \g2[0][17] , \g2[0][16] , \g2[0][15] , \g2[0][14] , 
        \g2[0][13] , \g2[0][12] , \g2[0][11] , \g2[0][10] , \g2[0][9] , 
        \g2[0][8] , \g2[0][7] , \g2[0][6] , \g2[0][5] , \g2[0][4] , \g2[0][3] , 
        \g2[0][2] , \g2[0][1] , \g2[0][0] }), .cout({\g2[14][63] , 
        \g2[14][62] , \g2[14][61] , \g2[14][60] , \g2[14][59] , \g2[14][58] , 
        \g2[14][57] , \g2[14][56] , \g2[14][55] , \g2[14][54] , \g2[14][53] , 
        \g2[14][52] , \g2[14][51] , \g2[14][50] , \g2[14][49] , \g2[14][48] , 
        \g2[14][47] , \g2[14][46] , \g2[14][45] , \g2[14][44] , \g2[14][43] , 
        \g2[14][42] , \g2[14][41] , \g2[14][40] , \g2[14][39] , \g2[14][38] , 
        \g2[14][37] , \g2[14][36] , \g2[14][35] , \g2[14][34] , \g2[14][33] , 
        \g2[14][32] , \g2[14][31] , \g2[14][30] , \g2[14][29] , \g2[14][28] , 
        \g2[14][27] , \g2[14][26] , \g2[14][25] , \g2[14][24] , \g2[14][23] , 
        \g2[14][22] , \g2[14][21] , \g2[14][20] , \g2[14][19] , \g2[14][18] , 
        \g2[14][17] , \g2[14][16] , \g2[14][15] , \g2[14][14] , \g2[14][13] , 
        \g2[14][12] , \g2[14][11] , \g2[14][10] , \g2[14][9] , \g2[14][8] , 
        \g2[14][7] , \g2[14][6] , \g2[14][5] , \g2[14][4] , \g2[14][3] , 
        \g2[14][2] , \g2[14][1] , SYNOPSYS_UNCONNECTED__21}) );
  FullAdder \level2[1].x5  ( .a({\g[3][63] , \g[3][62] , \g[3][61] , 
        \g[3][60] , \g[3][59] , \g[3][58] , \g[3][57] , \g[3][56] , \g[3][55] , 
        \g[3][54] , \g[3][53] , \g[3][52] , \g[3][51] , \g[3][50] , \g[3][49] , 
        \g[3][48] , \g[3][47] , \g[3][46] , \g[3][45] , \g[3][44] , \g[3][43] , 
        \g[3][42] , \g[3][41] , \g[3][40] , \g[3][39] , \g[3][38] , \g[3][37] , 
        \g[3][36] , \g[3][35] , \g[3][34] , \g[3][33] , \g[3][32] , \g[3][31] , 
        \g[3][30] , \g[3][29] , \g[3][28] , \g[3][27] , \g[3][26] , \g[3][25] , 
        \g[3][24] , \g[3][23] , \g[3][22] , \g[3][21] , \g[3][20] , \g[3][19] , 
        \g[3][18] , \g[3][17] , \g[3][16] , \g[3][15] , \g[3][14] , \g[3][13] , 
        \g[3][12] , \g[3][11] , \g[3][10] , \g[3][9] , \g[3][8] , \g[3][7] , 
        \g[3][6] , \g[3][5] , \g[3][4] , \g[3][3] , \g[3][2] , \g[3][1] , 
        \g[3][0] }), .b({\g[4][63] , \g[4][62] , \g[4][61] , \g[4][60] , 
        \g[4][59] , \g[4][58] , \g[4][57] , \g[4][56] , \g[4][55] , \g[4][54] , 
        \g[4][53] , \g[4][52] , \g[4][51] , \g[4][50] , \g[4][49] , \g[4][48] , 
        \g[4][47] , \g[4][46] , \g[4][45] , \g[4][44] , \g[4][43] , \g[4][42] , 
        \g[4][41] , \g[4][40] , \g[4][39] , \g[4][38] , \g[4][37] , \g[4][36] , 
        \g[4][35] , \g[4][34] , \g[4][33] , \g[4][32] , \g[4][31] , \g[4][30] , 
        \g[4][29] , \g[4][28] , \g[4][27] , \g[4][26] , \g[4][25] , \g[4][24] , 
        \g[4][23] , \g[4][22] , \g[4][21] , \g[4][20] , \g[4][19] , \g[4][18] , 
        \g[4][17] , \g[4][16] , \g[4][15] , \g[4][14] , \g[4][13] , \g[4][12] , 
        \g[4][11] , \g[4][10] , \g[4][9] , \g[4][8] , \g[4][7] , \g[4][6] , 
        \g[4][5] , \g[4][4] , \g[4][3] , \g[4][2] , \g[4][1] , \g[4][0] }), 
        .cin({\g[5][63] , \g[5][62] , \g[5][61] , \g[5][60] , \g[5][59] , 
        \g[5][58] , \g[5][57] , \g[5][56] , \g[5][55] , \g[5][54] , \g[5][53] , 
        \g[5][52] , \g[5][51] , \g[5][50] , \g[5][49] , \g[5][48] , \g[5][47] , 
        \g[5][46] , \g[5][45] , \g[5][44] , \g[5][43] , \g[5][42] , \g[5][41] , 
        \g[5][40] , \g[5][39] , \g[5][38] , \g[5][37] , \g[5][36] , \g[5][35] , 
        \g[5][34] , \g[5][33] , \g[5][32] , \g[5][31] , \g[5][30] , \g[5][29] , 
        \g[5][28] , \g[5][27] , \g[5][26] , \g[5][25] , \g[5][24] , \g[5][23] , 
        \g[5][22] , \g[5][21] , \g[5][20] , \g[5][19] , \g[5][18] , \g[5][17] , 
        \g[5][16] , \g[5][15] , \g[5][14] , \g[5][13] , \g[5][12] , \g[5][11] , 
        \g[5][10] , \g[5][9] , \g[5][8] , \g[5][7] , \g[5][6] , \g[5][5] , 
        \g[5][4] , \g[5][3] , \g[5][2] , \g[5][1] , \g[5][0] }), .sum({
        \g2[1][63] , \g2[1][62] , \g2[1][61] , \g2[1][60] , \g2[1][59] , 
        \g2[1][58] , \g2[1][57] , \g2[1][56] , \g2[1][55] , \g2[1][54] , 
        \g2[1][53] , \g2[1][52] , \g2[1][51] , \g2[1][50] , \g2[1][49] , 
        \g2[1][48] , \g2[1][47] , \g2[1][46] , \g2[1][45] , \g2[1][44] , 
        \g2[1][43] , \g2[1][42] , \g2[1][41] , \g2[1][40] , \g2[1][39] , 
        \g2[1][38] , \g2[1][37] , \g2[1][36] , \g2[1][35] , \g2[1][34] , 
        \g2[1][33] , \g2[1][32] , \g2[1][31] , \g2[1][30] , \g2[1][29] , 
        \g2[1][28] , \g2[1][27] , \g2[1][26] , \g2[1][25] , \g2[1][24] , 
        \g2[1][23] , \g2[1][22] , \g2[1][21] , \g2[1][20] , \g2[1][19] , 
        \g2[1][18] , \g2[1][17] , \g2[1][16] , \g2[1][15] , \g2[1][14] , 
        \g2[1][13] , \g2[1][12] , \g2[1][11] , \g2[1][10] , \g2[1][9] , 
        \g2[1][8] , \g2[1][7] , \g2[1][6] , \g2[1][5] , \g2[1][4] , \g2[1][3] , 
        \g2[1][2] , \g2[1][1] , \g2[1][0] }), .cout({\g2[15][63] , 
        \g2[15][62] , \g2[15][61] , \g2[15][60] , \g2[15][59] , \g2[15][58] , 
        \g2[15][57] , \g2[15][56] , \g2[15][55] , \g2[15][54] , \g2[15][53] , 
        \g2[15][52] , \g2[15][51] , \g2[15][50] , \g2[15][49] , \g2[15][48] , 
        \g2[15][47] , \g2[15][46] , \g2[15][45] , \g2[15][44] , \g2[15][43] , 
        \g2[15][42] , \g2[15][41] , \g2[15][40] , \g2[15][39] , \g2[15][38] , 
        \g2[15][37] , \g2[15][36] , \g2[15][35] , \g2[15][34] , \g2[15][33] , 
        \g2[15][32] , \g2[15][31] , \g2[15][30] , \g2[15][29] , \g2[15][28] , 
        \g2[15][27] , \g2[15][26] , \g2[15][25] , \g2[15][24] , \g2[15][23] , 
        \g2[15][22] , \g2[15][21] , \g2[15][20] , \g2[15][19] , \g2[15][18] , 
        \g2[15][17] , \g2[15][16] , \g2[15][15] , \g2[15][14] , \g2[15][13] , 
        \g2[15][12] , \g2[15][11] , \g2[15][10] , \g2[15][9] , \g2[15][8] , 
        \g2[15][7] , \g2[15][6] , \g2[15][5] , \g2[15][4] , \g2[15][3] , 
        \g2[15][2] , \g2[15][1] , SYNOPSYS_UNCONNECTED__22}) );
  FullAdder \level2[2].x5  ( .a({\g[6][63] , \g[6][62] , \g[6][61] , 
        \g[6][60] , \g[6][59] , \g[6][58] , \g[6][57] , \g[6][56] , \g[6][55] , 
        \g[6][54] , \g[6][53] , \g[6][52] , \g[6][51] , \g[6][50] , \g[6][49] , 
        \g[6][48] , \g[6][47] , \g[6][46] , \g[6][45] , \g[6][44] , \g[6][43] , 
        \g[6][42] , \g[6][41] , \g[6][40] , \g[6][39] , \g[6][38] , \g[6][37] , 
        \g[6][36] , \g[6][35] , \g[6][34] , \g[6][33] , \g[6][32] , \g[6][31] , 
        \g[6][30] , \g[6][29] , \g[6][28] , \g[6][27] , \g[6][26] , \g[6][25] , 
        \g[6][24] , \g[6][23] , \g[6][22] , \g[6][21] , \g[6][20] , \g[6][19] , 
        \g[6][18] , \g[6][17] , \g[6][16] , \g[6][15] , \g[6][14] , \g[6][13] , 
        \g[6][12] , \g[6][11] , \g[6][10] , \g[6][9] , \g[6][8] , \g[6][7] , 
        \g[6][6] , \g[6][5] , \g[6][4] , \g[6][3] , \g[6][2] , \g[6][1] , 
        \g[6][0] }), .b({\g[7][63] , \g[7][62] , \g[7][61] , \g[7][60] , 
        \g[7][59] , \g[7][58] , \g[7][57] , \g[7][56] , \g[7][55] , \g[7][54] , 
        \g[7][53] , \g[7][52] , \g[7][51] , \g[7][50] , \g[7][49] , \g[7][48] , 
        \g[7][47] , \g[7][46] , \g[7][45] , \g[7][44] , \g[7][43] , \g[7][42] , 
        \g[7][41] , \g[7][40] , \g[7][39] , \g[7][38] , \g[7][37] , \g[7][36] , 
        \g[7][35] , \g[7][34] , \g[7][33] , \g[7][32] , \g[7][31] , \g[7][30] , 
        \g[7][29] , \g[7][28] , \g[7][27] , \g[7][26] , \g[7][25] , \g[7][24] , 
        \g[7][23] , \g[7][22] , \g[7][21] , \g[7][20] , \g[7][19] , \g[7][18] , 
        \g[7][17] , \g[7][16] , \g[7][15] , \g[7][14] , \g[7][13] , \g[7][12] , 
        \g[7][11] , \g[7][10] , \g[7][9] , \g[7][8] , \g[7][7] , \g[7][6] , 
        \g[7][5] , \g[7][4] , \g[7][3] , \g[7][2] , \g[7][1] , \g[7][0] }), 
        .cin({\g[8][63] , \g[8][62] , \g[8][61] , \g[8][60] , \g[8][59] , 
        \g[8][58] , \g[8][57] , \g[8][56] , \g[8][55] , \g[8][54] , \g[8][53] , 
        \g[8][52] , \g[8][51] , \g[8][50] , \g[8][49] , \g[8][48] , \g[8][47] , 
        \g[8][46] , \g[8][45] , \g[8][44] , \g[8][43] , \g[8][42] , \g[8][41] , 
        \g[8][40] , \g[8][39] , \g[8][38] , \g[8][37] , \g[8][36] , \g[8][35] , 
        \g[8][34] , \g[8][33] , \g[8][32] , \g[8][31] , \g[8][30] , \g[8][29] , 
        \g[8][28] , \g[8][27] , \g[8][26] , \g[8][25] , \g[8][24] , \g[8][23] , 
        \g[8][22] , \g[8][21] , \g[8][20] , \g[8][19] , \g[8][18] , \g[8][17] , 
        \g[8][16] , \g[8][15] , \g[8][14] , \g[8][13] , \g[8][12] , \g[8][11] , 
        \g[8][10] , \g[8][9] , \g[8][8] , \g[8][7] , \g[8][6] , \g[8][5] , 
        \g[8][4] , \g[8][3] , \g[8][2] , \g[8][1] , \g[8][0] }), .sum({
        \g2[2][63] , \g2[2][62] , \g2[2][61] , \g2[2][60] , \g2[2][59] , 
        \g2[2][58] , \g2[2][57] , \g2[2][56] , \g2[2][55] , \g2[2][54] , 
        \g2[2][53] , \g2[2][52] , \g2[2][51] , \g2[2][50] , \g2[2][49] , 
        \g2[2][48] , \g2[2][47] , \g2[2][46] , \g2[2][45] , \g2[2][44] , 
        \g2[2][43] , \g2[2][42] , \g2[2][41] , \g2[2][40] , \g2[2][39] , 
        \g2[2][38] , \g2[2][37] , \g2[2][36] , \g2[2][35] , \g2[2][34] , 
        \g2[2][33] , \g2[2][32] , \g2[2][31] , \g2[2][30] , \g2[2][29] , 
        \g2[2][28] , \g2[2][27] , \g2[2][26] , \g2[2][25] , \g2[2][24] , 
        \g2[2][23] , \g2[2][22] , \g2[2][21] , \g2[2][20] , \g2[2][19] , 
        \g2[2][18] , \g2[2][17] , \g2[2][16] , \g2[2][15] , \g2[2][14] , 
        \g2[2][13] , \g2[2][12] , \g2[2][11] , \g2[2][10] , \g2[2][9] , 
        \g2[2][8] , \g2[2][7] , \g2[2][6] , \g2[2][5] , \g2[2][4] , \g2[2][3] , 
        \g2[2][2] , \g2[2][1] , \g2[2][0] }), .cout({\g2[16][63] , 
        \g2[16][62] , \g2[16][61] , \g2[16][60] , \g2[16][59] , \g2[16][58] , 
        \g2[16][57] , \g2[16][56] , \g2[16][55] , \g2[16][54] , \g2[16][53] , 
        \g2[16][52] , \g2[16][51] , \g2[16][50] , \g2[16][49] , \g2[16][48] , 
        \g2[16][47] , \g2[16][46] , \g2[16][45] , \g2[16][44] , \g2[16][43] , 
        \g2[16][42] , \g2[16][41] , \g2[16][40] , \g2[16][39] , \g2[16][38] , 
        \g2[16][37] , \g2[16][36] , \g2[16][35] , \g2[16][34] , \g2[16][33] , 
        \g2[16][32] , \g2[16][31] , \g2[16][30] , \g2[16][29] , \g2[16][28] , 
        \g2[16][27] , \g2[16][26] , \g2[16][25] , \g2[16][24] , \g2[16][23] , 
        \g2[16][22] , \g2[16][21] , \g2[16][20] , \g2[16][19] , \g2[16][18] , 
        \g2[16][17] , \g2[16][16] , \g2[16][15] , \g2[16][14] , \g2[16][13] , 
        \g2[16][12] , \g2[16][11] , \g2[16][10] , \g2[16][9] , \g2[16][8] , 
        \g2[16][7] , \g2[16][6] , \g2[16][5] , \g2[16][4] , \g2[16][3] , 
        \g2[16][2] , \g2[16][1] , SYNOPSYS_UNCONNECTED__23}) );
  FullAdder \level2[3].x5  ( .a({\g[9][63] , \g[9][62] , \g[9][61] , 
        \g[9][60] , \g[9][59] , \g[9][58] , \g[9][57] , \g[9][56] , \g[9][55] , 
        \g[9][54] , \g[9][53] , \g[9][52] , \g[9][51] , \g[9][50] , \g[9][49] , 
        \g[9][48] , \g[9][47] , \g[9][46] , \g[9][45] , \g[9][44] , \g[9][43] , 
        \g[9][42] , \g[9][41] , \g[9][40] , \g[9][39] , \g[9][38] , \g[9][37] , 
        \g[9][36] , \g[9][35] , \g[9][34] , \g[9][33] , \g[9][32] , \g[9][31] , 
        \g[9][30] , \g[9][29] , \g[9][28] , \g[9][27] , \g[9][26] , \g[9][25] , 
        \g[9][24] , \g[9][23] , \g[9][22] , \g[9][21] , \g[9][20] , \g[9][19] , 
        \g[9][18] , \g[9][17] , \g[9][16] , \g[9][15] , \g[9][14] , \g[9][13] , 
        \g[9][12] , \g[9][11] , \g[9][10] , \g[9][9] , \g[9][8] , \g[9][7] , 
        \g[9][6] , \g[9][5] , \g[9][4] , \g[9][3] , \g[9][2] , \g[9][1] , 
        \g[9][0] }), .b({\g[10][63] , \g[10][62] , \g[10][61] , \g[10][60] , 
        \g[10][59] , \g[10][58] , \g[10][57] , \g[10][56] , \g[10][55] , 
        \g[10][54] , \g[10][53] , \g[10][52] , \g[10][51] , \g[10][50] , 
        \g[10][49] , \g[10][48] , \g[10][47] , \g[10][46] , \g[10][45] , 
        \g[10][44] , \g[10][43] , \g[10][42] , \g[10][41] , \g[10][40] , 
        \g[10][39] , \g[10][38] , \g[10][37] , \g[10][36] , \g[10][35] , 
        \g[10][34] , \g[10][33] , \g[10][32] , \g[10][31] , \g[10][30] , 
        \g[10][29] , \g[10][28] , \g[10][27] , \g[10][26] , \g[10][25] , 
        \g[10][24] , \g[10][23] , \g[10][22] , \g[10][21] , \g[10][20] , 
        \g[10][19] , \g[10][18] , \g[10][17] , \g[10][16] , \g[10][15] , 
        \g[10][14] , \g[10][13] , \g[10][12] , \g[10][11] , \g[10][10] , 
        \g[10][9] , \g[10][8] , \g[10][7] , \g[10][6] , \g[10][5] , \g[10][4] , 
        \g[10][3] , \g[10][2] , \g[10][1] , \g[10][0] }), .cin({\g[11][63] , 
        \g[11][62] , \g[11][61] , \g[11][60] , \g[11][59] , \g[11][58] , 
        \g[11][57] , \g[11][56] , \g[11][55] , \g[11][54] , \g[11][53] , 
        \g[11][52] , \g[11][51] , \g[11][50] , \g[11][49] , \g[11][48] , 
        \g[11][47] , \g[11][46] , \g[11][45] , \g[11][44] , \g[11][43] , 
        \g[11][42] , \g[11][41] , \g[11][40] , \g[11][39] , \g[11][38] , 
        \g[11][37] , \g[11][36] , \g[11][35] , \g[11][34] , \g[11][33] , 
        \g[11][32] , \g[11][31] , \g[11][30] , \g[11][29] , \g[11][28] , 
        \g[11][27] , \g[11][26] , \g[11][25] , \g[11][24] , \g[11][23] , 
        \g[11][22] , \g[11][21] , \g[11][20] , \g[11][19] , \g[11][18] , 
        \g[11][17] , \g[11][16] , \g[11][15] , \g[11][14] , \g[11][13] , 
        \g[11][12] , \g[11][11] , \g[11][10] , \g[11][9] , \g[11][8] , 
        \g[11][7] , \g[11][6] , \g[11][5] , \g[11][4] , \g[11][3] , \g[11][2] , 
        \g[11][1] , \g[11][0] }), .sum({\g2[3][63] , \g2[3][62] , \g2[3][61] , 
        \g2[3][60] , \g2[3][59] , \g2[3][58] , \g2[3][57] , \g2[3][56] , 
        \g2[3][55] , \g2[3][54] , \g2[3][53] , \g2[3][52] , \g2[3][51] , 
        \g2[3][50] , \g2[3][49] , \g2[3][48] , \g2[3][47] , \g2[3][46] , 
        \g2[3][45] , \g2[3][44] , \g2[3][43] , \g2[3][42] , \g2[3][41] , 
        \g2[3][40] , \g2[3][39] , \g2[3][38] , \g2[3][37] , \g2[3][36] , 
        \g2[3][35] , \g2[3][34] , \g2[3][33] , \g2[3][32] , \g2[3][31] , 
        \g2[3][30] , \g2[3][29] , \g2[3][28] , \g2[3][27] , \g2[3][26] , 
        \g2[3][25] , \g2[3][24] , \g2[3][23] , \g2[3][22] , \g2[3][21] , 
        \g2[3][20] , \g2[3][19] , \g2[3][18] , \g2[3][17] , \g2[3][16] , 
        \g2[3][15] , \g2[3][14] , \g2[3][13] , \g2[3][12] , \g2[3][11] , 
        \g2[3][10] , \g2[3][9] , \g2[3][8] , \g2[3][7] , \g2[3][6] , 
        \g2[3][5] , \g2[3][4] , \g2[3][3] , \g2[3][2] , \g2[3][1] , \g2[3][0] }), .cout({\g2[17][63] , \g2[17][62] , \g2[17][61] , \g2[17][60] , \g2[17][59] , 
        \g2[17][58] , \g2[17][57] , \g2[17][56] , \g2[17][55] , \g2[17][54] , 
        \g2[17][53] , \g2[17][52] , \g2[17][51] , \g2[17][50] , \g2[17][49] , 
        \g2[17][48] , \g2[17][47] , \g2[17][46] , \g2[17][45] , \g2[17][44] , 
        \g2[17][43] , \g2[17][42] , \g2[17][41] , \g2[17][40] , \g2[17][39] , 
        \g2[17][38] , \g2[17][37] , \g2[17][36] , \g2[17][35] , \g2[17][34] , 
        \g2[17][33] , \g2[17][32] , \g2[17][31] , \g2[17][30] , \g2[17][29] , 
        \g2[17][28] , \g2[17][27] , \g2[17][26] , \g2[17][25] , \g2[17][24] , 
        \g2[17][23] , \g2[17][22] , \g2[17][21] , \g2[17][20] , \g2[17][19] , 
        \g2[17][18] , \g2[17][17] , \g2[17][16] , \g2[17][15] , \g2[17][14] , 
        \g2[17][13] , \g2[17][12] , \g2[17][11] , \g2[17][10] , \g2[17][9] , 
        \g2[17][8] , \g2[17][7] , \g2[17][6] , \g2[17][5] , \g2[17][4] , 
        \g2[17][3] , \g2[17][2] , \g2[17][1] , SYNOPSYS_UNCONNECTED__24}) );
  FullAdder \level2[4].x5  ( .a({\g[12][63] , \g[12][62] , \g[12][61] , 
        \g[12][60] , \g[12][59] , \g[12][58] , \g[12][57] , \g[12][56] , 
        \g[12][55] , \g[12][54] , \g[12][53] , \g[12][52] , \g[12][51] , 
        \g[12][50] , \g[12][49] , \g[12][48] , \g[12][47] , \g[12][46] , 
        \g[12][45] , \g[12][44] , \g[12][43] , \g[12][42] , \g[12][41] , 
        \g[12][40] , \g[12][39] , \g[12][38] , \g[12][37] , \g[12][36] , 
        \g[12][35] , \g[12][34] , \g[12][33] , \g[12][32] , \g[12][31] , 
        \g[12][30] , \g[12][29] , \g[12][28] , \g[12][27] , \g[12][26] , 
        \g[12][25] , \g[12][24] , \g[12][23] , \g[12][22] , \g[12][21] , 
        \g[12][20] , \g[12][19] , \g[12][18] , \g[12][17] , \g[12][16] , 
        \g[12][15] , \g[12][14] , \g[12][13] , \g[12][12] , \g[12][11] , 
        \g[12][10] , \g[12][9] , \g[12][8] , \g[12][7] , \g[12][6] , 
        \g[12][5] , \g[12][4] , \g[12][3] , \g[12][2] , \g[12][1] , \g[12][0] }), .b({\g[13][63] , \g[13][62] , \g[13][61] , \g[13][60] , \g[13][59] , 
        \g[13][58] , \g[13][57] , \g[13][56] , \g[13][55] , \g[13][54] , 
        \g[13][53] , \g[13][52] , \g[13][51] , \g[13][50] , \g[13][49] , 
        \g[13][48] , \g[13][47] , \g[13][46] , \g[13][45] , \g[13][44] , 
        \g[13][43] , \g[13][42] , \g[13][41] , \g[13][40] , \g[13][39] , 
        \g[13][38] , \g[13][37] , \g[13][36] , \g[13][35] , \g[13][34] , 
        \g[13][33] , \g[13][32] , \g[13][31] , \g[13][30] , \g[13][29] , 
        \g[13][28] , \g[13][27] , \g[13][26] , \g[13][25] , \g[13][24] , 
        \g[13][23] , \g[13][22] , \g[13][21] , \g[13][20] , \g[13][19] , 
        \g[13][18] , \g[13][17] , \g[13][16] , \g[13][15] , \g[13][14] , 
        \g[13][13] , \g[13][12] , \g[13][11] , \g[13][10] , \g[13][9] , 
        \g[13][8] , \g[13][7] , \g[13][6] , \g[13][5] , \g[13][4] , \g[13][3] , 
        \g[13][2] , \g[13][1] , \g[13][0] }), .cin({\g[14][63] , \g[14][62] , 
        \g[14][61] , \g[14][60] , \g[14][59] , \g[14][58] , \g[14][57] , 
        \g[14][56] , \g[14][55] , \g[14][54] , \g[14][53] , \g[14][52] , 
        \g[14][51] , \g[14][50] , \g[14][49] , \g[14][48] , \g[14][47] , 
        \g[14][46] , \g[14][45] , \g[14][44] , \g[14][43] , \g[14][42] , 
        \g[14][41] , \g[14][40] , \g[14][39] , \g[14][38] , \g[14][37] , 
        \g[14][36] , \g[14][35] , \g[14][34] , \g[14][33] , \g[14][32] , 
        \g[14][31] , \g[14][30] , \g[14][29] , \g[14][28] , \g[14][27] , 
        \g[14][26] , \g[14][25] , \g[14][24] , \g[14][23] , \g[14][22] , 
        \g[14][21] , \g[14][20] , \g[14][19] , \g[14][18] , \g[14][17] , 
        \g[14][16] , \g[14][15] , \g[14][14] , \g[14][13] , \g[14][12] , 
        \g[14][11] , \g[14][10] , \g[14][9] , \g[14][8] , \g[14][7] , 
        \g[14][6] , \g[14][5] , \g[14][4] , \g[14][3] , \g[14][2] , \g[14][1] , 
        \g[14][0] }), .sum({\g2[4][63] , \g2[4][62] , \g2[4][61] , \g2[4][60] , 
        \g2[4][59] , \g2[4][58] , \g2[4][57] , \g2[4][56] , \g2[4][55] , 
        \g2[4][54] , \g2[4][53] , \g2[4][52] , \g2[4][51] , \g2[4][50] , 
        \g2[4][49] , \g2[4][48] , \g2[4][47] , \g2[4][46] , \g2[4][45] , 
        \g2[4][44] , \g2[4][43] , \g2[4][42] , \g2[4][41] , \g2[4][40] , 
        \g2[4][39] , \g2[4][38] , \g2[4][37] , \g2[4][36] , \g2[4][35] , 
        \g2[4][34] , \g2[4][33] , \g2[4][32] , \g2[4][31] , \g2[4][30] , 
        \g2[4][29] , \g2[4][28] , \g2[4][27] , \g2[4][26] , \g2[4][25] , 
        \g2[4][24] , \g2[4][23] , \g2[4][22] , \g2[4][21] , \g2[4][20] , 
        \g2[4][19] , \g2[4][18] , \g2[4][17] , \g2[4][16] , \g2[4][15] , 
        \g2[4][14] , \g2[4][13] , \g2[4][12] , \g2[4][11] , \g2[4][10] , 
        \g2[4][9] , \g2[4][8] , \g2[4][7] , \g2[4][6] , \g2[4][5] , \g2[4][4] , 
        \g2[4][3] , \g2[4][2] , \g2[4][1] , \g2[4][0] }), .cout({\g2[18][63] , 
        \g2[18][62] , \g2[18][61] , \g2[18][60] , \g2[18][59] , \g2[18][58] , 
        \g2[18][57] , \g2[18][56] , \g2[18][55] , \g2[18][54] , \g2[18][53] , 
        \g2[18][52] , \g2[18][51] , \g2[18][50] , \g2[18][49] , \g2[18][48] , 
        \g2[18][47] , \g2[18][46] , \g2[18][45] , \g2[18][44] , \g2[18][43] , 
        \g2[18][42] , \g2[18][41] , \g2[18][40] , \g2[18][39] , \g2[18][38] , 
        \g2[18][37] , \g2[18][36] , \g2[18][35] , \g2[18][34] , \g2[18][33] , 
        \g2[18][32] , \g2[18][31] , \g2[18][30] , \g2[18][29] , \g2[18][28] , 
        \g2[18][27] , \g2[18][26] , \g2[18][25] , \g2[18][24] , \g2[18][23] , 
        \g2[18][22] , \g2[18][21] , \g2[18][20] , \g2[18][19] , \g2[18][18] , 
        \g2[18][17] , \g2[18][16] , \g2[18][15] , \g2[18][14] , \g2[18][13] , 
        \g2[18][12] , \g2[18][11] , \g2[18][10] , \g2[18][9] , \g2[18][8] , 
        \g2[18][7] , \g2[18][6] , \g2[18][5] , \g2[18][4] , \g2[18][3] , 
        \g2[18][2] , \g2[18][1] , SYNOPSYS_UNCONNECTED__25}) );
  FullAdder \level2[5].x5  ( .a({\g[15][63] , \g[15][62] , \g[15][61] , 
        \g[15][60] , \g[15][59] , \g[15][58] , \g[15][57] , \g[15][56] , 
        \g[15][55] , \g[15][54] , \g[15][53] , \g[15][52] , \g[15][51] , 
        \g[15][50] , \g[15][49] , \g[15][48] , \g[15][47] , \g[15][46] , 
        \g[15][45] , \g[15][44] , \g[15][43] , \g[15][42] , \g[15][41] , 
        \g[15][40] , \g[15][39] , \g[15][38] , \g[15][37] , \g[15][36] , 
        \g[15][35] , \g[15][34] , \g[15][33] , \g[15][32] , \g[15][31] , 
        \g[15][30] , \g[15][29] , \g[15][28] , \g[15][27] , \g[15][26] , 
        \g[15][25] , \g[15][24] , \g[15][23] , \g[15][22] , \g[15][21] , 
        \g[15][20] , \g[15][19] , \g[15][18] , \g[15][17] , \g[15][16] , 
        \g[15][15] , \g[15][14] , \g[15][13] , \g[15][12] , \g[15][11] , 
        \g[15][10] , \g[15][9] , \g[15][8] , \g[15][7] , \g[15][6] , 
        \g[15][5] , \g[15][4] , \g[15][3] , \g[15][2] , \g[15][1] , \g[15][0] }), .b({\g[16][63] , \g[16][62] , \g[16][61] , \g[16][60] , \g[16][59] , 
        \g[16][58] , \g[16][57] , \g[16][56] , \g[16][55] , \g[16][54] , 
        \g[16][53] , \g[16][52] , \g[16][51] , \g[16][50] , \g[16][49] , 
        \g[16][48] , \g[16][47] , \g[16][46] , \g[16][45] , \g[16][44] , 
        \g[16][43] , \g[16][42] , \g[16][41] , \g[16][40] , \g[16][39] , 
        \g[16][38] , \g[16][37] , \g[16][36] , \g[16][35] , \g[16][34] , 
        \g[16][33] , \g[16][32] , \g[16][31] , \g[16][30] , \g[16][29] , 
        \g[16][28] , \g[16][27] , \g[16][26] , \g[16][25] , \g[16][24] , 
        \g[16][23] , \g[16][22] , \g[16][21] , \g[16][20] , \g[16][19] , 
        \g[16][18] , \g[16][17] , \g[16][16] , \g[16][15] , \g[16][14] , 
        \g[16][13] , \g[16][12] , \g[16][11] , \g[16][10] , \g[16][9] , 
        \g[16][8] , \g[16][7] , \g[16][6] , \g[16][5] , \g[16][4] , \g[16][3] , 
        \g[16][2] , \g[16][1] , \g[16][0] }), .cin({\g[17][63] , \g[17][62] , 
        \g[17][61] , \g[17][60] , \g[17][59] , \g[17][58] , \g[17][57] , 
        \g[17][56] , \g[17][55] , \g[17][54] , \g[17][53] , \g[17][52] , 
        \g[17][51] , \g[17][50] , \g[17][49] , \g[17][48] , \g[17][47] , 
        \g[17][46] , \g[17][45] , \g[17][44] , \g[17][43] , \g[17][42] , 
        \g[17][41] , \g[17][40] , \g[17][39] , \g[17][38] , \g[17][37] , 
        \g[17][36] , \g[17][35] , \g[17][34] , \g[17][33] , \g[17][32] , 
        \g[17][31] , \g[17][30] , \g[17][29] , \g[17][28] , \g[17][27] , 
        \g[17][26] , \g[17][25] , \g[17][24] , \g[17][23] , \g[17][22] , 
        \g[17][21] , \g[17][20] , \g[17][19] , \g[17][18] , \g[17][17] , 
        \g[17][16] , \g[17][15] , \g[17][14] , \g[17][13] , \g[17][12] , 
        \g[17][11] , \g[17][10] , \g[17][9] , \g[17][8] , \g[17][7] , 
        \g[17][6] , \g[17][5] , \g[17][4] , \g[17][3] , \g[17][2] , \g[17][1] , 
        \g[17][0] }), .sum({\g2[5][63] , \g2[5][62] , \g2[5][61] , \g2[5][60] , 
        \g2[5][59] , \g2[5][58] , \g2[5][57] , \g2[5][56] , \g2[5][55] , 
        \g2[5][54] , \g2[5][53] , \g2[5][52] , \g2[5][51] , \g2[5][50] , 
        \g2[5][49] , \g2[5][48] , \g2[5][47] , \g2[5][46] , \g2[5][45] , 
        \g2[5][44] , \g2[5][43] , \g2[5][42] , \g2[5][41] , \g2[5][40] , 
        \g2[5][39] , \g2[5][38] , \g2[5][37] , \g2[5][36] , \g2[5][35] , 
        \g2[5][34] , \g2[5][33] , \g2[5][32] , \g2[5][31] , \g2[5][30] , 
        \g2[5][29] , \g2[5][28] , \g2[5][27] , \g2[5][26] , \g2[5][25] , 
        \g2[5][24] , \g2[5][23] , \g2[5][22] , \g2[5][21] , \g2[5][20] , 
        \g2[5][19] , \g2[5][18] , \g2[5][17] , \g2[5][16] , \g2[5][15] , 
        \g2[5][14] , \g2[5][13] , \g2[5][12] , \g2[5][11] , \g2[5][10] , 
        \g2[5][9] , \g2[5][8] , \g2[5][7] , \g2[5][6] , \g2[5][5] , \g2[5][4] , 
        \g2[5][3] , \g2[5][2] , \g2[5][1] , \g2[5][0] }), .cout({\g2[19][63] , 
        \g2[19][62] , \g2[19][61] , \g2[19][60] , \g2[19][59] , \g2[19][58] , 
        \g2[19][57] , \g2[19][56] , \g2[19][55] , \g2[19][54] , \g2[19][53] , 
        \g2[19][52] , \g2[19][51] , \g2[19][50] , \g2[19][49] , \g2[19][48] , 
        \g2[19][47] , \g2[19][46] , \g2[19][45] , \g2[19][44] , \g2[19][43] , 
        \g2[19][42] , \g2[19][41] , \g2[19][40] , \g2[19][39] , \g2[19][38] , 
        \g2[19][37] , \g2[19][36] , \g2[19][35] , \g2[19][34] , \g2[19][33] , 
        \g2[19][32] , \g2[19][31] , \g2[19][30] , \g2[19][29] , \g2[19][28] , 
        \g2[19][27] , \g2[19][26] , \g2[19][25] , \g2[19][24] , \g2[19][23] , 
        \g2[19][22] , \g2[19][21] , \g2[19][20] , \g2[19][19] , \g2[19][18] , 
        \g2[19][17] , \g2[19][16] , \g2[19][15] , \g2[19][14] , \g2[19][13] , 
        \g2[19][12] , \g2[19][11] , \g2[19][10] , \g2[19][9] , \g2[19][8] , 
        \g2[19][7] , \g2[19][6] , \g2[19][5] , \g2[19][4] , \g2[19][3] , 
        \g2[19][2] , \g2[19][1] , SYNOPSYS_UNCONNECTED__26}) );
  FullAdder \level2[6].x5  ( .a({\g[18][63] , \g[18][62] , \g[18][61] , 
        \g[18][60] , \g[18][59] , \g[18][58] , \g[18][57] , \g[18][56] , 
        \g[18][55] , \g[18][54] , \g[18][53] , \g[18][52] , \g[18][51] , 
        \g[18][50] , \g[18][49] , \g[18][48] , \g[18][47] , \g[18][46] , 
        \g[18][45] , \g[18][44] , \g[18][43] , \g[18][42] , \g[18][41] , 
        \g[18][40] , \g[18][39] , \g[18][38] , \g[18][37] , \g[18][36] , 
        \g[18][35] , \g[18][34] , \g[18][33] , \g[18][32] , \g[18][31] , 
        \g[18][30] , \g[18][29] , \g[18][28] , \g[18][27] , \g[18][26] , 
        \g[18][25] , \g[18][24] , \g[18][23] , \g[18][22] , \g[18][21] , 
        \g[18][20] , \g[18][19] , \g[18][18] , \g[18][17] , \g[18][16] , 
        \g[18][15] , \g[18][14] , \g[18][13] , \g[18][12] , \g[18][11] , 
        \g[18][10] , \g[18][9] , \g[18][8] , \g[18][7] , \g[18][6] , 
        \g[18][5] , \g[18][4] , \g[18][3] , \g[18][2] , \g[18][1] , \g[18][0] }), .b({\g[19][63] , \g[19][62] , \g[19][61] , \g[19][60] , \g[19][59] , 
        \g[19][58] , \g[19][57] , \g[19][56] , \g[19][55] , \g[19][54] , 
        \g[19][53] , \g[19][52] , \g[19][51] , \g[19][50] , \g[19][49] , 
        \g[19][48] , \g[19][47] , \g[19][46] , \g[19][45] , \g[19][44] , 
        \g[19][43] , \g[19][42] , \g[19][41] , \g[19][40] , \g[19][39] , 
        \g[19][38] , \g[19][37] , \g[19][36] , \g[19][35] , \g[19][34] , 
        \g[19][33] , \g[19][32] , \g[19][31] , \g[19][30] , \g[19][29] , 
        \g[19][28] , \g[19][27] , \g[19][26] , \g[19][25] , \g[19][24] , 
        \g[19][23] , \g[19][22] , \g[19][21] , \g[19][20] , \g[19][19] , 
        \g[19][18] , \g[19][17] , \g[19][16] , \g[19][15] , \g[19][14] , 
        \g[19][13] , \g[19][12] , \g[19][11] , \g[19][10] , \g[19][9] , 
        \g[19][8] , \g[19][7] , \g[19][6] , \g[19][5] , \g[19][4] , \g[19][3] , 
        \g[19][2] , \g[19][1] , \g[19][0] }), .cin({\g[20][63] , \g[20][62] , 
        \g[20][61] , \g[20][60] , \g[20][59] , \g[20][58] , \g[20][57] , 
        \g[20][56] , \g[20][55] , \g[20][54] , \g[20][53] , \g[20][52] , 
        \g[20][51] , \g[20][50] , \g[20][49] , \g[20][48] , \g[20][47] , 
        \g[20][46] , \g[20][45] , \g[20][44] , \g[20][43] , \g[20][42] , 
        \g[20][41] , \g[20][40] , \g[20][39] , \g[20][38] , \g[20][37] , 
        \g[20][36] , \g[20][35] , \g[20][34] , \g[20][33] , \g[20][32] , 
        \g[20][31] , \g[20][30] , \g[20][29] , \g[20][28] , \g[20][27] , 
        \g[20][26] , \g[20][25] , \g[20][24] , \g[20][23] , \g[20][22] , 
        \g[20][21] , \g[20][20] , \g[20][19] , \g[20][18] , \g[20][17] , 
        \g[20][16] , \g[20][15] , \g[20][14] , \g[20][13] , \g[20][12] , 
        \g[20][11] , \g[20][10] , \g[20][9] , \g[20][8] , \g[20][7] , 
        \g[20][6] , \g[20][5] , \g[20][4] , \g[20][3] , \g[20][2] , \g[20][1] , 
        \g[20][0] }), .sum({\g2[6][63] , \g2[6][62] , \g2[6][61] , \g2[6][60] , 
        \g2[6][59] , \g2[6][58] , \g2[6][57] , \g2[6][56] , \g2[6][55] , 
        \g2[6][54] , \g2[6][53] , \g2[6][52] , \g2[6][51] , \g2[6][50] , 
        \g2[6][49] , \g2[6][48] , \g2[6][47] , \g2[6][46] , \g2[6][45] , 
        \g2[6][44] , \g2[6][43] , \g2[6][42] , \g2[6][41] , \g2[6][40] , 
        \g2[6][39] , \g2[6][38] , \g2[6][37] , \g2[6][36] , \g2[6][35] , 
        \g2[6][34] , \g2[6][33] , \g2[6][32] , \g2[6][31] , \g2[6][30] , 
        \g2[6][29] , \g2[6][28] , \g2[6][27] , \g2[6][26] , \g2[6][25] , 
        \g2[6][24] , \g2[6][23] , \g2[6][22] , \g2[6][21] , \g2[6][20] , 
        \g2[6][19] , \g2[6][18] , \g2[6][17] , \g2[6][16] , \g2[6][15] , 
        \g2[6][14] , \g2[6][13] , \g2[6][12] , \g2[6][11] , \g2[6][10] , 
        \g2[6][9] , \g2[6][8] , \g2[6][7] , \g2[6][6] , \g2[6][5] , \g2[6][4] , 
        \g2[6][3] , \g2[6][2] , \g2[6][1] , \g2[6][0] }), .cout({\g2[20][63] , 
        \g2[20][62] , \g2[20][61] , \g2[20][60] , \g2[20][59] , \g2[20][58] , 
        \g2[20][57] , \g2[20][56] , \g2[20][55] , \g2[20][54] , \g2[20][53] , 
        \g2[20][52] , \g2[20][51] , \g2[20][50] , \g2[20][49] , \g2[20][48] , 
        \g2[20][47] , \g2[20][46] , \g2[20][45] , \g2[20][44] , \g2[20][43] , 
        \g2[20][42] , \g2[20][41] , \g2[20][40] , \g2[20][39] , \g2[20][38] , 
        \g2[20][37] , \g2[20][36] , \g2[20][35] , \g2[20][34] , \g2[20][33] , 
        \g2[20][32] , \g2[20][31] , \g2[20][30] , \g2[20][29] , \g2[20][28] , 
        \g2[20][27] , \g2[20][26] , \g2[20][25] , \g2[20][24] , \g2[20][23] , 
        \g2[20][22] , \g2[20][21] , \g2[20][20] , \g2[20][19] , \g2[20][18] , 
        \g2[20][17] , \g2[20][16] , \g2[20][15] , \g2[20][14] , \g2[20][13] , 
        \g2[20][12] , \g2[20][11] , \g2[20][10] , \g2[20][9] , \g2[20][8] , 
        \g2[20][7] , \g2[20][6] , \g2[20][5] , \g2[20][4] , \g2[20][3] , 
        \g2[20][2] , \g2[20][1] , SYNOPSYS_UNCONNECTED__27}) );
  FullAdder \level2[7].x5  ( .a({\g[21][63] , \g[21][62] , \g[21][61] , 
        \g[21][60] , \g[21][59] , \g[21][58] , \g[21][57] , \g[21][56] , 
        \g[21][55] , \g[21][54] , \g[21][53] , \g[21][52] , \g[21][51] , 
        \g[21][50] , \g[21][49] , \g[21][48] , \g[21][47] , \g[21][46] , 
        \g[21][45] , \g[21][44] , \g[21][43] , \g[21][42] , \g[21][41] , 
        \g[21][40] , \g[21][39] , \g[21][38] , \g[21][37] , \g[21][36] , 
        \g[21][35] , \g[21][34] , \g[21][33] , \g[21][32] , \g[21][31] , 
        \g[21][30] , \g[21][29] , \g[21][28] , \g[21][27] , \g[21][26] , 
        \g[21][25] , \g[21][24] , \g[21][23] , \g[21][22] , \g[21][21] , 
        \g[21][20] , \g[21][19] , \g[21][18] , \g[21][17] , \g[21][16] , 
        \g[21][15] , \g[21][14] , \g[21][13] , \g[21][12] , \g[21][11] , 
        \g[21][10] , \g[21][9] , \g[21][8] , \g[21][7] , \g[21][6] , 
        \g[21][5] , \g[21][4] , \g[21][3] , \g[21][2] , \g[21][1] , 1'b0}), 
        .b({\g[22][63] , \g[22][62] , \g[22][61] , \g[22][60] , \g[22][59] , 
        \g[22][58] , \g[22][57] , \g[22][56] , \g[22][55] , \g[22][54] , 
        \g[22][53] , \g[22][52] , \g[22][51] , \g[22][50] , \g[22][49] , 
        \g[22][48] , \g[22][47] , \g[22][46] , \g[22][45] , \g[22][44] , 
        \g[22][43] , \g[22][42] , \g[22][41] , \g[22][40] , \g[22][39] , 
        \g[22][38] , \g[22][37] , \g[22][36] , \g[22][35] , \g[22][34] , 
        \g[22][33] , \g[22][32] , \g[22][31] , \g[22][30] , \g[22][29] , 
        \g[22][28] , \g[22][27] , \g[22][26] , \g[22][25] , \g[22][24] , 
        \g[22][23] , \g[22][22] , \g[22][21] , \g[22][20] , \g[22][19] , 
        \g[22][18] , \g[22][17] , \g[22][16] , \g[22][15] , \g[22][14] , 
        \g[22][13] , \g[22][12] , \g[22][11] , \g[22][10] , \g[22][9] , 
        \g[22][8] , \g[22][7] , \g[22][6] , \g[22][5] , \g[22][4] , \g[22][3] , 
        \g[22][2] , \g[22][1] , 1'b0}), .cin({\g[23][63] , \g[23][62] , 
        \g[23][61] , \g[23][60] , \g[23][59] , \g[23][58] , \g[23][57] , 
        \g[23][56] , \g[23][55] , \g[23][54] , \g[23][53] , \g[23][52] , 
        \g[23][51] , \g[23][50] , \g[23][49] , \g[23][48] , \g[23][47] , 
        \g[23][46] , \g[23][45] , \g[23][44] , \g[23][43] , \g[23][42] , 
        \g[23][41] , \g[23][40] , \g[23][39] , \g[23][38] , \g[23][37] , 
        \g[23][36] , \g[23][35] , \g[23][34] , \g[23][33] , \g[23][32] , 
        \g[23][31] , \g[23][30] , \g[23][29] , \g[23][28] , \g[23][27] , 
        \g[23][26] , \g[23][25] , \g[23][24] , \g[23][23] , \g[23][22] , 
        \g[23][21] , \g[23][20] , \g[23][19] , \g[23][18] , \g[23][17] , 
        \g[23][16] , \g[23][15] , \g[23][14] , \g[23][13] , \g[23][12] , 
        \g[23][11] , \g[23][10] , \g[23][9] , \g[23][8] , \g[23][7] , 
        \g[23][6] , \g[23][5] , \g[23][4] , \g[23][3] , \g[23][2] , \g[23][1] , 
        1'b0}), .sum({\g2[7][63] , \g2[7][62] , \g2[7][61] , \g2[7][60] , 
        \g2[7][59] , \g2[7][58] , \g2[7][57] , \g2[7][56] , \g2[7][55] , 
        \g2[7][54] , \g2[7][53] , \g2[7][52] , \g2[7][51] , \g2[7][50] , 
        \g2[7][49] , \g2[7][48] , \g2[7][47] , \g2[7][46] , \g2[7][45] , 
        \g2[7][44] , \g2[7][43] , \g2[7][42] , \g2[7][41] , \g2[7][40] , 
        \g2[7][39] , \g2[7][38] , \g2[7][37] , \g2[7][36] , \g2[7][35] , 
        \g2[7][34] , \g2[7][33] , \g2[7][32] , \g2[7][31] , \g2[7][30] , 
        \g2[7][29] , \g2[7][28] , \g2[7][27] , \g2[7][26] , \g2[7][25] , 
        \g2[7][24] , \g2[7][23] , \g2[7][22] , \g2[7][21] , \g2[7][20] , 
        \g2[7][19] , \g2[7][18] , \g2[7][17] , \g2[7][16] , \g2[7][15] , 
        \g2[7][14] , \g2[7][13] , \g2[7][12] , \g2[7][11] , \g2[7][10] , 
        \g2[7][9] , \g2[7][8] , \g2[7][7] , \g2[7][6] , \g2[7][5] , \g2[7][4] , 
        \g2[7][3] , \g2[7][2] , \g2[7][1] , \g2[7][0] }), .cout({\g2[21][63] , 
        \g2[21][62] , \g2[21][61] , \g2[21][60] , \g2[21][59] , \g2[21][58] , 
        \g2[21][57] , \g2[21][56] , \g2[21][55] , \g2[21][54] , \g2[21][53] , 
        \g2[21][52] , \g2[21][51] , \g2[21][50] , \g2[21][49] , \g2[21][48] , 
        \g2[21][47] , \g2[21][46] , \g2[21][45] , \g2[21][44] , \g2[21][43] , 
        \g2[21][42] , \g2[21][41] , \g2[21][40] , \g2[21][39] , \g2[21][38] , 
        \g2[21][37] , \g2[21][36] , \g2[21][35] , \g2[21][34] , \g2[21][33] , 
        \g2[21][32] , \g2[21][31] , \g2[21][30] , \g2[21][29] , \g2[21][28] , 
        \g2[21][27] , \g2[21][26] , \g2[21][25] , \g2[21][24] , \g2[21][23] , 
        \g2[21][22] , \g2[21][21] , \g2[21][20] , \g2[21][19] , \g2[21][18] , 
        \g2[21][17] , \g2[21][16] , \g2[21][15] , \g2[21][14] , \g2[21][13] , 
        \g2[21][12] , \g2[21][11] , \g2[21][10] , \g2[21][9] , \g2[21][8] , 
        \g2[21][7] , \g2[21][6] , \g2[21][5] , \g2[21][4] , \g2[21][3] , 
        \g2[21][2] , \g2[21][1] , SYNOPSYS_UNCONNECTED__28}) );
  FullAdder \level2[8].x5  ( .a({\g[24][63] , \g[24][62] , \g[24][61] , 
        \g[24][60] , \g[24][59] , \g[24][58] , \g[24][57] , \g[24][56] , 
        \g[24][55] , \g[24][54] , \g[24][53] , \g[24][52] , \g[24][51] , 
        \g[24][50] , \g[24][49] , \g[24][48] , \g[24][47] , \g[24][46] , 
        \g[24][45] , \g[24][44] , \g[24][43] , \g[24][42] , \g[24][41] , 
        \g[24][40] , \g[24][39] , \g[24][38] , \g[24][37] , \g[24][36] , 
        \g[24][35] , \g[24][34] , \g[24][33] , \g[24][32] , \g[24][31] , 
        \g[24][30] , \g[24][29] , \g[24][28] , \g[24][27] , \g[24][26] , 
        \g[24][25] , \g[24][24] , \g[24][23] , \g[24][22] , \g[24][21] , 
        \g[24][20] , \g[24][19] , \g[24][18] , \g[24][17] , \g[24][16] , 
        \g[24][15] , \g[24][14] , \g[24][13] , \g[24][12] , \g[24][11] , 
        \g[24][10] , \g[24][9] , \g[24][8] , \g[24][7] , \g[24][6] , 
        \g[24][5] , \g[24][4] , \g[24][3] , \g[24][2] , \g[24][1] , 1'b0}), 
        .b({\g[25][63] , \g[25][62] , \g[25][61] , \g[25][60] , \g[25][59] , 
        \g[25][58] , \g[25][57] , \g[25][56] , \g[25][55] , \g[25][54] , 
        \g[25][53] , \g[25][52] , \g[25][51] , \g[25][50] , \g[25][49] , 
        \g[25][48] , \g[25][47] , \g[25][46] , \g[25][45] , \g[25][44] , 
        \g[25][43] , \g[25][42] , \g[25][41] , \g[25][40] , \g[25][39] , 
        \g[25][38] , \g[25][37] , \g[25][36] , \g[25][35] , \g[25][34] , 
        \g[25][33] , \g[25][32] , \g[25][31] , \g[25][30] , \g[25][29] , 
        \g[25][28] , \g[25][27] , \g[25][26] , \g[25][25] , \g[25][24] , 
        \g[25][23] , \g[25][22] , \g[25][21] , \g[25][20] , \g[25][19] , 
        \g[25][18] , \g[25][17] , \g[25][16] , \g[25][15] , \g[25][14] , 
        \g[25][13] , \g[25][12] , \g[25][11] , \g[25][10] , \g[25][9] , 
        \g[25][8] , \g[25][7] , \g[25][6] , \g[25][5] , \g[25][4] , \g[25][3] , 
        \g[25][2] , \g[25][1] , 1'b0}), .cin({\g[26][63] , \g[26][62] , 
        \g[26][61] , \g[26][60] , \g[26][59] , \g[26][58] , \g[26][57] , 
        \g[26][56] , \g[26][55] , \g[26][54] , \g[26][53] , \g[26][52] , 
        \g[26][51] , \g[26][50] , \g[26][49] , \g[26][48] , \g[26][47] , 
        \g[26][46] , \g[26][45] , \g[26][44] , \g[26][43] , \g[26][42] , 
        \g[26][41] , \g[26][40] , \g[26][39] , \g[26][38] , \g[26][37] , 
        \g[26][36] , \g[26][35] , \g[26][34] , \g[26][33] , \g[26][32] , 
        \g[26][31] , \g[26][30] , \g[26][29] , \g[26][28] , \g[26][27] , 
        \g[26][26] , \g[26][25] , \g[26][24] , \g[26][23] , \g[26][22] , 
        \g[26][21] , \g[26][20] , \g[26][19] , \g[26][18] , \g[26][17] , 
        \g[26][16] , \g[26][15] , \g[26][14] , \g[26][13] , \g[26][12] , 
        \g[26][11] , \g[26][10] , \g[26][9] , \g[26][8] , \g[26][7] , 
        \g[26][6] , \g[26][5] , \g[26][4] , \g[26][3] , \g[26][2] , \g[26][1] , 
        1'b0}), .sum({\g2[8][63] , \g2[8][62] , \g2[8][61] , \g2[8][60] , 
        \g2[8][59] , \g2[8][58] , \g2[8][57] , \g2[8][56] , \g2[8][55] , 
        \g2[8][54] , \g2[8][53] , \g2[8][52] , \g2[8][51] , \g2[8][50] , 
        \g2[8][49] , \g2[8][48] , \g2[8][47] , \g2[8][46] , \g2[8][45] , 
        \g2[8][44] , \g2[8][43] , \g2[8][42] , \g2[8][41] , \g2[8][40] , 
        \g2[8][39] , \g2[8][38] , \g2[8][37] , \g2[8][36] , \g2[8][35] , 
        \g2[8][34] , \g2[8][33] , \g2[8][32] , \g2[8][31] , \g2[8][30] , 
        \g2[8][29] , \g2[8][28] , \g2[8][27] , \g2[8][26] , \g2[8][25] , 
        \g2[8][24] , \g2[8][23] , \g2[8][22] , \g2[8][21] , \g2[8][20] , 
        \g2[8][19] , \g2[8][18] , \g2[8][17] , \g2[8][16] , \g2[8][15] , 
        \g2[8][14] , \g2[8][13] , \g2[8][12] , \g2[8][11] , \g2[8][10] , 
        \g2[8][9] , \g2[8][8] , \g2[8][7] , \g2[8][6] , \g2[8][5] , \g2[8][4] , 
        \g2[8][3] , \g2[8][2] , \g2[8][1] , \g2[8][0] }), .cout({\g2[22][63] , 
        \g2[22][62] , \g2[22][61] , \g2[22][60] , \g2[22][59] , \g2[22][58] , 
        \g2[22][57] , \g2[22][56] , \g2[22][55] , \g2[22][54] , \g2[22][53] , 
        \g2[22][52] , \g2[22][51] , \g2[22][50] , \g2[22][49] , \g2[22][48] , 
        \g2[22][47] , \g2[22][46] , \g2[22][45] , \g2[22][44] , \g2[22][43] , 
        \g2[22][42] , \g2[22][41] , \g2[22][40] , \g2[22][39] , \g2[22][38] , 
        \g2[22][37] , \g2[22][36] , \g2[22][35] , \g2[22][34] , \g2[22][33] , 
        \g2[22][32] , \g2[22][31] , \g2[22][30] , \g2[22][29] , \g2[22][28] , 
        \g2[22][27] , \g2[22][26] , \g2[22][25] , \g2[22][24] , \g2[22][23] , 
        \g2[22][22] , \g2[22][21] , \g2[22][20] , \g2[22][19] , \g2[22][18] , 
        \g2[22][17] , \g2[22][16] , \g2[22][15] , \g2[22][14] , \g2[22][13] , 
        \g2[22][12] , \g2[22][11] , \g2[22][10] , \g2[22][9] , \g2[22][8] , 
        \g2[22][7] , \g2[22][6] , \g2[22][5] , \g2[22][4] , \g2[22][3] , 
        \g2[22][2] , \g2[22][1] , SYNOPSYS_UNCONNECTED__29}) );
  FullAdder \level2[9].x5  ( .a({\g[27][63] , \g[27][62] , \g[27][61] , 
        \g[27][60] , \g[27][59] , \g[27][58] , \g[27][57] , \g[27][56] , 
        \g[27][55] , \g[27][54] , \g[27][53] , \g[27][52] , \g[27][51] , 
        \g[27][50] , \g[27][49] , \g[27][48] , \g[27][47] , \g[27][46] , 
        \g[27][45] , \g[27][44] , \g[27][43] , \g[27][42] , \g[27][41] , 
        \g[27][40] , \g[27][39] , \g[27][38] , \g[27][37] , \g[27][36] , 
        \g[27][35] , \g[27][34] , \g[27][33] , \g[27][32] , \g[27][31] , 
        \g[27][30] , \g[27][29] , \g[27][28] , \g[27][27] , \g[27][26] , 
        \g[27][25] , \g[27][24] , \g[27][23] , \g[27][22] , \g[27][21] , 
        \g[27][20] , \g[27][19] , \g[27][18] , \g[27][17] , \g[27][16] , 
        \g[27][15] , \g[27][14] , \g[27][13] , \g[27][12] , \g[27][11] , 
        \g[27][10] , \g[27][9] , \g[27][8] , \g[27][7] , \g[27][6] , 
        \g[27][5] , \g[27][4] , \g[27][3] , \g[27][2] , \g[27][1] , 1'b0}), 
        .b({\g[28][63] , \g[28][62] , \g[28][61] , \g[28][60] , \g[28][59] , 
        \g[28][58] , \g[28][57] , \g[28][56] , \g[28][55] , \g[28][54] , 
        \g[28][53] , \g[28][52] , \g[28][51] , \g[28][50] , \g[28][49] , 
        \g[28][48] , \g[28][47] , \g[28][46] , \g[28][45] , \g[28][44] , 
        \g[28][43] , \g[28][42] , \g[28][41] , \g[28][40] , \g[28][39] , 
        \g[28][38] , \g[28][37] , \g[28][36] , \g[28][35] , \g[28][34] , 
        \g[28][33] , \g[28][32] , \g[28][31] , \g[28][30] , \g[28][29] , 
        \g[28][28] , \g[28][27] , \g[28][26] , \g[28][25] , \g[28][24] , 
        \g[28][23] , \g[28][22] , \g[28][21] , \g[28][20] , \g[28][19] , 
        \g[28][18] , \g[28][17] , \g[28][16] , \g[28][15] , \g[28][14] , 
        \g[28][13] , \g[28][12] , \g[28][11] , \g[28][10] , \g[28][9] , 
        \g[28][8] , \g[28][7] , \g[28][6] , \g[28][5] , \g[28][4] , \g[28][3] , 
        \g[28][2] , \g[28][1] , 1'b0}), .cin({\g[29][63] , \g[29][62] , 
        \g[29][61] , \g[29][60] , \g[29][59] , \g[29][58] , \g[29][57] , 
        \g[29][56] , \g[29][55] , \g[29][54] , \g[29][53] , \g[29][52] , 
        \g[29][51] , \g[29][50] , \g[29][49] , \g[29][48] , \g[29][47] , 
        \g[29][46] , \g[29][45] , \g[29][44] , \g[29][43] , \g[29][42] , 
        \g[29][41] , \g[29][40] , \g[29][39] , \g[29][38] , \g[29][37] , 
        \g[29][36] , \g[29][35] , \g[29][34] , \g[29][33] , \g[29][32] , 
        \g[29][31] , \g[29][30] , \g[29][29] , \g[29][28] , \g[29][27] , 
        \g[29][26] , \g[29][25] , \g[29][24] , \g[29][23] , \g[29][22] , 
        \g[29][21] , \g[29][20] , \g[29][19] , \g[29][18] , \g[29][17] , 
        \g[29][16] , \g[29][15] , \g[29][14] , \g[29][13] , \g[29][12] , 
        \g[29][11] , \g[29][10] , \g[29][9] , \g[29][8] , \g[29][7] , 
        \g[29][6] , \g[29][5] , \g[29][4] , \g[29][3] , \g[29][2] , \g[29][1] , 
        1'b0}), .sum({\g2[9][63] , \g2[9][62] , \g2[9][61] , \g2[9][60] , 
        \g2[9][59] , \g2[9][58] , \g2[9][57] , \g2[9][56] , \g2[9][55] , 
        \g2[9][54] , \g2[9][53] , \g2[9][52] , \g2[9][51] , \g2[9][50] , 
        \g2[9][49] , \g2[9][48] , \g2[9][47] , \g2[9][46] , \g2[9][45] , 
        \g2[9][44] , \g2[9][43] , \g2[9][42] , \g2[9][41] , \g2[9][40] , 
        \g2[9][39] , \g2[9][38] , \g2[9][37] , \g2[9][36] , \g2[9][35] , 
        \g2[9][34] , \g2[9][33] , \g2[9][32] , \g2[9][31] , \g2[9][30] , 
        \g2[9][29] , \g2[9][28] , \g2[9][27] , \g2[9][26] , \g2[9][25] , 
        \g2[9][24] , \g2[9][23] , \g2[9][22] , \g2[9][21] , \g2[9][20] , 
        \g2[9][19] , \g2[9][18] , \g2[9][17] , \g2[9][16] , \g2[9][15] , 
        \g2[9][14] , \g2[9][13] , \g2[9][12] , \g2[9][11] , \g2[9][10] , 
        \g2[9][9] , \g2[9][8] , \g2[9][7] , \g2[9][6] , \g2[9][5] , \g2[9][4] , 
        \g2[9][3] , \g2[9][2] , \g2[9][1] , \g2[9][0] }), .cout({\g2[23][63] , 
        \g2[23][62] , \g2[23][61] , \g2[23][60] , \g2[23][59] , \g2[23][58] , 
        \g2[23][57] , \g2[23][56] , \g2[23][55] , \g2[23][54] , \g2[23][53] , 
        \g2[23][52] , \g2[23][51] , \g2[23][50] , \g2[23][49] , \g2[23][48] , 
        \g2[23][47] , \g2[23][46] , \g2[23][45] , \g2[23][44] , \g2[23][43] , 
        \g2[23][42] , \g2[23][41] , \g2[23][40] , \g2[23][39] , \g2[23][38] , 
        \g2[23][37] , \g2[23][36] , \g2[23][35] , \g2[23][34] , \g2[23][33] , 
        \g2[23][32] , \g2[23][31] , \g2[23][30] , \g2[23][29] , \g2[23][28] , 
        \g2[23][27] , \g2[23][26] , \g2[23][25] , \g2[23][24] , \g2[23][23] , 
        \g2[23][22] , \g2[23][21] , \g2[23][20] , \g2[23][19] , \g2[23][18] , 
        \g2[23][17] , \g2[23][16] , \g2[23][15] , \g2[23][14] , \g2[23][13] , 
        \g2[23][12] , \g2[23][11] , \g2[23][10] , \g2[23][9] , \g2[23][8] , 
        \g2[23][7] , \g2[23][6] , \g2[23][5] , \g2[23][4] , \g2[23][3] , 
        \g2[23][2] , \g2[23][1] , SYNOPSYS_UNCONNECTED__30}) );
  FullAdder \level2[10].x5  ( .a({\g[30][63] , \g[30][62] , \g[30][61] , 
        \g[30][60] , \g[30][59] , \g[30][58] , \g[30][57] , \g[30][56] , 
        \g[30][55] , \g[30][54] , \g[30][53] , \g[30][52] , \g[30][51] , 
        \g[30][50] , \g[30][49] , \g[30][48] , \g[30][47] , \g[30][46] , 
        \g[30][45] , \g[30][44] , \g[30][43] , \g[30][42] , \g[30][41] , 
        \g[30][40] , \g[30][39] , \g[30][38] , \g[30][37] , \g[30][36] , 
        \g[30][35] , \g[30][34] , \g[30][33] , \g[30][32] , \g[30][31] , 
        \g[30][30] , \g[30][29] , \g[30][28] , \g[30][27] , \g[30][26] , 
        \g[30][25] , \g[30][24] , \g[30][23] , \g[30][22] , \g[30][21] , 
        \g[30][20] , \g[30][19] , \g[30][18] , \g[30][17] , \g[30][16] , 
        \g[30][15] , \g[30][14] , \g[30][13] , \g[30][12] , \g[30][11] , 
        \g[30][10] , \g[30][9] , \g[30][8] , \g[30][7] , \g[30][6] , 
        \g[30][5] , \g[30][4] , \g[30][3] , \g[30][2] , \g[30][1] , 1'b0}), 
        .b({\g[31][63] , \g[31][62] , \g[31][61] , \g[31][60] , \g[31][59] , 
        \g[31][58] , \g[31][57] , \g[31][56] , \g[31][55] , \g[31][54] , 
        \g[31][53] , \g[31][52] , \g[31][51] , \g[31][50] , \g[31][49] , 
        \g[31][48] , \g[31][47] , \g[31][46] , \g[31][45] , \g[31][44] , 
        \g[31][43] , \g[31][42] , \g[31][41] , \g[31][40] , \g[31][39] , 
        \g[31][38] , \g[31][37] , \g[31][36] , \g[31][35] , \g[31][34] , 
        \g[31][33] , \g[31][32] , \g[31][31] , \g[31][30] , \g[31][29] , 
        \g[31][28] , \g[31][27] , \g[31][26] , \g[31][25] , \g[31][24] , 
        \g[31][23] , \g[31][22] , \g[31][21] , \g[31][20] , \g[31][19] , 
        \g[31][18] , \g[31][17] , \g[31][16] , \g[31][15] , \g[31][14] , 
        \g[31][13] , \g[31][12] , \g[31][11] , \g[31][10] , \g[31][9] , 
        \g[31][8] , \g[31][7] , \g[31][6] , \g[31][5] , \g[31][4] , \g[31][3] , 
        \g[31][2] , \g[31][1] , 1'b0}), .cin({\g[32][63] , \g[32][62] , 
        \g[32][61] , \g[32][60] , \g[32][59] , \g[32][58] , \g[32][57] , 
        \g[32][56] , \g[32][55] , \g[32][54] , \g[32][53] , \g[32][52] , 
        \g[32][51] , \g[32][50] , \g[32][49] , \g[32][48] , \g[32][47] , 
        \g[32][46] , \g[32][45] , \g[32][44] , \g[32][43] , \g[32][42] , 
        \g[32][41] , \g[32][40] , \g[32][39] , \g[32][38] , \g[32][37] , 
        \g[32][36] , \g[32][35] , \g[32][34] , \g[32][33] , \g[32][32] , 
        \g[32][31] , \g[32][30] , \g[32][29] , \g[32][28] , \g[32][27] , 
        \g[32][26] , \g[32][25] , \g[32][24] , \g[32][23] , \g[32][22] , 
        \g[32][21] , \g[32][20] , \g[32][19] , \g[32][18] , \g[32][17] , 
        \g[32][16] , \g[32][15] , \g[32][14] , \g[32][13] , \g[32][12] , 
        \g[32][11] , \g[32][10] , \g[32][9] , \g[32][8] , \g[32][7] , 
        \g[32][6] , \g[32][5] , \g[32][4] , \g[32][3] , \g[32][2] , \g[32][1] , 
        1'b0}), .sum({\g2[10][63] , \g2[10][62] , \g2[10][61] , \g2[10][60] , 
        \g2[10][59] , \g2[10][58] , \g2[10][57] , \g2[10][56] , \g2[10][55] , 
        \g2[10][54] , \g2[10][53] , \g2[10][52] , \g2[10][51] , \g2[10][50] , 
        \g2[10][49] , \g2[10][48] , \g2[10][47] , \g2[10][46] , \g2[10][45] , 
        \g2[10][44] , \g2[10][43] , \g2[10][42] , \g2[10][41] , \g2[10][40] , 
        \g2[10][39] , \g2[10][38] , \g2[10][37] , \g2[10][36] , \g2[10][35] , 
        \g2[10][34] , \g2[10][33] , \g2[10][32] , \g2[10][31] , \g2[10][30] , 
        \g2[10][29] , \g2[10][28] , \g2[10][27] , \g2[10][26] , \g2[10][25] , 
        \g2[10][24] , \g2[10][23] , \g2[10][22] , \g2[10][21] , \g2[10][20] , 
        \g2[10][19] , \g2[10][18] , \g2[10][17] , \g2[10][16] , \g2[10][15] , 
        \g2[10][14] , \g2[10][13] , \g2[10][12] , \g2[10][11] , \g2[10][10] , 
        \g2[10][9] , \g2[10][8] , \g2[10][7] , \g2[10][6] , \g2[10][5] , 
        \g2[10][4] , \g2[10][3] , \g2[10][2] , \g2[10][1] , \g2[10][0] }), 
        .cout({\g2[24][63] , \g2[24][62] , \g2[24][61] , \g2[24][60] , 
        \g2[24][59] , \g2[24][58] , \g2[24][57] , \g2[24][56] , \g2[24][55] , 
        \g2[24][54] , \g2[24][53] , \g2[24][52] , \g2[24][51] , \g2[24][50] , 
        \g2[24][49] , \g2[24][48] , \g2[24][47] , \g2[24][46] , \g2[24][45] , 
        \g2[24][44] , \g2[24][43] , \g2[24][42] , \g2[24][41] , \g2[24][40] , 
        \g2[24][39] , \g2[24][38] , \g2[24][37] , \g2[24][36] , \g2[24][35] , 
        \g2[24][34] , \g2[24][33] , \g2[24][32] , \g2[24][31] , \g2[24][30] , 
        \g2[24][29] , \g2[24][28] , \g2[24][27] , \g2[24][26] , \g2[24][25] , 
        \g2[24][24] , \g2[24][23] , \g2[24][22] , \g2[24][21] , \g2[24][20] , 
        \g2[24][19] , \g2[24][18] , \g2[24][17] , \g2[24][16] , \g2[24][15] , 
        \g2[24][14] , \g2[24][13] , \g2[24][12] , \g2[24][11] , \g2[24][10] , 
        \g2[24][9] , \g2[24][8] , \g2[24][7] , \g2[24][6] , \g2[24][5] , 
        \g2[24][4] , \g2[24][3] , \g2[24][2] , \g2[24][1] , 
        SYNOPSYS_UNCONNECTED__31}) );
  FullAdder \level2[11].x5  ( .a({\g[33][63] , \g[33][62] , \g[33][61] , 
        \g[33][60] , \g[33][59] , \g[33][58] , \g[33][57] , \g[33][56] , 
        \g[33][55] , \g[33][54] , \g[33][53] , \g[33][52] , \g[33][51] , 
        \g[33][50] , \g[33][49] , \g[33][48] , \g[33][47] , \g[33][46] , 
        \g[33][45] , \g[33][44] , \g[33][43] , \g[33][42] , \g[33][41] , 
        \g[33][40] , \g[33][39] , \g[33][38] , \g[33][37] , \g[33][36] , 
        \g[33][35] , \g[33][34] , \g[33][33] , \g[33][32] , \g[33][31] , 
        \g[33][30] , \g[33][29] , \g[33][28] , \g[33][27] , \g[33][26] , 
        \g[33][25] , \g[33][24] , \g[33][23] , \g[33][22] , \g[33][21] , 
        \g[33][20] , \g[33][19] , \g[33][18] , \g[33][17] , \g[33][16] , 
        \g[33][15] , \g[33][14] , \g[33][13] , \g[33][12] , \g[33][11] , 
        \g[33][10] , \g[33][9] , \g[33][8] , \g[33][7] , \g[33][6] , 
        \g[33][5] , \g[33][4] , \g[33][3] , \g[33][2] , \g[33][1] , 1'b0}), 
        .b({\g[34][63] , \g[34][62] , \g[34][61] , \g[34][60] , \g[34][59] , 
        \g[34][58] , \g[34][57] , \g[34][56] , \g[34][55] , \g[34][54] , 
        \g[34][53] , \g[34][52] , \g[34][51] , \g[34][50] , \g[34][49] , 
        \g[34][48] , \g[34][47] , \g[34][46] , \g[34][45] , \g[34][44] , 
        \g[34][43] , \g[34][42] , \g[34][41] , \g[34][40] , \g[34][39] , 
        \g[34][38] , \g[34][37] , \g[34][36] , \g[34][35] , \g[34][34] , 
        \g[34][33] , \g[34][32] , \g[34][31] , \g[34][30] , \g[34][29] , 
        \g[34][28] , \g[34][27] , \g[34][26] , \g[34][25] , \g[34][24] , 
        \g[34][23] , \g[34][22] , \g[34][21] , \g[34][20] , \g[34][19] , 
        \g[34][18] , \g[34][17] , \g[34][16] , \g[34][15] , \g[34][14] , 
        \g[34][13] , \g[34][12] , \g[34][11] , \g[34][10] , \g[34][9] , 
        \g[34][8] , \g[34][7] , \g[34][6] , \g[34][5] , \g[34][4] , \g[34][3] , 
        \g[34][2] , \g[34][1] , 1'b0}), .cin({\g[35][63] , \g[35][62] , 
        \g[35][61] , \g[35][60] , \g[35][59] , \g[35][58] , \g[35][57] , 
        \g[35][56] , \g[35][55] , \g[35][54] , \g[35][53] , \g[35][52] , 
        \g[35][51] , \g[35][50] , \g[35][49] , \g[35][48] , \g[35][47] , 
        \g[35][46] , \g[35][45] , \g[35][44] , \g[35][43] , \g[35][42] , 
        \g[35][41] , \g[35][40] , \g[35][39] , \g[35][38] , \g[35][37] , 
        \g[35][36] , \g[35][35] , \g[35][34] , \g[35][33] , \g[35][32] , 
        \g[35][31] , \g[35][30] , \g[35][29] , \g[35][28] , \g[35][27] , 
        \g[35][26] , \g[35][25] , \g[35][24] , \g[35][23] , \g[35][22] , 
        \g[35][21] , \g[35][20] , \g[35][19] , \g[35][18] , \g[35][17] , 
        \g[35][16] , \g[35][15] , \g[35][14] , \g[35][13] , \g[35][12] , 
        \g[35][11] , \g[35][10] , \g[35][9] , \g[35][8] , \g[35][7] , 
        \g[35][6] , \g[35][5] , \g[35][4] , \g[35][3] , \g[35][2] , \g[35][1] , 
        1'b0}), .sum({\g2[11][63] , \g2[11][62] , \g2[11][61] , \g2[11][60] , 
        \g2[11][59] , \g2[11][58] , \g2[11][57] , \g2[11][56] , \g2[11][55] , 
        \g2[11][54] , \g2[11][53] , \g2[11][52] , \g2[11][51] , \g2[11][50] , 
        \g2[11][49] , \g2[11][48] , \g2[11][47] , \g2[11][46] , \g2[11][45] , 
        \g2[11][44] , \g2[11][43] , \g2[11][42] , \g2[11][41] , \g2[11][40] , 
        \g2[11][39] , \g2[11][38] , \g2[11][37] , \g2[11][36] , \g2[11][35] , 
        \g2[11][34] , \g2[11][33] , \g2[11][32] , \g2[11][31] , \g2[11][30] , 
        \g2[11][29] , \g2[11][28] , \g2[11][27] , \g2[11][26] , \g2[11][25] , 
        \g2[11][24] , \g2[11][23] , \g2[11][22] , \g2[11][21] , \g2[11][20] , 
        \g2[11][19] , \g2[11][18] , \g2[11][17] , \g2[11][16] , \g2[11][15] , 
        \g2[11][14] , \g2[11][13] , \g2[11][12] , \g2[11][11] , \g2[11][10] , 
        \g2[11][9] , \g2[11][8] , \g2[11][7] , \g2[11][6] , \g2[11][5] , 
        \g2[11][4] , \g2[11][3] , \g2[11][2] , \g2[11][1] , \g2[11][0] }), 
        .cout({\g2[25][63] , \g2[25][62] , \g2[25][61] , \g2[25][60] , 
        \g2[25][59] , \g2[25][58] , \g2[25][57] , \g2[25][56] , \g2[25][55] , 
        \g2[25][54] , \g2[25][53] , \g2[25][52] , \g2[25][51] , \g2[25][50] , 
        \g2[25][49] , \g2[25][48] , \g2[25][47] , \g2[25][46] , \g2[25][45] , 
        \g2[25][44] , \g2[25][43] , \g2[25][42] , \g2[25][41] , \g2[25][40] , 
        \g2[25][39] , \g2[25][38] , \g2[25][37] , \g2[25][36] , \g2[25][35] , 
        \g2[25][34] , \g2[25][33] , \g2[25][32] , \g2[25][31] , \g2[25][30] , 
        \g2[25][29] , \g2[25][28] , \g2[25][27] , \g2[25][26] , \g2[25][25] , 
        \g2[25][24] , \g2[25][23] , \g2[25][22] , \g2[25][21] , \g2[25][20] , 
        \g2[25][19] , \g2[25][18] , \g2[25][17] , \g2[25][16] , \g2[25][15] , 
        \g2[25][14] , \g2[25][13] , \g2[25][12] , \g2[25][11] , \g2[25][10] , 
        \g2[25][9] , \g2[25][8] , \g2[25][7] , \g2[25][6] , \g2[25][5] , 
        \g2[25][4] , \g2[25][3] , \g2[25][2] , \g2[25][1] , 
        SYNOPSYS_UNCONNECTED__32}) );
  FullAdder \level2[12].x5  ( .a({\g[36][63] , \g[36][62] , \g[36][61] , 
        \g[36][60] , \g[36][59] , \g[36][58] , \g[36][57] , \g[36][56] , 
        \g[36][55] , \g[36][54] , \g[36][53] , \g[36][52] , \g[36][51] , 
        \g[36][50] , \g[36][49] , \g[36][48] , \g[36][47] , \g[36][46] , 
        \g[36][45] , \g[36][44] , \g[36][43] , \g[36][42] , \g[36][41] , 
        \g[36][40] , \g[36][39] , \g[36][38] , \g[36][37] , \g[36][36] , 
        \g[36][35] , \g[36][34] , \g[36][33] , \g[36][32] , \g[36][31] , 
        \g[36][30] , \g[36][29] , \g[36][28] , \g[36][27] , \g[36][26] , 
        \g[36][25] , \g[36][24] , \g[36][23] , \g[36][22] , \g[36][21] , 
        \g[36][20] , \g[36][19] , \g[36][18] , \g[36][17] , \g[36][16] , 
        \g[36][15] , \g[36][14] , \g[36][13] , \g[36][12] , \g[36][11] , 
        \g[36][10] , \g[36][9] , \g[36][8] , \g[36][7] , \g[36][6] , 
        \g[36][5] , \g[36][4] , \g[36][3] , \g[36][2] , \g[36][1] , 1'b0}), 
        .b({\g[37][63] , \g[37][62] , \g[37][61] , \g[37][60] , \g[37][59] , 
        \g[37][58] , \g[37][57] , \g[37][56] , \g[37][55] , \g[37][54] , 
        \g[37][53] , \g[37][52] , \g[37][51] , \g[37][50] , \g[37][49] , 
        \g[37][48] , \g[37][47] , \g[37][46] , \g[37][45] , \g[37][44] , 
        \g[37][43] , \g[37][42] , \g[37][41] , \g[37][40] , \g[37][39] , 
        \g[37][38] , \g[37][37] , \g[37][36] , \g[37][35] , \g[37][34] , 
        \g[37][33] , \g[37][32] , \g[37][31] , \g[37][30] , \g[37][29] , 
        \g[37][28] , \g[37][27] , \g[37][26] , \g[37][25] , \g[37][24] , 
        \g[37][23] , \g[37][22] , \g[37][21] , \g[37][20] , \g[37][19] , 
        \g[37][18] , \g[37][17] , \g[37][16] , \g[37][15] , \g[37][14] , 
        \g[37][13] , \g[37][12] , \g[37][11] , \g[37][10] , \g[37][9] , 
        \g[37][8] , \g[37][7] , \g[37][6] , \g[37][5] , \g[37][4] , \g[37][3] , 
        \g[37][2] , \g[37][1] , 1'b0}), .cin({\g[38][63] , \g[38][62] , 
        \g[38][61] , \g[38][60] , \g[38][59] , \g[38][58] , \g[38][57] , 
        \g[38][56] , \g[38][55] , \g[38][54] , \g[38][53] , \g[38][52] , 
        \g[38][51] , \g[38][50] , \g[38][49] , \g[38][48] , \g[38][47] , 
        \g[38][46] , \g[38][45] , \g[38][44] , \g[38][43] , \g[38][42] , 
        \g[38][41] , \g[38][40] , \g[38][39] , \g[38][38] , \g[38][37] , 
        \g[38][36] , \g[38][35] , \g[38][34] , \g[38][33] , \g[38][32] , 
        \g[38][31] , \g[38][30] , \g[38][29] , \g[38][28] , \g[38][27] , 
        \g[38][26] , \g[38][25] , \g[38][24] , \g[38][23] , \g[38][22] , 
        \g[38][21] , \g[38][20] , \g[38][19] , \g[38][18] , \g[38][17] , 
        \g[38][16] , \g[38][15] , \g[38][14] , \g[38][13] , \g[38][12] , 
        \g[38][11] , \g[38][10] , \g[38][9] , \g[38][8] , \g[38][7] , 
        \g[38][6] , \g[38][5] , \g[38][4] , \g[38][3] , \g[38][2] , \g[38][1] , 
        1'b0}), .sum({\g2[12][63] , \g2[12][62] , \g2[12][61] , \g2[12][60] , 
        \g2[12][59] , \g2[12][58] , \g2[12][57] , \g2[12][56] , \g2[12][55] , 
        \g2[12][54] , \g2[12][53] , \g2[12][52] , \g2[12][51] , \g2[12][50] , 
        \g2[12][49] , \g2[12][48] , \g2[12][47] , \g2[12][46] , \g2[12][45] , 
        \g2[12][44] , \g2[12][43] , \g2[12][42] , \g2[12][41] , \g2[12][40] , 
        \g2[12][39] , \g2[12][38] , \g2[12][37] , \g2[12][36] , \g2[12][35] , 
        \g2[12][34] , \g2[12][33] , \g2[12][32] , \g2[12][31] , \g2[12][30] , 
        \g2[12][29] , \g2[12][28] , \g2[12][27] , \g2[12][26] , \g2[12][25] , 
        \g2[12][24] , \g2[12][23] , \g2[12][22] , \g2[12][21] , \g2[12][20] , 
        \g2[12][19] , \g2[12][18] , \g2[12][17] , \g2[12][16] , \g2[12][15] , 
        \g2[12][14] , \g2[12][13] , \g2[12][12] , \g2[12][11] , \g2[12][10] , 
        \g2[12][9] , \g2[12][8] , \g2[12][7] , \g2[12][6] , \g2[12][5] , 
        \g2[12][4] , \g2[12][3] , \g2[12][2] , \g2[12][1] , \g2[12][0] }), 
        .cout({\g2[26][63] , \g2[26][62] , \g2[26][61] , \g2[26][60] , 
        \g2[26][59] , \g2[26][58] , \g2[26][57] , \g2[26][56] , \g2[26][55] , 
        \g2[26][54] , \g2[26][53] , \g2[26][52] , \g2[26][51] , \g2[26][50] , 
        \g2[26][49] , \g2[26][48] , \g2[26][47] , \g2[26][46] , \g2[26][45] , 
        \g2[26][44] , \g2[26][43] , \g2[26][42] , \g2[26][41] , \g2[26][40] , 
        \g2[26][39] , \g2[26][38] , \g2[26][37] , \g2[26][36] , \g2[26][35] , 
        \g2[26][34] , \g2[26][33] , \g2[26][32] , \g2[26][31] , \g2[26][30] , 
        \g2[26][29] , \g2[26][28] , \g2[26][27] , \g2[26][26] , \g2[26][25] , 
        \g2[26][24] , \g2[26][23] , \g2[26][22] , \g2[26][21] , \g2[26][20] , 
        \g2[26][19] , \g2[26][18] , \g2[26][17] , \g2[26][16] , \g2[26][15] , 
        \g2[26][14] , \g2[26][13] , \g2[26][12] , \g2[26][11] , \g2[26][10] , 
        \g2[26][9] , \g2[26][8] , \g2[26][7] , \g2[26][6] , \g2[26][5] , 
        \g2[26][4] , \g2[26][3] , \g2[26][2] , \g2[26][1] , 
        SYNOPSYS_UNCONNECTED__33}) );
  FullAdder \level2[13].x5  ( .a({\g[39][63] , \g[39][62] , \g[39][61] , 
        \g[39][60] , \g[39][59] , \g[39][58] , \g[39][57] , \g[39][56] , 
        \g[39][55] , \g[39][54] , \g[39][53] , \g[39][52] , \g[39][51] , 
        \g[39][50] , \g[39][49] , \g[39][48] , \g[39][47] , \g[39][46] , 
        \g[39][45] , \g[39][44] , \g[39][43] , \g[39][42] , \g[39][41] , 
        \g[39][40] , \g[39][39] , \g[39][38] , \g[39][37] , \g[39][36] , 
        \g[39][35] , \g[39][34] , \g[39][33] , \g[39][32] , \g[39][31] , 
        \g[39][30] , \g[39][29] , \g[39][28] , \g[39][27] , \g[39][26] , 
        \g[39][25] , \g[39][24] , \g[39][23] , \g[39][22] , \g[39][21] , 
        \g[39][20] , \g[39][19] , \g[39][18] , \g[39][17] , \g[39][16] , 
        \g[39][15] , \g[39][14] , \g[39][13] , \g[39][12] , \g[39][11] , 
        \g[39][10] , \g[39][9] , \g[39][8] , \g[39][7] , \g[39][6] , 
        \g[39][5] , \g[39][4] , \g[39][3] , \g[39][2] , \g[39][1] , 1'b0}), 
        .b({\g[40][63] , \g[40][62] , \g[40][61] , \g[40][60] , \g[40][59] , 
        \g[40][58] , \g[40][57] , \g[40][56] , \g[40][55] , \g[40][54] , 
        \g[40][53] , \g[40][52] , \g[40][51] , \g[40][50] , \g[40][49] , 
        \g[40][48] , \g[40][47] , \g[40][46] , \g[40][45] , \g[40][44] , 
        \g[40][43] , \g[40][42] , \g[40][41] , \g[40][40] , \g[40][39] , 
        \g[40][38] , \g[40][37] , \g[40][36] , \g[40][35] , \g[40][34] , 
        \g[40][33] , \g[40][32] , \g[40][31] , \g[40][30] , \g[40][29] , 
        \g[40][28] , \g[40][27] , \g[40][26] , \g[40][25] , \g[40][24] , 
        \g[40][23] , \g[40][22] , \g[40][21] , \g[40][20] , \g[40][19] , 
        \g[40][18] , \g[40][17] , \g[40][16] , \g[40][15] , \g[40][14] , 
        \g[40][13] , \g[40][12] , \g[40][11] , \g[40][10] , \g[40][9] , 
        \g[40][8] , \g[40][7] , \g[40][6] , \g[40][5] , \g[40][4] , \g[40][3] , 
        \g[40][2] , \g[40][1] , 1'b0}), .cin({\g[41][63] , \g[41][62] , 
        \g[41][61] , \g[41][60] , \g[41][59] , \g[41][58] , \g[41][57] , 
        \g[41][56] , \g[41][55] , \g[41][54] , \g[41][53] , \g[41][52] , 
        \g[41][51] , \g[41][50] , \g[41][49] , \g[41][48] , \g[41][47] , 
        \g[41][46] , \g[41][45] , \g[41][44] , \g[41][43] , \g[41][42] , 
        \g[41][41] , \g[41][40] , \g[41][39] , \g[41][38] , \g[41][37] , 
        \g[41][36] , \g[41][35] , \g[41][34] , \g[41][33] , \g[41][32] , 
        \g[41][31] , \g[41][30] , \g[41][29] , \g[41][28] , \g[41][27] , 
        \g[41][26] , \g[41][25] , \g[41][24] , \g[41][23] , \g[41][22] , 
        \g[41][21] , \g[41][20] , \g[41][19] , \g[41][18] , \g[41][17] , 
        \g[41][16] , \g[41][15] , \g[41][14] , \g[41][13] , \g[41][12] , 
        \g[41][11] , \g[41][10] , \g[41][9] , \g[41][8] , \g[41][7] , 
        \g[41][6] , \g[41][5] , \g[41][4] , \g[41][3] , \g[41][2] , \g[41][1] , 
        1'b0}), .sum({\g2[13][63] , \g2[13][62] , \g2[13][61] , \g2[13][60] , 
        \g2[13][59] , \g2[13][58] , \g2[13][57] , \g2[13][56] , \g2[13][55] , 
        \g2[13][54] , \g2[13][53] , \g2[13][52] , \g2[13][51] , \g2[13][50] , 
        \g2[13][49] , \g2[13][48] , \g2[13][47] , \g2[13][46] , \g2[13][45] , 
        \g2[13][44] , \g2[13][43] , \g2[13][42] , \g2[13][41] , \g2[13][40] , 
        \g2[13][39] , \g2[13][38] , \g2[13][37] , \g2[13][36] , \g2[13][35] , 
        \g2[13][34] , \g2[13][33] , \g2[13][32] , \g2[13][31] , \g2[13][30] , 
        \g2[13][29] , \g2[13][28] , \g2[13][27] , \g2[13][26] , \g2[13][25] , 
        \g2[13][24] , \g2[13][23] , \g2[13][22] , \g2[13][21] , \g2[13][20] , 
        \g2[13][19] , \g2[13][18] , \g2[13][17] , \g2[13][16] , \g2[13][15] , 
        \g2[13][14] , \g2[13][13] , \g2[13][12] , \g2[13][11] , \g2[13][10] , 
        \g2[13][9] , \g2[13][8] , \g2[13][7] , \g2[13][6] , \g2[13][5] , 
        \g2[13][4] , \g2[13][3] , \g2[13][2] , \g2[13][1] , \g2[13][0] }), 
        .cout({\g2[27][63] , \g2[27][62] , \g2[27][61] , \g2[27][60] , 
        \g2[27][59] , \g2[27][58] , \g2[27][57] , \g2[27][56] , \g2[27][55] , 
        \g2[27][54] , \g2[27][53] , \g2[27][52] , \g2[27][51] , \g2[27][50] , 
        \g2[27][49] , \g2[27][48] , \g2[27][47] , \g2[27][46] , \g2[27][45] , 
        \g2[27][44] , \g2[27][43] , \g2[27][42] , \g2[27][41] , \g2[27][40] , 
        \g2[27][39] , \g2[27][38] , \g2[27][37] , \g2[27][36] , \g2[27][35] , 
        \g2[27][34] , \g2[27][33] , \g2[27][32] , \g2[27][31] , \g2[27][30] , 
        \g2[27][29] , \g2[27][28] , \g2[27][27] , \g2[27][26] , \g2[27][25] , 
        \g2[27][24] , \g2[27][23] , \g2[27][22] , \g2[27][21] , \g2[27][20] , 
        \g2[27][19] , \g2[27][18] , \g2[27][17] , \g2[27][16] , \g2[27][15] , 
        \g2[27][14] , \g2[27][13] , \g2[27][12] , \g2[27][11] , \g2[27][10] , 
        \g2[27][9] , \g2[27][8] , \g2[27][7] , \g2[27][6] , \g2[27][5] , 
        \g2[27][4] , \g2[27][3] , \g2[27][2] , \g2[27][1] , 
        SYNOPSYS_UNCONNECTED__34}) );
  FullAdder \level3[0].x0  ( .a({\g2[0][63] , \g2[0][62] , \g2[0][61] , 
        \g2[0][60] , \g2[0][59] , \g2[0][58] , \g2[0][57] , \g2[0][56] , 
        \g2[0][55] , \g2[0][54] , \g2[0][53] , \g2[0][52] , \g2[0][51] , 
        \g2[0][50] , \g2[0][49] , \g2[0][48] , \g2[0][47] , \g2[0][46] , 
        \g2[0][45] , \g2[0][44] , \g2[0][43] , \g2[0][42] , \g2[0][41] , 
        \g2[0][40] , \g2[0][39] , \g2[0][38] , \g2[0][37] , \g2[0][36] , 
        \g2[0][35] , \g2[0][34] , \g2[0][33] , \g2[0][32] , \g2[0][31] , 
        \g2[0][30] , \g2[0][29] , \g2[0][28] , \g2[0][27] , \g2[0][26] , 
        \g2[0][25] , \g2[0][24] , \g2[0][23] , \g2[0][22] , \g2[0][21] , 
        \g2[0][20] , \g2[0][19] , \g2[0][18] , \g2[0][17] , \g2[0][16] , 
        \g2[0][15] , \g2[0][14] , \g2[0][13] , \g2[0][12] , \g2[0][11] , 
        \g2[0][10] , \g2[0][9] , \g2[0][8] , \g2[0][7] , \g2[0][6] , 
        \g2[0][5] , \g2[0][4] , \g2[0][3] , \g2[0][2] , \g2[0][1] , \g2[0][0] }), .b({\g2[1][63] , \g2[1][62] , \g2[1][61] , \g2[1][60] , \g2[1][59] , 
        \g2[1][58] , \g2[1][57] , \g2[1][56] , \g2[1][55] , \g2[1][54] , 
        \g2[1][53] , \g2[1][52] , \g2[1][51] , \g2[1][50] , \g2[1][49] , 
        \g2[1][48] , \g2[1][47] , \g2[1][46] , \g2[1][45] , \g2[1][44] , 
        \g2[1][43] , \g2[1][42] , \g2[1][41] , \g2[1][40] , \g2[1][39] , 
        \g2[1][38] , \g2[1][37] , \g2[1][36] , \g2[1][35] , \g2[1][34] , 
        \g2[1][33] , \g2[1][32] , \g2[1][31] , \g2[1][30] , \g2[1][29] , 
        \g2[1][28] , \g2[1][27] , \g2[1][26] , \g2[1][25] , \g2[1][24] , 
        \g2[1][23] , \g2[1][22] , \g2[1][21] , \g2[1][20] , \g2[1][19] , 
        \g2[1][18] , \g2[1][17] , \g2[1][16] , \g2[1][15] , \g2[1][14] , 
        \g2[1][13] , \g2[1][12] , \g2[1][11] , \g2[1][10] , \g2[1][9] , 
        \g2[1][8] , \g2[1][7] , \g2[1][6] , \g2[1][5] , \g2[1][4] , \g2[1][3] , 
        \g2[1][2] , \g2[1][1] , \g2[1][0] }), .cin({\g2[2][63] , \g2[2][62] , 
        \g2[2][61] , \g2[2][60] , \g2[2][59] , \g2[2][58] , \g2[2][57] , 
        \g2[2][56] , \g2[2][55] , \g2[2][54] , \g2[2][53] , \g2[2][52] , 
        \g2[2][51] , \g2[2][50] , \g2[2][49] , \g2[2][48] , \g2[2][47] , 
        \g2[2][46] , \g2[2][45] , \g2[2][44] , \g2[2][43] , \g2[2][42] , 
        \g2[2][41] , \g2[2][40] , \g2[2][39] , \g2[2][38] , \g2[2][37] , 
        \g2[2][36] , \g2[2][35] , \g2[2][34] , \g2[2][33] , \g2[2][32] , 
        \g2[2][31] , \g2[2][30] , \g2[2][29] , \g2[2][28] , \g2[2][27] , 
        \g2[2][26] , \g2[2][25] , \g2[2][24] , \g2[2][23] , \g2[2][22] , 
        \g2[2][21] , \g2[2][20] , \g2[2][19] , \g2[2][18] , \g2[2][17] , 
        \g2[2][16] , \g2[2][15] , \g2[2][14] , \g2[2][13] , \g2[2][12] , 
        \g2[2][11] , \g2[2][10] , \g2[2][9] , \g2[2][8] , \g2[2][7] , 
        \g2[2][6] , \g2[2][5] , \g2[2][4] , \g2[2][3] , \g2[2][2] , \g2[2][1] , 
        \g2[2][0] }), .sum({\g3[0][63] , \g3[0][62] , \g3[0][61] , \g3[0][60] , 
        \g3[0][59] , \g3[0][58] , \g3[0][57] , \g3[0][56] , \g3[0][55] , 
        \g3[0][54] , \g3[0][53] , \g3[0][52] , \g3[0][51] , \g3[0][50] , 
        \g3[0][49] , \g3[0][48] , \g3[0][47] , \g3[0][46] , \g3[0][45] , 
        \g3[0][44] , \g3[0][43] , \g3[0][42] , \g3[0][41] , \g3[0][40] , 
        \g3[0][39] , \g3[0][38] , \g3[0][37] , \g3[0][36] , \g3[0][35] , 
        \g3[0][34] , \g3[0][33] , \g3[0][32] , \g3[0][31] , \g3[0][30] , 
        \g3[0][29] , \g3[0][28] , \g3[0][27] , \g3[0][26] , \g3[0][25] , 
        \g3[0][24] , \g3[0][23] , \g3[0][22] , \g3[0][21] , \g3[0][20] , 
        \g3[0][19] , \g3[0][18] , \g3[0][17] , \g3[0][16] , \g3[0][15] , 
        \g3[0][14] , \g3[0][13] , \g3[0][12] , \g3[0][11] , \g3[0][10] , 
        \g3[0][9] , \g3[0][8] , \g3[0][7] , \g3[0][6] , \g3[0][5] , \g3[0][4] , 
        \g3[0][3] , \g3[0][2] , \g3[0][1] , \g3[0][0] }), .cout({\g3[9][63] , 
        \g3[9][62] , \g3[9][61] , \g3[9][60] , \g3[9][59] , \g3[9][58] , 
        \g3[9][57] , \g3[9][56] , \g3[9][55] , \g3[9][54] , \g3[9][53] , 
        \g3[9][52] , \g3[9][51] , \g3[9][50] , \g3[9][49] , \g3[9][48] , 
        \g3[9][47] , \g3[9][46] , \g3[9][45] , \g3[9][44] , \g3[9][43] , 
        \g3[9][42] , \g3[9][41] , \g3[9][40] , \g3[9][39] , \g3[9][38] , 
        \g3[9][37] , \g3[9][36] , \g3[9][35] , \g3[9][34] , \g3[9][33] , 
        \g3[9][32] , \g3[9][31] , \g3[9][30] , \g3[9][29] , \g3[9][28] , 
        \g3[9][27] , \g3[9][26] , \g3[9][25] , \g3[9][24] , \g3[9][23] , 
        \g3[9][22] , \g3[9][21] , \g3[9][20] , \g3[9][19] , \g3[9][18] , 
        \g3[9][17] , \g3[9][16] , \g3[9][15] , \g3[9][14] , \g3[9][13] , 
        \g3[9][12] , \g3[9][11] , \g3[9][10] , \g3[9][9] , \g3[9][8] , 
        \g3[9][7] , \g3[9][6] , \g3[9][5] , \g3[9][4] , \g3[9][3] , \g3[9][2] , 
        \g3[9][1] , SYNOPSYS_UNCONNECTED__35}) );
  FullAdder \level3[1].x0  ( .a({\g2[3][63] , \g2[3][62] , \g2[3][61] , 
        \g2[3][60] , \g2[3][59] , \g2[3][58] , \g2[3][57] , \g2[3][56] , 
        \g2[3][55] , \g2[3][54] , \g2[3][53] , \g2[3][52] , \g2[3][51] , 
        \g2[3][50] , \g2[3][49] , \g2[3][48] , \g2[3][47] , \g2[3][46] , 
        \g2[3][45] , \g2[3][44] , \g2[3][43] , \g2[3][42] , \g2[3][41] , 
        \g2[3][40] , \g2[3][39] , \g2[3][38] , \g2[3][37] , \g2[3][36] , 
        \g2[3][35] , \g2[3][34] , \g2[3][33] , \g2[3][32] , \g2[3][31] , 
        \g2[3][30] , \g2[3][29] , \g2[3][28] , \g2[3][27] , \g2[3][26] , 
        \g2[3][25] , \g2[3][24] , \g2[3][23] , \g2[3][22] , \g2[3][21] , 
        \g2[3][20] , \g2[3][19] , \g2[3][18] , \g2[3][17] , \g2[3][16] , 
        \g2[3][15] , \g2[3][14] , \g2[3][13] , \g2[3][12] , \g2[3][11] , 
        \g2[3][10] , \g2[3][9] , \g2[3][8] , \g2[3][7] , \g2[3][6] , 
        \g2[3][5] , \g2[3][4] , \g2[3][3] , \g2[3][2] , \g2[3][1] , \g2[3][0] }), .b({\g2[4][63] , \g2[4][62] , \g2[4][61] , \g2[4][60] , \g2[4][59] , 
        \g2[4][58] , \g2[4][57] , \g2[4][56] , \g2[4][55] , \g2[4][54] , 
        \g2[4][53] , \g2[4][52] , \g2[4][51] , \g2[4][50] , \g2[4][49] , 
        \g2[4][48] , \g2[4][47] , \g2[4][46] , \g2[4][45] , \g2[4][44] , 
        \g2[4][43] , \g2[4][42] , \g2[4][41] , \g2[4][40] , \g2[4][39] , 
        \g2[4][38] , \g2[4][37] , \g2[4][36] , \g2[4][35] , \g2[4][34] , 
        \g2[4][33] , \g2[4][32] , \g2[4][31] , \g2[4][30] , \g2[4][29] , 
        \g2[4][28] , \g2[4][27] , \g2[4][26] , \g2[4][25] , \g2[4][24] , 
        \g2[4][23] , \g2[4][22] , \g2[4][21] , \g2[4][20] , \g2[4][19] , 
        \g2[4][18] , \g2[4][17] , \g2[4][16] , \g2[4][15] , \g2[4][14] , 
        \g2[4][13] , \g2[4][12] , \g2[4][11] , \g2[4][10] , \g2[4][9] , 
        \g2[4][8] , \g2[4][7] , \g2[4][6] , \g2[4][5] , \g2[4][4] , \g2[4][3] , 
        \g2[4][2] , \g2[4][1] , \g2[4][0] }), .cin({\g2[5][63] , \g2[5][62] , 
        \g2[5][61] , \g2[5][60] , \g2[5][59] , \g2[5][58] , \g2[5][57] , 
        \g2[5][56] , \g2[5][55] , \g2[5][54] , \g2[5][53] , \g2[5][52] , 
        \g2[5][51] , \g2[5][50] , \g2[5][49] , \g2[5][48] , \g2[5][47] , 
        \g2[5][46] , \g2[5][45] , \g2[5][44] , \g2[5][43] , \g2[5][42] , 
        \g2[5][41] , \g2[5][40] , \g2[5][39] , \g2[5][38] , \g2[5][37] , 
        \g2[5][36] , \g2[5][35] , \g2[5][34] , \g2[5][33] , \g2[5][32] , 
        \g2[5][31] , \g2[5][30] , \g2[5][29] , \g2[5][28] , \g2[5][27] , 
        \g2[5][26] , \g2[5][25] , \g2[5][24] , \g2[5][23] , \g2[5][22] , 
        \g2[5][21] , \g2[5][20] , \g2[5][19] , \g2[5][18] , \g2[5][17] , 
        \g2[5][16] , \g2[5][15] , \g2[5][14] , \g2[5][13] , \g2[5][12] , 
        \g2[5][11] , \g2[5][10] , \g2[5][9] , \g2[5][8] , \g2[5][7] , 
        \g2[5][6] , \g2[5][5] , \g2[5][4] , \g2[5][3] , \g2[5][2] , \g2[5][1] , 
        \g2[5][0] }), .sum({\g3[1][63] , \g3[1][62] , \g3[1][61] , \g3[1][60] , 
        \g3[1][59] , \g3[1][58] , \g3[1][57] , \g3[1][56] , \g3[1][55] , 
        \g3[1][54] , \g3[1][53] , \g3[1][52] , \g3[1][51] , \g3[1][50] , 
        \g3[1][49] , \g3[1][48] , \g3[1][47] , \g3[1][46] , \g3[1][45] , 
        \g3[1][44] , \g3[1][43] , \g3[1][42] , \g3[1][41] , \g3[1][40] , 
        \g3[1][39] , \g3[1][38] , \g3[1][37] , \g3[1][36] , \g3[1][35] , 
        \g3[1][34] , \g3[1][33] , \g3[1][32] , \g3[1][31] , \g3[1][30] , 
        \g3[1][29] , \g3[1][28] , \g3[1][27] , \g3[1][26] , \g3[1][25] , 
        \g3[1][24] , \g3[1][23] , \g3[1][22] , \g3[1][21] , \g3[1][20] , 
        \g3[1][19] , \g3[1][18] , \g3[1][17] , \g3[1][16] , \g3[1][15] , 
        \g3[1][14] , \g3[1][13] , \g3[1][12] , \g3[1][11] , \g3[1][10] , 
        \g3[1][9] , \g3[1][8] , \g3[1][7] , \g3[1][6] , \g3[1][5] , \g3[1][4] , 
        \g3[1][3] , \g3[1][2] , \g3[1][1] , \g3[1][0] }), .cout({\g3[10][63] , 
        \g3[10][62] , \g3[10][61] , \g3[10][60] , \g3[10][59] , \g3[10][58] , 
        \g3[10][57] , \g3[10][56] , \g3[10][55] , \g3[10][54] , \g3[10][53] , 
        \g3[10][52] , \g3[10][51] , \g3[10][50] , \g3[10][49] , \g3[10][48] , 
        \g3[10][47] , \g3[10][46] , \g3[10][45] , \g3[10][44] , \g3[10][43] , 
        \g3[10][42] , \g3[10][41] , \g3[10][40] , \g3[10][39] , \g3[10][38] , 
        \g3[10][37] , \g3[10][36] , \g3[10][35] , \g3[10][34] , \g3[10][33] , 
        \g3[10][32] , \g3[10][31] , \g3[10][30] , \g3[10][29] , \g3[10][28] , 
        \g3[10][27] , \g3[10][26] , \g3[10][25] , \g3[10][24] , \g3[10][23] , 
        \g3[10][22] , \g3[10][21] , \g3[10][20] , \g3[10][19] , \g3[10][18] , 
        \g3[10][17] , \g3[10][16] , \g3[10][15] , \g3[10][14] , \g3[10][13] , 
        \g3[10][12] , \g3[10][11] , \g3[10][10] , \g3[10][9] , \g3[10][8] , 
        \g3[10][7] , \g3[10][6] , \g3[10][5] , \g3[10][4] , \g3[10][3] , 
        \g3[10][2] , \g3[10][1] , SYNOPSYS_UNCONNECTED__36}) );
  FullAdder \level3[2].x0  ( .a({\g2[6][63] , \g2[6][62] , \g2[6][61] , 
        \g2[6][60] , \g2[6][59] , \g2[6][58] , \g2[6][57] , \g2[6][56] , 
        \g2[6][55] , \g2[6][54] , \g2[6][53] , \g2[6][52] , \g2[6][51] , 
        \g2[6][50] , \g2[6][49] , \g2[6][48] , \g2[6][47] , \g2[6][46] , 
        \g2[6][45] , \g2[6][44] , \g2[6][43] , \g2[6][42] , \g2[6][41] , 
        \g2[6][40] , \g2[6][39] , \g2[6][38] , \g2[6][37] , \g2[6][36] , 
        \g2[6][35] , \g2[6][34] , \g2[6][33] , \g2[6][32] , \g2[6][31] , 
        \g2[6][30] , \g2[6][29] , \g2[6][28] , \g2[6][27] , \g2[6][26] , 
        \g2[6][25] , \g2[6][24] , \g2[6][23] , \g2[6][22] , \g2[6][21] , 
        \g2[6][20] , \g2[6][19] , \g2[6][18] , \g2[6][17] , \g2[6][16] , 
        \g2[6][15] , \g2[6][14] , \g2[6][13] , \g2[6][12] , \g2[6][11] , 
        \g2[6][10] , \g2[6][9] , \g2[6][8] , \g2[6][7] , \g2[6][6] , 
        \g2[6][5] , \g2[6][4] , \g2[6][3] , \g2[6][2] , \g2[6][1] , \g2[6][0] }), .b({\g2[7][63] , \g2[7][62] , \g2[7][61] , \g2[7][60] , \g2[7][59] , 
        \g2[7][58] , \g2[7][57] , \g2[7][56] , \g2[7][55] , \g2[7][54] , 
        \g2[7][53] , \g2[7][52] , \g2[7][51] , \g2[7][50] , \g2[7][49] , 
        \g2[7][48] , \g2[7][47] , \g2[7][46] , \g2[7][45] , \g2[7][44] , 
        \g2[7][43] , \g2[7][42] , \g2[7][41] , \g2[7][40] , \g2[7][39] , 
        \g2[7][38] , \g2[7][37] , \g2[7][36] , \g2[7][35] , \g2[7][34] , 
        \g2[7][33] , \g2[7][32] , \g2[7][31] , \g2[7][30] , \g2[7][29] , 
        \g2[7][28] , \g2[7][27] , \g2[7][26] , \g2[7][25] , \g2[7][24] , 
        \g2[7][23] , \g2[7][22] , \g2[7][21] , \g2[7][20] , \g2[7][19] , 
        \g2[7][18] , \g2[7][17] , \g2[7][16] , \g2[7][15] , \g2[7][14] , 
        \g2[7][13] , \g2[7][12] , \g2[7][11] , \g2[7][10] , \g2[7][9] , 
        \g2[7][8] , \g2[7][7] , \g2[7][6] , \g2[7][5] , \g2[7][4] , \g2[7][3] , 
        \g2[7][2] , \g2[7][1] , \g2[7][0] }), .cin({\g2[8][63] , \g2[8][62] , 
        \g2[8][61] , \g2[8][60] , \g2[8][59] , \g2[8][58] , \g2[8][57] , 
        \g2[8][56] , \g2[8][55] , \g2[8][54] , \g2[8][53] , \g2[8][52] , 
        \g2[8][51] , \g2[8][50] , \g2[8][49] , \g2[8][48] , \g2[8][47] , 
        \g2[8][46] , \g2[8][45] , \g2[8][44] , \g2[8][43] , \g2[8][42] , 
        \g2[8][41] , \g2[8][40] , \g2[8][39] , \g2[8][38] , \g2[8][37] , 
        \g2[8][36] , \g2[8][35] , \g2[8][34] , \g2[8][33] , \g2[8][32] , 
        \g2[8][31] , \g2[8][30] , \g2[8][29] , \g2[8][28] , \g2[8][27] , 
        \g2[8][26] , \g2[8][25] , \g2[8][24] , \g2[8][23] , \g2[8][22] , 
        \g2[8][21] , \g2[8][20] , \g2[8][19] , \g2[8][18] , \g2[8][17] , 
        \g2[8][16] , \g2[8][15] , \g2[8][14] , \g2[8][13] , \g2[8][12] , 
        \g2[8][11] , \g2[8][10] , \g2[8][9] , \g2[8][8] , \g2[8][7] , 
        \g2[8][6] , \g2[8][5] , \g2[8][4] , \g2[8][3] , \g2[8][2] , \g2[8][1] , 
        \g2[8][0] }), .sum({\g3[2][63] , \g3[2][62] , \g3[2][61] , \g3[2][60] , 
        \g3[2][59] , \g3[2][58] , \g3[2][57] , \g3[2][56] , \g3[2][55] , 
        \g3[2][54] , \g3[2][53] , \g3[2][52] , \g3[2][51] , \g3[2][50] , 
        \g3[2][49] , \g3[2][48] , \g3[2][47] , \g3[2][46] , \g3[2][45] , 
        \g3[2][44] , \g3[2][43] , \g3[2][42] , \g3[2][41] , \g3[2][40] , 
        \g3[2][39] , \g3[2][38] , \g3[2][37] , \g3[2][36] , \g3[2][35] , 
        \g3[2][34] , \g3[2][33] , \g3[2][32] , \g3[2][31] , \g3[2][30] , 
        \g3[2][29] , \g3[2][28] , \g3[2][27] , \g3[2][26] , \g3[2][25] , 
        \g3[2][24] , \g3[2][23] , \g3[2][22] , \g3[2][21] , \g3[2][20] , 
        \g3[2][19] , \g3[2][18] , \g3[2][17] , \g3[2][16] , \g3[2][15] , 
        \g3[2][14] , \g3[2][13] , \g3[2][12] , \g3[2][11] , \g3[2][10] , 
        \g3[2][9] , \g3[2][8] , \g3[2][7] , \g3[2][6] , \g3[2][5] , \g3[2][4] , 
        \g3[2][3] , \g3[2][2] , \g3[2][1] , \g3[2][0] }), .cout({\g3[11][63] , 
        \g3[11][62] , \g3[11][61] , \g3[11][60] , \g3[11][59] , \g3[11][58] , 
        \g3[11][57] , \g3[11][56] , \g3[11][55] , \g3[11][54] , \g3[11][53] , 
        \g3[11][52] , \g3[11][51] , \g3[11][50] , \g3[11][49] , \g3[11][48] , 
        \g3[11][47] , \g3[11][46] , \g3[11][45] , \g3[11][44] , \g3[11][43] , 
        \g3[11][42] , \g3[11][41] , \g3[11][40] , \g3[11][39] , \g3[11][38] , 
        \g3[11][37] , \g3[11][36] , \g3[11][35] , \g3[11][34] , \g3[11][33] , 
        \g3[11][32] , \g3[11][31] , \g3[11][30] , \g3[11][29] , \g3[11][28] , 
        \g3[11][27] , \g3[11][26] , \g3[11][25] , \g3[11][24] , \g3[11][23] , 
        \g3[11][22] , \g3[11][21] , \g3[11][20] , \g3[11][19] , \g3[11][18] , 
        \g3[11][17] , \g3[11][16] , \g3[11][15] , \g3[11][14] , \g3[11][13] , 
        \g3[11][12] , \g3[11][11] , \g3[11][10] , \g3[11][9] , \g3[11][8] , 
        \g3[11][7] , \g3[11][6] , \g3[11][5] , \g3[11][4] , \g3[11][3] , 
        \g3[11][2] , \g3[11][1] , SYNOPSYS_UNCONNECTED__37}) );
  FullAdder \level3[3].x0  ( .a({\g2[9][63] , \g2[9][62] , \g2[9][61] , 
        \g2[9][60] , \g2[9][59] , \g2[9][58] , \g2[9][57] , \g2[9][56] , 
        \g2[9][55] , \g2[9][54] , \g2[9][53] , \g2[9][52] , \g2[9][51] , 
        \g2[9][50] , \g2[9][49] , \g2[9][48] , \g2[9][47] , \g2[9][46] , 
        \g2[9][45] , \g2[9][44] , \g2[9][43] , \g2[9][42] , \g2[9][41] , 
        \g2[9][40] , \g2[9][39] , \g2[9][38] , \g2[9][37] , \g2[9][36] , 
        \g2[9][35] , \g2[9][34] , \g2[9][33] , \g2[9][32] , \g2[9][31] , 
        \g2[9][30] , \g2[9][29] , \g2[9][28] , \g2[9][27] , \g2[9][26] , 
        \g2[9][25] , \g2[9][24] , \g2[9][23] , \g2[9][22] , \g2[9][21] , 
        \g2[9][20] , \g2[9][19] , \g2[9][18] , \g2[9][17] , \g2[9][16] , 
        \g2[9][15] , \g2[9][14] , \g2[9][13] , \g2[9][12] , \g2[9][11] , 
        \g2[9][10] , \g2[9][9] , \g2[9][8] , \g2[9][7] , \g2[9][6] , 
        \g2[9][5] , \g2[9][4] , \g2[9][3] , \g2[9][2] , \g2[9][1] , \g2[9][0] }), .b({\g2[10][63] , \g2[10][62] , \g2[10][61] , \g2[10][60] , \g2[10][59] , 
        \g2[10][58] , \g2[10][57] , \g2[10][56] , \g2[10][55] , \g2[10][54] , 
        \g2[10][53] , \g2[10][52] , \g2[10][51] , \g2[10][50] , \g2[10][49] , 
        \g2[10][48] , \g2[10][47] , \g2[10][46] , \g2[10][45] , \g2[10][44] , 
        \g2[10][43] , \g2[10][42] , \g2[10][41] , \g2[10][40] , \g2[10][39] , 
        \g2[10][38] , \g2[10][37] , \g2[10][36] , \g2[10][35] , \g2[10][34] , 
        \g2[10][33] , \g2[10][32] , \g2[10][31] , \g2[10][30] , \g2[10][29] , 
        \g2[10][28] , \g2[10][27] , \g2[10][26] , \g2[10][25] , \g2[10][24] , 
        \g2[10][23] , \g2[10][22] , \g2[10][21] , \g2[10][20] , \g2[10][19] , 
        \g2[10][18] , \g2[10][17] , \g2[10][16] , \g2[10][15] , \g2[10][14] , 
        \g2[10][13] , \g2[10][12] , \g2[10][11] , \g2[10][10] , \g2[10][9] , 
        \g2[10][8] , \g2[10][7] , \g2[10][6] , \g2[10][5] , \g2[10][4] , 
        \g2[10][3] , \g2[10][2] , \g2[10][1] , \g2[10][0] }), .cin({
        \g2[11][63] , \g2[11][62] , \g2[11][61] , \g2[11][60] , \g2[11][59] , 
        \g2[11][58] , \g2[11][57] , \g2[11][56] , \g2[11][55] , \g2[11][54] , 
        \g2[11][53] , \g2[11][52] , \g2[11][51] , \g2[11][50] , \g2[11][49] , 
        \g2[11][48] , \g2[11][47] , \g2[11][46] , \g2[11][45] , \g2[11][44] , 
        \g2[11][43] , \g2[11][42] , \g2[11][41] , \g2[11][40] , \g2[11][39] , 
        \g2[11][38] , \g2[11][37] , \g2[11][36] , \g2[11][35] , \g2[11][34] , 
        \g2[11][33] , \g2[11][32] , \g2[11][31] , \g2[11][30] , \g2[11][29] , 
        \g2[11][28] , \g2[11][27] , \g2[11][26] , \g2[11][25] , \g2[11][24] , 
        \g2[11][23] , \g2[11][22] , \g2[11][21] , \g2[11][20] , \g2[11][19] , 
        \g2[11][18] , \g2[11][17] , \g2[11][16] , \g2[11][15] , \g2[11][14] , 
        \g2[11][13] , \g2[11][12] , \g2[11][11] , \g2[11][10] , \g2[11][9] , 
        \g2[11][8] , \g2[11][7] , \g2[11][6] , \g2[11][5] , \g2[11][4] , 
        \g2[11][3] , \g2[11][2] , \g2[11][1] , \g2[11][0] }), .sum({
        \g3[3][63] , \g3[3][62] , \g3[3][61] , \g3[3][60] , \g3[3][59] , 
        \g3[3][58] , \g3[3][57] , \g3[3][56] , \g3[3][55] , \g3[3][54] , 
        \g3[3][53] , \g3[3][52] , \g3[3][51] , \g3[3][50] , \g3[3][49] , 
        \g3[3][48] , \g3[3][47] , \g3[3][46] , \g3[3][45] , \g3[3][44] , 
        \g3[3][43] , \g3[3][42] , \g3[3][41] , \g3[3][40] , \g3[3][39] , 
        \g3[3][38] , \g3[3][37] , \g3[3][36] , \g3[3][35] , \g3[3][34] , 
        \g3[3][33] , \g3[3][32] , \g3[3][31] , \g3[3][30] , \g3[3][29] , 
        \g3[3][28] , \g3[3][27] , \g3[3][26] , \g3[3][25] , \g3[3][24] , 
        \g3[3][23] , \g3[3][22] , \g3[3][21] , \g3[3][20] , \g3[3][19] , 
        \g3[3][18] , \g3[3][17] , \g3[3][16] , \g3[3][15] , \g3[3][14] , 
        \g3[3][13] , \g3[3][12] , \g3[3][11] , \g3[3][10] , \g3[3][9] , 
        \g3[3][8] , \g3[3][7] , \g3[3][6] , \g3[3][5] , \g3[3][4] , \g3[3][3] , 
        \g3[3][2] , \g3[3][1] , \g3[3][0] }), .cout({\g3[12][63] , 
        \g3[12][62] , \g3[12][61] , \g3[12][60] , \g3[12][59] , \g3[12][58] , 
        \g3[12][57] , \g3[12][56] , \g3[12][55] , \g3[12][54] , \g3[12][53] , 
        \g3[12][52] , \g3[12][51] , \g3[12][50] , \g3[12][49] , \g3[12][48] , 
        \g3[12][47] , \g3[12][46] , \g3[12][45] , \g3[12][44] , \g3[12][43] , 
        \g3[12][42] , \g3[12][41] , \g3[12][40] , \g3[12][39] , \g3[12][38] , 
        \g3[12][37] , \g3[12][36] , \g3[12][35] , \g3[12][34] , \g3[12][33] , 
        \g3[12][32] , \g3[12][31] , \g3[12][30] , \g3[12][29] , \g3[12][28] , 
        \g3[12][27] , \g3[12][26] , \g3[12][25] , \g3[12][24] , \g3[12][23] , 
        \g3[12][22] , \g3[12][21] , \g3[12][20] , \g3[12][19] , \g3[12][18] , 
        \g3[12][17] , \g3[12][16] , \g3[12][15] , \g3[12][14] , \g3[12][13] , 
        \g3[12][12] , \g3[12][11] , \g3[12][10] , \g3[12][9] , \g3[12][8] , 
        \g3[12][7] , \g3[12][6] , \g3[12][5] , \g3[12][4] , \g3[12][3] , 
        \g3[12][2] , \g3[12][1] , SYNOPSYS_UNCONNECTED__38}) );
  FullAdder \level3[4].x0  ( .a({\g2[12][63] , \g2[12][62] , \g2[12][61] , 
        \g2[12][60] , \g2[12][59] , \g2[12][58] , \g2[12][57] , \g2[12][56] , 
        \g2[12][55] , \g2[12][54] , \g2[12][53] , \g2[12][52] , \g2[12][51] , 
        \g2[12][50] , \g2[12][49] , \g2[12][48] , \g2[12][47] , \g2[12][46] , 
        \g2[12][45] , \g2[12][44] , \g2[12][43] , \g2[12][42] , \g2[12][41] , 
        \g2[12][40] , \g2[12][39] , \g2[12][38] , \g2[12][37] , \g2[12][36] , 
        \g2[12][35] , \g2[12][34] , \g2[12][33] , \g2[12][32] , \g2[12][31] , 
        \g2[12][30] , \g2[12][29] , \g2[12][28] , \g2[12][27] , \g2[12][26] , 
        \g2[12][25] , \g2[12][24] , \g2[12][23] , \g2[12][22] , \g2[12][21] , 
        \g2[12][20] , \g2[12][19] , \g2[12][18] , \g2[12][17] , \g2[12][16] , 
        \g2[12][15] , \g2[12][14] , \g2[12][13] , \g2[12][12] , \g2[12][11] , 
        \g2[12][10] , \g2[12][9] , \g2[12][8] , \g2[12][7] , \g2[12][6] , 
        \g2[12][5] , \g2[12][4] , \g2[12][3] , \g2[12][2] , \g2[12][1] , 
        \g2[12][0] }), .b({\g2[13][63] , \g2[13][62] , \g2[13][61] , 
        \g2[13][60] , \g2[13][59] , \g2[13][58] , \g2[13][57] , \g2[13][56] , 
        \g2[13][55] , \g2[13][54] , \g2[13][53] , \g2[13][52] , \g2[13][51] , 
        \g2[13][50] , \g2[13][49] , \g2[13][48] , \g2[13][47] , \g2[13][46] , 
        \g2[13][45] , \g2[13][44] , \g2[13][43] , \g2[13][42] , \g2[13][41] , 
        \g2[13][40] , \g2[13][39] , \g2[13][38] , \g2[13][37] , \g2[13][36] , 
        \g2[13][35] , \g2[13][34] , \g2[13][33] , \g2[13][32] , \g2[13][31] , 
        \g2[13][30] , \g2[13][29] , \g2[13][28] , \g2[13][27] , \g2[13][26] , 
        \g2[13][25] , \g2[13][24] , \g2[13][23] , \g2[13][22] , \g2[13][21] , 
        \g2[13][20] , \g2[13][19] , \g2[13][18] , \g2[13][17] , \g2[13][16] , 
        \g2[13][15] , \g2[13][14] , \g2[13][13] , \g2[13][12] , \g2[13][11] , 
        \g2[13][10] , \g2[13][9] , \g2[13][8] , \g2[13][7] , \g2[13][6] , 
        \g2[13][5] , \g2[13][4] , \g2[13][3] , \g2[13][2] , \g2[13][1] , 
        \g2[13][0] }), .cin({\g2[14][63] , \g2[14][62] , \g2[14][61] , 
        \g2[14][60] , \g2[14][59] , \g2[14][58] , \g2[14][57] , \g2[14][56] , 
        \g2[14][55] , \g2[14][54] , \g2[14][53] , \g2[14][52] , \g2[14][51] , 
        \g2[14][50] , \g2[14][49] , \g2[14][48] , \g2[14][47] , \g2[14][46] , 
        \g2[14][45] , \g2[14][44] , \g2[14][43] , \g2[14][42] , \g2[14][41] , 
        \g2[14][40] , \g2[14][39] , \g2[14][38] , \g2[14][37] , \g2[14][36] , 
        \g2[14][35] , \g2[14][34] , \g2[14][33] , \g2[14][32] , \g2[14][31] , 
        \g2[14][30] , \g2[14][29] , \g2[14][28] , \g2[14][27] , \g2[14][26] , 
        \g2[14][25] , \g2[14][24] , \g2[14][23] , \g2[14][22] , \g2[14][21] , 
        \g2[14][20] , \g2[14][19] , \g2[14][18] , \g2[14][17] , \g2[14][16] , 
        \g2[14][15] , \g2[14][14] , \g2[14][13] , \g2[14][12] , \g2[14][11] , 
        \g2[14][10] , \g2[14][9] , \g2[14][8] , \g2[14][7] , \g2[14][6] , 
        \g2[14][5] , \g2[14][4] , \g2[14][3] , \g2[14][2] , \g2[14][1] , 1'b0}), .sum({\g3[4][63] , \g3[4][62] , \g3[4][61] , \g3[4][60] , \g3[4][59] , 
        \g3[4][58] , \g3[4][57] , \g3[4][56] , \g3[4][55] , \g3[4][54] , 
        \g3[4][53] , \g3[4][52] , \g3[4][51] , \g3[4][50] , \g3[4][49] , 
        \g3[4][48] , \g3[4][47] , \g3[4][46] , \g3[4][45] , \g3[4][44] , 
        \g3[4][43] , \g3[4][42] , \g3[4][41] , \g3[4][40] , \g3[4][39] , 
        \g3[4][38] , \g3[4][37] , \g3[4][36] , \g3[4][35] , \g3[4][34] , 
        \g3[4][33] , \g3[4][32] , \g3[4][31] , \g3[4][30] , \g3[4][29] , 
        \g3[4][28] , \g3[4][27] , \g3[4][26] , \g3[4][25] , \g3[4][24] , 
        \g3[4][23] , \g3[4][22] , \g3[4][21] , \g3[4][20] , \g3[4][19] , 
        \g3[4][18] , \g3[4][17] , \g3[4][16] , \g3[4][15] , \g3[4][14] , 
        \g3[4][13] , \g3[4][12] , \g3[4][11] , \g3[4][10] , \g3[4][9] , 
        \g3[4][8] , \g3[4][7] , \g3[4][6] , \g3[4][5] , \g3[4][4] , \g3[4][3] , 
        \g3[4][2] , \g3[4][1] , \g3[4][0] }), .cout({\g3[13][63] , 
        \g3[13][62] , \g3[13][61] , \g3[13][60] , \g3[13][59] , \g3[13][58] , 
        \g3[13][57] , \g3[13][56] , \g3[13][55] , \g3[13][54] , \g3[13][53] , 
        \g3[13][52] , \g3[13][51] , \g3[13][50] , \g3[13][49] , \g3[13][48] , 
        \g3[13][47] , \g3[13][46] , \g3[13][45] , \g3[13][44] , \g3[13][43] , 
        \g3[13][42] , \g3[13][41] , \g3[13][40] , \g3[13][39] , \g3[13][38] , 
        \g3[13][37] , \g3[13][36] , \g3[13][35] , \g3[13][34] , \g3[13][33] , 
        \g3[13][32] , \g3[13][31] , \g3[13][30] , \g3[13][29] , \g3[13][28] , 
        \g3[13][27] , \g3[13][26] , \g3[13][25] , \g3[13][24] , \g3[13][23] , 
        \g3[13][22] , \g3[13][21] , \g3[13][20] , \g3[13][19] , \g3[13][18] , 
        \g3[13][17] , \g3[13][16] , \g3[13][15] , \g3[13][14] , \g3[13][13] , 
        \g3[13][12] , \g3[13][11] , \g3[13][10] , \g3[13][9] , \g3[13][8] , 
        \g3[13][7] , \g3[13][6] , \g3[13][5] , \g3[13][4] , \g3[13][3] , 
        \g3[13][2] , \g3[13][1] , SYNOPSYS_UNCONNECTED__39}) );
  FullAdder \level3[5].x0  ( .a({\g2[15][63] , \g2[15][62] , \g2[15][61] , 
        \g2[15][60] , \g2[15][59] , \g2[15][58] , \g2[15][57] , \g2[15][56] , 
        \g2[15][55] , \g2[15][54] , \g2[15][53] , \g2[15][52] , \g2[15][51] , 
        \g2[15][50] , \g2[15][49] , \g2[15][48] , \g2[15][47] , \g2[15][46] , 
        \g2[15][45] , \g2[15][44] , \g2[15][43] , \g2[15][42] , \g2[15][41] , 
        \g2[15][40] , \g2[15][39] , \g2[15][38] , \g2[15][37] , \g2[15][36] , 
        \g2[15][35] , \g2[15][34] , \g2[15][33] , \g2[15][32] , \g2[15][31] , 
        \g2[15][30] , \g2[15][29] , \g2[15][28] , \g2[15][27] , \g2[15][26] , 
        \g2[15][25] , \g2[15][24] , \g2[15][23] , \g2[15][22] , \g2[15][21] , 
        \g2[15][20] , \g2[15][19] , \g2[15][18] , \g2[15][17] , \g2[15][16] , 
        \g2[15][15] , \g2[15][14] , \g2[15][13] , \g2[15][12] , \g2[15][11] , 
        \g2[15][10] , \g2[15][9] , \g2[15][8] , \g2[15][7] , \g2[15][6] , 
        \g2[15][5] , \g2[15][4] , \g2[15][3] , \g2[15][2] , \g2[15][1] , 1'b0}), .b({\g2[16][63] , \g2[16][62] , \g2[16][61] , \g2[16][60] , \g2[16][59] , 
        \g2[16][58] , \g2[16][57] , \g2[16][56] , \g2[16][55] , \g2[16][54] , 
        \g2[16][53] , \g2[16][52] , \g2[16][51] , \g2[16][50] , \g2[16][49] , 
        \g2[16][48] , \g2[16][47] , \g2[16][46] , \g2[16][45] , \g2[16][44] , 
        \g2[16][43] , \g2[16][42] , \g2[16][41] , \g2[16][40] , \g2[16][39] , 
        \g2[16][38] , \g2[16][37] , \g2[16][36] , \g2[16][35] , \g2[16][34] , 
        \g2[16][33] , \g2[16][32] , \g2[16][31] , \g2[16][30] , \g2[16][29] , 
        \g2[16][28] , \g2[16][27] , \g2[16][26] , \g2[16][25] , \g2[16][24] , 
        \g2[16][23] , \g2[16][22] , \g2[16][21] , \g2[16][20] , \g2[16][19] , 
        \g2[16][18] , \g2[16][17] , \g2[16][16] , \g2[16][15] , \g2[16][14] , 
        \g2[16][13] , \g2[16][12] , \g2[16][11] , \g2[16][10] , \g2[16][9] , 
        \g2[16][8] , \g2[16][7] , \g2[16][6] , \g2[16][5] , \g2[16][4] , 
        \g2[16][3] , \g2[16][2] , \g2[16][1] , 1'b0}), .cin({\g2[17][63] , 
        \g2[17][62] , \g2[17][61] , \g2[17][60] , \g2[17][59] , \g2[17][58] , 
        \g2[17][57] , \g2[17][56] , \g2[17][55] , \g2[17][54] , \g2[17][53] , 
        \g2[17][52] , \g2[17][51] , \g2[17][50] , \g2[17][49] , \g2[17][48] , 
        \g2[17][47] , \g2[17][46] , \g2[17][45] , \g2[17][44] , \g2[17][43] , 
        \g2[17][42] , \g2[17][41] , \g2[17][40] , \g2[17][39] , \g2[17][38] , 
        \g2[17][37] , \g2[17][36] , \g2[17][35] , \g2[17][34] , \g2[17][33] , 
        \g2[17][32] , \g2[17][31] , \g2[17][30] , \g2[17][29] , \g2[17][28] , 
        \g2[17][27] , \g2[17][26] , \g2[17][25] , \g2[17][24] , \g2[17][23] , 
        \g2[17][22] , \g2[17][21] , \g2[17][20] , \g2[17][19] , \g2[17][18] , 
        \g2[17][17] , \g2[17][16] , \g2[17][15] , \g2[17][14] , \g2[17][13] , 
        \g2[17][12] , \g2[17][11] , \g2[17][10] , \g2[17][9] , \g2[17][8] , 
        \g2[17][7] , \g2[17][6] , \g2[17][5] , \g2[17][4] , \g2[17][3] , 
        \g2[17][2] , \g2[17][1] , 1'b0}), .sum({\g3[5][63] , \g3[5][62] , 
        \g3[5][61] , \g3[5][60] , \g3[5][59] , \g3[5][58] , \g3[5][57] , 
        \g3[5][56] , \g3[5][55] , \g3[5][54] , \g3[5][53] , \g3[5][52] , 
        \g3[5][51] , \g3[5][50] , \g3[5][49] , \g3[5][48] , \g3[5][47] , 
        \g3[5][46] , \g3[5][45] , \g3[5][44] , \g3[5][43] , \g3[5][42] , 
        \g3[5][41] , \g3[5][40] , \g3[5][39] , \g3[5][38] , \g3[5][37] , 
        \g3[5][36] , \g3[5][35] , \g3[5][34] , \g3[5][33] , \g3[5][32] , 
        \g3[5][31] , \g3[5][30] , \g3[5][29] , \g3[5][28] , \g3[5][27] , 
        \g3[5][26] , \g3[5][25] , \g3[5][24] , \g3[5][23] , \g3[5][22] , 
        \g3[5][21] , \g3[5][20] , \g3[5][19] , \g3[5][18] , \g3[5][17] , 
        \g3[5][16] , \g3[5][15] , \g3[5][14] , \g3[5][13] , \g3[5][12] , 
        \g3[5][11] , \g3[5][10] , \g3[5][9] , \g3[5][8] , \g3[5][7] , 
        \g3[5][6] , \g3[5][5] , \g3[5][4] , \g3[5][3] , \g3[5][2] , \g3[5][1] , 
        \g3[5][0] }), .cout({\g3[14][63] , \g3[14][62] , \g3[14][61] , 
        \g3[14][60] , \g3[14][59] , \g3[14][58] , \g3[14][57] , \g3[14][56] , 
        \g3[14][55] , \g3[14][54] , \g3[14][53] , \g3[14][52] , \g3[14][51] , 
        \g3[14][50] , \g3[14][49] , \g3[14][48] , \g3[14][47] , \g3[14][46] , 
        \g3[14][45] , \g3[14][44] , \g3[14][43] , \g3[14][42] , \g3[14][41] , 
        \g3[14][40] , \g3[14][39] , \g3[14][38] , \g3[14][37] , \g3[14][36] , 
        \g3[14][35] , \g3[14][34] , \g3[14][33] , \g3[14][32] , \g3[14][31] , 
        \g3[14][30] , \g3[14][29] , \g3[14][28] , \g3[14][27] , \g3[14][26] , 
        \g3[14][25] , \g3[14][24] , \g3[14][23] , \g3[14][22] , \g3[14][21] , 
        \g3[14][20] , \g3[14][19] , \g3[14][18] , \g3[14][17] , \g3[14][16] , 
        \g3[14][15] , \g3[14][14] , \g3[14][13] , \g3[14][12] , \g3[14][11] , 
        \g3[14][10] , \g3[14][9] , \g3[14][8] , \g3[14][7] , \g3[14][6] , 
        \g3[14][5] , \g3[14][4] , \g3[14][3] , \g3[14][2] , \g3[14][1] , 
        SYNOPSYS_UNCONNECTED__40}) );
  FullAdder \level3[6].x0  ( .a({\g2[18][63] , \g2[18][62] , \g2[18][61] , 
        \g2[18][60] , \g2[18][59] , \g2[18][58] , \g2[18][57] , \g2[18][56] , 
        \g2[18][55] , \g2[18][54] , \g2[18][53] , \g2[18][52] , \g2[18][51] , 
        \g2[18][50] , \g2[18][49] , \g2[18][48] , \g2[18][47] , \g2[18][46] , 
        \g2[18][45] , \g2[18][44] , \g2[18][43] , \g2[18][42] , \g2[18][41] , 
        \g2[18][40] , \g2[18][39] , \g2[18][38] , \g2[18][37] , \g2[18][36] , 
        \g2[18][35] , \g2[18][34] , \g2[18][33] , \g2[18][32] , \g2[18][31] , 
        \g2[18][30] , \g2[18][29] , \g2[18][28] , \g2[18][27] , \g2[18][26] , 
        \g2[18][25] , \g2[18][24] , \g2[18][23] , \g2[18][22] , \g2[18][21] , 
        \g2[18][20] , \g2[18][19] , \g2[18][18] , \g2[18][17] , \g2[18][16] , 
        \g2[18][15] , \g2[18][14] , \g2[18][13] , \g2[18][12] , \g2[18][11] , 
        \g2[18][10] , \g2[18][9] , \g2[18][8] , \g2[18][7] , \g2[18][6] , 
        \g2[18][5] , \g2[18][4] , \g2[18][3] , \g2[18][2] , \g2[18][1] , 1'b0}), .b({\g2[19][63] , \g2[19][62] , \g2[19][61] , \g2[19][60] , \g2[19][59] , 
        \g2[19][58] , \g2[19][57] , \g2[19][56] , \g2[19][55] , \g2[19][54] , 
        \g2[19][53] , \g2[19][52] , \g2[19][51] , \g2[19][50] , \g2[19][49] , 
        \g2[19][48] , \g2[19][47] , \g2[19][46] , \g2[19][45] , \g2[19][44] , 
        \g2[19][43] , \g2[19][42] , \g2[19][41] , \g2[19][40] , \g2[19][39] , 
        \g2[19][38] , \g2[19][37] , \g2[19][36] , \g2[19][35] , \g2[19][34] , 
        \g2[19][33] , \g2[19][32] , \g2[19][31] , \g2[19][30] , \g2[19][29] , 
        \g2[19][28] , \g2[19][27] , \g2[19][26] , \g2[19][25] , \g2[19][24] , 
        \g2[19][23] , \g2[19][22] , \g2[19][21] , \g2[19][20] , \g2[19][19] , 
        \g2[19][18] , \g2[19][17] , \g2[19][16] , \g2[19][15] , \g2[19][14] , 
        \g2[19][13] , \g2[19][12] , \g2[19][11] , \g2[19][10] , \g2[19][9] , 
        \g2[19][8] , \g2[19][7] , \g2[19][6] , \g2[19][5] , \g2[19][4] , 
        \g2[19][3] , \g2[19][2] , \g2[19][1] , 1'b0}), .cin({\g2[20][63] , 
        \g2[20][62] , \g2[20][61] , \g2[20][60] , \g2[20][59] , \g2[20][58] , 
        \g2[20][57] , \g2[20][56] , \g2[20][55] , \g2[20][54] , \g2[20][53] , 
        \g2[20][52] , \g2[20][51] , \g2[20][50] , \g2[20][49] , \g2[20][48] , 
        \g2[20][47] , \g2[20][46] , \g2[20][45] , \g2[20][44] , \g2[20][43] , 
        \g2[20][42] , \g2[20][41] , \g2[20][40] , \g2[20][39] , \g2[20][38] , 
        \g2[20][37] , \g2[20][36] , \g2[20][35] , \g2[20][34] , \g2[20][33] , 
        \g2[20][32] , \g2[20][31] , \g2[20][30] , \g2[20][29] , \g2[20][28] , 
        \g2[20][27] , \g2[20][26] , \g2[20][25] , \g2[20][24] , \g2[20][23] , 
        \g2[20][22] , \g2[20][21] , \g2[20][20] , \g2[20][19] , \g2[20][18] , 
        \g2[20][17] , \g2[20][16] , \g2[20][15] , \g2[20][14] , \g2[20][13] , 
        \g2[20][12] , \g2[20][11] , \g2[20][10] , \g2[20][9] , \g2[20][8] , 
        \g2[20][7] , \g2[20][6] , \g2[20][5] , \g2[20][4] , \g2[20][3] , 
        \g2[20][2] , \g2[20][1] , 1'b0}), .sum({\g3[6][63] , \g3[6][62] , 
        \g3[6][61] , \g3[6][60] , \g3[6][59] , \g3[6][58] , \g3[6][57] , 
        \g3[6][56] , \g3[6][55] , \g3[6][54] , \g3[6][53] , \g3[6][52] , 
        \g3[6][51] , \g3[6][50] , \g3[6][49] , \g3[6][48] , \g3[6][47] , 
        \g3[6][46] , \g3[6][45] , \g3[6][44] , \g3[6][43] , \g3[6][42] , 
        \g3[6][41] , \g3[6][40] , \g3[6][39] , \g3[6][38] , \g3[6][37] , 
        \g3[6][36] , \g3[6][35] , \g3[6][34] , \g3[6][33] , \g3[6][32] , 
        \g3[6][31] , \g3[6][30] , \g3[6][29] , \g3[6][28] , \g3[6][27] , 
        \g3[6][26] , \g3[6][25] , \g3[6][24] , \g3[6][23] , \g3[6][22] , 
        \g3[6][21] , \g3[6][20] , \g3[6][19] , \g3[6][18] , \g3[6][17] , 
        \g3[6][16] , \g3[6][15] , \g3[6][14] , \g3[6][13] , \g3[6][12] , 
        \g3[6][11] , \g3[6][10] , \g3[6][9] , \g3[6][8] , \g3[6][7] , 
        \g3[6][6] , \g3[6][5] , \g3[6][4] , \g3[6][3] , \g3[6][2] , \g3[6][1] , 
        \g3[6][0] }), .cout({\g3[15][63] , \g3[15][62] , \g3[15][61] , 
        \g3[15][60] , \g3[15][59] , \g3[15][58] , \g3[15][57] , \g3[15][56] , 
        \g3[15][55] , \g3[15][54] , \g3[15][53] , \g3[15][52] , \g3[15][51] , 
        \g3[15][50] , \g3[15][49] , \g3[15][48] , \g3[15][47] , \g3[15][46] , 
        \g3[15][45] , \g3[15][44] , \g3[15][43] , \g3[15][42] , \g3[15][41] , 
        \g3[15][40] , \g3[15][39] , \g3[15][38] , \g3[15][37] , \g3[15][36] , 
        \g3[15][35] , \g3[15][34] , \g3[15][33] , \g3[15][32] , \g3[15][31] , 
        \g3[15][30] , \g3[15][29] , \g3[15][28] , \g3[15][27] , \g3[15][26] , 
        \g3[15][25] , \g3[15][24] , \g3[15][23] , \g3[15][22] , \g3[15][21] , 
        \g3[15][20] , \g3[15][19] , \g3[15][18] , \g3[15][17] , \g3[15][16] , 
        \g3[15][15] , \g3[15][14] , \g3[15][13] , \g3[15][12] , \g3[15][11] , 
        \g3[15][10] , \g3[15][9] , \g3[15][8] , \g3[15][7] , \g3[15][6] , 
        \g3[15][5] , \g3[15][4] , \g3[15][3] , \g3[15][2] , \g3[15][1] , 
        SYNOPSYS_UNCONNECTED__41}) );
  FullAdder \level3[7].x0  ( .a({\g2[21][63] , \g2[21][62] , \g2[21][61] , 
        \g2[21][60] , \g2[21][59] , \g2[21][58] , \g2[21][57] , \g2[21][56] , 
        \g2[21][55] , \g2[21][54] , \g2[21][53] , \g2[21][52] , \g2[21][51] , 
        \g2[21][50] , \g2[21][49] , \g2[21][48] , \g2[21][47] , \g2[21][46] , 
        \g2[21][45] , \g2[21][44] , \g2[21][43] , \g2[21][42] , \g2[21][41] , 
        \g2[21][40] , \g2[21][39] , \g2[21][38] , \g2[21][37] , \g2[21][36] , 
        \g2[21][35] , \g2[21][34] , \g2[21][33] , \g2[21][32] , \g2[21][31] , 
        \g2[21][30] , \g2[21][29] , \g2[21][28] , \g2[21][27] , \g2[21][26] , 
        \g2[21][25] , \g2[21][24] , \g2[21][23] , \g2[21][22] , \g2[21][21] , 
        \g2[21][20] , \g2[21][19] , \g2[21][18] , \g2[21][17] , \g2[21][16] , 
        \g2[21][15] , \g2[21][14] , \g2[21][13] , \g2[21][12] , \g2[21][11] , 
        \g2[21][10] , \g2[21][9] , \g2[21][8] , \g2[21][7] , \g2[21][6] , 
        \g2[21][5] , \g2[21][4] , \g2[21][3] , \g2[21][2] , \g2[21][1] , 1'b0}), .b({\g2[22][63] , \g2[22][62] , \g2[22][61] , \g2[22][60] , \g2[22][59] , 
        \g2[22][58] , \g2[22][57] , \g2[22][56] , \g2[22][55] , \g2[22][54] , 
        \g2[22][53] , \g2[22][52] , \g2[22][51] , \g2[22][50] , \g2[22][49] , 
        \g2[22][48] , \g2[22][47] , \g2[22][46] , \g2[22][45] , \g2[22][44] , 
        \g2[22][43] , \g2[22][42] , \g2[22][41] , \g2[22][40] , \g2[22][39] , 
        \g2[22][38] , \g2[22][37] , \g2[22][36] , \g2[22][35] , \g2[22][34] , 
        \g2[22][33] , \g2[22][32] , \g2[22][31] , \g2[22][30] , \g2[22][29] , 
        \g2[22][28] , \g2[22][27] , \g2[22][26] , \g2[22][25] , \g2[22][24] , 
        \g2[22][23] , \g2[22][22] , \g2[22][21] , \g2[22][20] , \g2[22][19] , 
        \g2[22][18] , \g2[22][17] , \g2[22][16] , \g2[22][15] , \g2[22][14] , 
        \g2[22][13] , \g2[22][12] , \g2[22][11] , \g2[22][10] , \g2[22][9] , 
        \g2[22][8] , \g2[22][7] , \g2[22][6] , \g2[22][5] , \g2[22][4] , 
        \g2[22][3] , \g2[22][2] , \g2[22][1] , 1'b0}), .cin({\g2[23][63] , 
        \g2[23][62] , \g2[23][61] , \g2[23][60] , \g2[23][59] , \g2[23][58] , 
        \g2[23][57] , \g2[23][56] , \g2[23][55] , \g2[23][54] , \g2[23][53] , 
        \g2[23][52] , \g2[23][51] , \g2[23][50] , \g2[23][49] , \g2[23][48] , 
        \g2[23][47] , \g2[23][46] , \g2[23][45] , \g2[23][44] , \g2[23][43] , 
        \g2[23][42] , \g2[23][41] , \g2[23][40] , \g2[23][39] , \g2[23][38] , 
        \g2[23][37] , \g2[23][36] , \g2[23][35] , \g2[23][34] , \g2[23][33] , 
        \g2[23][32] , \g2[23][31] , \g2[23][30] , \g2[23][29] , \g2[23][28] , 
        \g2[23][27] , \g2[23][26] , \g2[23][25] , \g2[23][24] , \g2[23][23] , 
        \g2[23][22] , \g2[23][21] , \g2[23][20] , \g2[23][19] , \g2[23][18] , 
        \g2[23][17] , \g2[23][16] , \g2[23][15] , \g2[23][14] , \g2[23][13] , 
        \g2[23][12] , \g2[23][11] , \g2[23][10] , \g2[23][9] , \g2[23][8] , 
        \g2[23][7] , \g2[23][6] , \g2[23][5] , \g2[23][4] , \g2[23][3] , 
        \g2[23][2] , \g2[23][1] , 1'b0}), .sum({\g3[7][63] , \g3[7][62] , 
        \g3[7][61] , \g3[7][60] , \g3[7][59] , \g3[7][58] , \g3[7][57] , 
        \g3[7][56] , \g3[7][55] , \g3[7][54] , \g3[7][53] , \g3[7][52] , 
        \g3[7][51] , \g3[7][50] , \g3[7][49] , \g3[7][48] , \g3[7][47] , 
        \g3[7][46] , \g3[7][45] , \g3[7][44] , \g3[7][43] , \g3[7][42] , 
        \g3[7][41] , \g3[7][40] , \g3[7][39] , \g3[7][38] , \g3[7][37] , 
        \g3[7][36] , \g3[7][35] , \g3[7][34] , \g3[7][33] , \g3[7][32] , 
        \g3[7][31] , \g3[7][30] , \g3[7][29] , \g3[7][28] , \g3[7][27] , 
        \g3[7][26] , \g3[7][25] , \g3[7][24] , \g3[7][23] , \g3[7][22] , 
        \g3[7][21] , \g3[7][20] , \g3[7][19] , \g3[7][18] , \g3[7][17] , 
        \g3[7][16] , \g3[7][15] , \g3[7][14] , \g3[7][13] , \g3[7][12] , 
        \g3[7][11] , \g3[7][10] , \g3[7][9] , \g3[7][8] , \g3[7][7] , 
        \g3[7][6] , \g3[7][5] , \g3[7][4] , \g3[7][3] , \g3[7][2] , \g3[7][1] , 
        \g3[7][0] }), .cout({\g3[16][63] , \g3[16][62] , \g3[16][61] , 
        \g3[16][60] , \g3[16][59] , \g3[16][58] , \g3[16][57] , \g3[16][56] , 
        \g3[16][55] , \g3[16][54] , \g3[16][53] , \g3[16][52] , \g3[16][51] , 
        \g3[16][50] , \g3[16][49] , \g3[16][48] , \g3[16][47] , \g3[16][46] , 
        \g3[16][45] , \g3[16][44] , \g3[16][43] , \g3[16][42] , \g3[16][41] , 
        \g3[16][40] , \g3[16][39] , \g3[16][38] , \g3[16][37] , \g3[16][36] , 
        \g3[16][35] , \g3[16][34] , \g3[16][33] , \g3[16][32] , \g3[16][31] , 
        \g3[16][30] , \g3[16][29] , \g3[16][28] , \g3[16][27] , \g3[16][26] , 
        \g3[16][25] , \g3[16][24] , \g3[16][23] , \g3[16][22] , \g3[16][21] , 
        \g3[16][20] , \g3[16][19] , \g3[16][18] , \g3[16][17] , \g3[16][16] , 
        \g3[16][15] , \g3[16][14] , \g3[16][13] , \g3[16][12] , \g3[16][11] , 
        \g3[16][10] , \g3[16][9] , \g3[16][8] , \g3[16][7] , \g3[16][6] , 
        \g3[16][5] , \g3[16][4] , \g3[16][3] , \g3[16][2] , \g3[16][1] , 
        SYNOPSYS_UNCONNECTED__42}) );
  FullAdder \level3[8].x0  ( .a({\g2[24][63] , \g2[24][62] , \g2[24][61] , 
        \g2[24][60] , \g2[24][59] , \g2[24][58] , \g2[24][57] , \g2[24][56] , 
        \g2[24][55] , \g2[24][54] , \g2[24][53] , \g2[24][52] , \g2[24][51] , 
        \g2[24][50] , \g2[24][49] , \g2[24][48] , \g2[24][47] , \g2[24][46] , 
        \g2[24][45] , \g2[24][44] , \g2[24][43] , \g2[24][42] , \g2[24][41] , 
        \g2[24][40] , \g2[24][39] , \g2[24][38] , \g2[24][37] , \g2[24][36] , 
        \g2[24][35] , \g2[24][34] , \g2[24][33] , \g2[24][32] , \g2[24][31] , 
        \g2[24][30] , \g2[24][29] , \g2[24][28] , \g2[24][27] , \g2[24][26] , 
        \g2[24][25] , \g2[24][24] , \g2[24][23] , \g2[24][22] , \g2[24][21] , 
        \g2[24][20] , \g2[24][19] , \g2[24][18] , \g2[24][17] , \g2[24][16] , 
        \g2[24][15] , \g2[24][14] , \g2[24][13] , \g2[24][12] , \g2[24][11] , 
        \g2[24][10] , \g2[24][9] , \g2[24][8] , \g2[24][7] , \g2[24][6] , 
        \g2[24][5] , \g2[24][4] , \g2[24][3] , \g2[24][2] , \g2[24][1] , 1'b0}), .b({\g2[25][63] , \g2[25][62] , \g2[25][61] , \g2[25][60] , \g2[25][59] , 
        \g2[25][58] , \g2[25][57] , \g2[25][56] , \g2[25][55] , \g2[25][54] , 
        \g2[25][53] , \g2[25][52] , \g2[25][51] , \g2[25][50] , \g2[25][49] , 
        \g2[25][48] , \g2[25][47] , \g2[25][46] , \g2[25][45] , \g2[25][44] , 
        \g2[25][43] , \g2[25][42] , \g2[25][41] , \g2[25][40] , \g2[25][39] , 
        \g2[25][38] , \g2[25][37] , \g2[25][36] , \g2[25][35] , \g2[25][34] , 
        \g2[25][33] , \g2[25][32] , \g2[25][31] , \g2[25][30] , \g2[25][29] , 
        \g2[25][28] , \g2[25][27] , \g2[25][26] , \g2[25][25] , \g2[25][24] , 
        \g2[25][23] , \g2[25][22] , \g2[25][21] , \g2[25][20] , \g2[25][19] , 
        \g2[25][18] , \g2[25][17] , \g2[25][16] , \g2[25][15] , \g2[25][14] , 
        \g2[25][13] , \g2[25][12] , \g2[25][11] , \g2[25][10] , \g2[25][9] , 
        \g2[25][8] , \g2[25][7] , \g2[25][6] , \g2[25][5] , \g2[25][4] , 
        \g2[25][3] , \g2[25][2] , \g2[25][1] , 1'b0}), .cin({\g2[26][63] , 
        \g2[26][62] , \g2[26][61] , \g2[26][60] , \g2[26][59] , \g2[26][58] , 
        \g2[26][57] , \g2[26][56] , \g2[26][55] , \g2[26][54] , \g2[26][53] , 
        \g2[26][52] , \g2[26][51] , \g2[26][50] , \g2[26][49] , \g2[26][48] , 
        \g2[26][47] , \g2[26][46] , \g2[26][45] , \g2[26][44] , \g2[26][43] , 
        \g2[26][42] , \g2[26][41] , \g2[26][40] , \g2[26][39] , \g2[26][38] , 
        \g2[26][37] , \g2[26][36] , \g2[26][35] , \g2[26][34] , \g2[26][33] , 
        \g2[26][32] , \g2[26][31] , \g2[26][30] , \g2[26][29] , \g2[26][28] , 
        \g2[26][27] , \g2[26][26] , \g2[26][25] , \g2[26][24] , \g2[26][23] , 
        \g2[26][22] , \g2[26][21] , \g2[26][20] , \g2[26][19] , \g2[26][18] , 
        \g2[26][17] , \g2[26][16] , \g2[26][15] , \g2[26][14] , \g2[26][13] , 
        \g2[26][12] , \g2[26][11] , \g2[26][10] , \g2[26][9] , \g2[26][8] , 
        \g2[26][7] , \g2[26][6] , \g2[26][5] , \g2[26][4] , \g2[26][3] , 
        \g2[26][2] , \g2[26][1] , 1'b0}), .sum({\g3[8][63] , \g3[8][62] , 
        \g3[8][61] , \g3[8][60] , \g3[8][59] , \g3[8][58] , \g3[8][57] , 
        \g3[8][56] , \g3[8][55] , \g3[8][54] , \g3[8][53] , \g3[8][52] , 
        \g3[8][51] , \g3[8][50] , \g3[8][49] , \g3[8][48] , \g3[8][47] , 
        \g3[8][46] , \g3[8][45] , \g3[8][44] , \g3[8][43] , \g3[8][42] , 
        \g3[8][41] , \g3[8][40] , \g3[8][39] , \g3[8][38] , \g3[8][37] , 
        \g3[8][36] , \g3[8][35] , \g3[8][34] , \g3[8][33] , \g3[8][32] , 
        \g3[8][31] , \g3[8][30] , \g3[8][29] , \g3[8][28] , \g3[8][27] , 
        \g3[8][26] , \g3[8][25] , \g3[8][24] , \g3[8][23] , \g3[8][22] , 
        \g3[8][21] , \g3[8][20] , \g3[8][19] , \g3[8][18] , \g3[8][17] , 
        \g3[8][16] , \g3[8][15] , \g3[8][14] , \g3[8][13] , \g3[8][12] , 
        \g3[8][11] , \g3[8][10] , \g3[8][9] , \g3[8][8] , \g3[8][7] , 
        \g3[8][6] , \g3[8][5] , \g3[8][4] , \g3[8][3] , \g3[8][2] , \g3[8][1] , 
        \g3[8][0] }), .cout({\g3[17][63] , \g3[17][62] , \g3[17][61] , 
        \g3[17][60] , \g3[17][59] , \g3[17][58] , \g3[17][57] , \g3[17][56] , 
        \g3[17][55] , \g3[17][54] , \g3[17][53] , \g3[17][52] , \g3[17][51] , 
        \g3[17][50] , \g3[17][49] , \g3[17][48] , \g3[17][47] , \g3[17][46] , 
        \g3[17][45] , \g3[17][44] , \g3[17][43] , \g3[17][42] , \g3[17][41] , 
        \g3[17][40] , \g3[17][39] , \g3[17][38] , \g3[17][37] , \g3[17][36] , 
        \g3[17][35] , \g3[17][34] , \g3[17][33] , \g3[17][32] , \g3[17][31] , 
        \g3[17][30] , \g3[17][29] , \g3[17][28] , \g3[17][27] , \g3[17][26] , 
        \g3[17][25] , \g3[17][24] , \g3[17][23] , \g3[17][22] , \g3[17][21] , 
        \g3[17][20] , \g3[17][19] , \g3[17][18] , \g3[17][17] , \g3[17][16] , 
        \g3[17][15] , \g3[17][14] , \g3[17][13] , \g3[17][12] , \g3[17][11] , 
        \g3[17][10] , \g3[17][9] , \g3[17][8] , \g3[17][7] , \g3[17][6] , 
        \g3[17][5] , \g3[17][4] , \g3[17][3] , \g3[17][2] , \g3[17][1] , 
        SYNOPSYS_UNCONNECTED__43}) );
  FullAdder \level4[0].x1  ( .a({\g3[0][63] , \g3[0][62] , \g3[0][61] , 
        \g3[0][60] , \g3[0][59] , \g3[0][58] , \g3[0][57] , \g3[0][56] , 
        \g3[0][55] , \g3[0][54] , \g3[0][53] , \g3[0][52] , \g3[0][51] , 
        \g3[0][50] , \g3[0][49] , \g3[0][48] , \g3[0][47] , \g3[0][46] , 
        \g3[0][45] , \g3[0][44] , \g3[0][43] , \g3[0][42] , \g3[0][41] , 
        \g3[0][40] , \g3[0][39] , \g3[0][38] , \g3[0][37] , \g3[0][36] , 
        \g3[0][35] , \g3[0][34] , \g3[0][33] , \g3[0][32] , \g3[0][31] , 
        \g3[0][30] , \g3[0][29] , \g3[0][28] , \g3[0][27] , \g3[0][26] , 
        \g3[0][25] , \g3[0][24] , \g3[0][23] , \g3[0][22] , \g3[0][21] , 
        \g3[0][20] , \g3[0][19] , \g3[0][18] , \g3[0][17] , \g3[0][16] , 
        \g3[0][15] , \g3[0][14] , \g3[0][13] , \g3[0][12] , \g3[0][11] , 
        \g3[0][10] , \g3[0][9] , \g3[0][8] , \g3[0][7] , \g3[0][6] , 
        \g3[0][5] , \g3[0][4] , \g3[0][3] , \g3[0][2] , \g3[0][1] , \g3[0][0] }), .b({\g3[1][63] , \g3[1][62] , \g3[1][61] , \g3[1][60] , \g3[1][59] , 
        \g3[1][58] , \g3[1][57] , \g3[1][56] , \g3[1][55] , \g3[1][54] , 
        \g3[1][53] , \g3[1][52] , \g3[1][51] , \g3[1][50] , \g3[1][49] , 
        \g3[1][48] , \g3[1][47] , \g3[1][46] , \g3[1][45] , \g3[1][44] , 
        \g3[1][43] , \g3[1][42] , \g3[1][41] , \g3[1][40] , \g3[1][39] , 
        \g3[1][38] , \g3[1][37] , \g3[1][36] , \g3[1][35] , \g3[1][34] , 
        \g3[1][33] , \g3[1][32] , \g3[1][31] , \g3[1][30] , \g3[1][29] , 
        \g3[1][28] , \g3[1][27] , \g3[1][26] , \g3[1][25] , \g3[1][24] , 
        \g3[1][23] , \g3[1][22] , \g3[1][21] , \g3[1][20] , \g3[1][19] , 
        \g3[1][18] , \g3[1][17] , \g3[1][16] , \g3[1][15] , \g3[1][14] , 
        \g3[1][13] , \g3[1][12] , \g3[1][11] , \g3[1][10] , \g3[1][9] , 
        \g3[1][8] , \g3[1][7] , \g3[1][6] , \g3[1][5] , \g3[1][4] , \g3[1][3] , 
        \g3[1][2] , \g3[1][1] , \g3[1][0] }), .cin({\g3[2][63] , \g3[2][62] , 
        \g3[2][61] , \g3[2][60] , \g3[2][59] , \g3[2][58] , \g3[2][57] , 
        \g3[2][56] , \g3[2][55] , \g3[2][54] , \g3[2][53] , \g3[2][52] , 
        \g3[2][51] , \g3[2][50] , \g3[2][49] , \g3[2][48] , \g3[2][47] , 
        \g3[2][46] , \g3[2][45] , \g3[2][44] , \g3[2][43] , \g3[2][42] , 
        \g3[2][41] , \g3[2][40] , \g3[2][39] , \g3[2][38] , \g3[2][37] , 
        \g3[2][36] , \g3[2][35] , \g3[2][34] , \g3[2][33] , \g3[2][32] , 
        \g3[2][31] , \g3[2][30] , \g3[2][29] , \g3[2][28] , \g3[2][27] , 
        \g3[2][26] , \g3[2][25] , \g3[2][24] , \g3[2][23] , \g3[2][22] , 
        \g3[2][21] , \g3[2][20] , \g3[2][19] , \g3[2][18] , \g3[2][17] , 
        \g3[2][16] , \g3[2][15] , \g3[2][14] , \g3[2][13] , \g3[2][12] , 
        \g3[2][11] , \g3[2][10] , \g3[2][9] , \g3[2][8] , \g3[2][7] , 
        \g3[2][6] , \g3[2][5] , \g3[2][4] , \g3[2][3] , \g3[2][2] , \g3[2][1] , 
        \g3[2][0] }), .sum({\g4[0][63] , \g4[0][62] , \g4[0][61] , \g4[0][60] , 
        \g4[0][59] , \g4[0][58] , \g4[0][57] , \g4[0][56] , \g4[0][55] , 
        \g4[0][54] , \g4[0][53] , \g4[0][52] , \g4[0][51] , \g4[0][50] , 
        \g4[0][49] , \g4[0][48] , \g4[0][47] , \g4[0][46] , \g4[0][45] , 
        \g4[0][44] , \g4[0][43] , \g4[0][42] , \g4[0][41] , \g4[0][40] , 
        \g4[0][39] , \g4[0][38] , \g4[0][37] , \g4[0][36] , \g4[0][35] , 
        \g4[0][34] , \g4[0][33] , \g4[0][32] , \g4[0][31] , \g4[0][30] , 
        \g4[0][29] , \g4[0][28] , \g4[0][27] , \g4[0][26] , \g4[0][25] , 
        \g4[0][24] , \g4[0][23] , \g4[0][22] , \g4[0][21] , \g4[0][20] , 
        \g4[0][19] , \g4[0][18] , \g4[0][17] , \g4[0][16] , \g4[0][15] , 
        \g4[0][14] , \g4[0][13] , \g4[0][12] , \g4[0][11] , \g4[0][10] , 
        \g4[0][9] , \g4[0][8] , \g4[0][7] , \g4[0][6] , \g4[0][5] , \g4[0][4] , 
        \g4[0][3] , \g4[0][2] , \g4[0][1] , \g4[0][0] }), .cout({\g4[6][63] , 
        \g4[6][62] , \g4[6][61] , \g4[6][60] , \g4[6][59] , \g4[6][58] , 
        \g4[6][57] , \g4[6][56] , \g4[6][55] , \g4[6][54] , \g4[6][53] , 
        \g4[6][52] , \g4[6][51] , \g4[6][50] , \g4[6][49] , \g4[6][48] , 
        \g4[6][47] , \g4[6][46] , \g4[6][45] , \g4[6][44] , \g4[6][43] , 
        \g4[6][42] , \g4[6][41] , \g4[6][40] , \g4[6][39] , \g4[6][38] , 
        \g4[6][37] , \g4[6][36] , \g4[6][35] , \g4[6][34] , \g4[6][33] , 
        \g4[6][32] , \g4[6][31] , \g4[6][30] , \g4[6][29] , \g4[6][28] , 
        \g4[6][27] , \g4[6][26] , \g4[6][25] , \g4[6][24] , \g4[6][23] , 
        \g4[6][22] , \g4[6][21] , \g4[6][20] , \g4[6][19] , \g4[6][18] , 
        \g4[6][17] , \g4[6][16] , \g4[6][15] , \g4[6][14] , \g4[6][13] , 
        \g4[6][12] , \g4[6][11] , \g4[6][10] , \g4[6][9] , \g4[6][8] , 
        \g4[6][7] , \g4[6][6] , \g4[6][5] , \g4[6][4] , \g4[6][3] , \g4[6][2] , 
        \g4[6][1] , SYNOPSYS_UNCONNECTED__44}) );
  FullAdder \level4[1].x1  ( .a({\g3[3][63] , \g3[3][62] , \g3[3][61] , 
        \g3[3][60] , \g3[3][59] , \g3[3][58] , \g3[3][57] , \g3[3][56] , 
        \g3[3][55] , \g3[3][54] , \g3[3][53] , \g3[3][52] , \g3[3][51] , 
        \g3[3][50] , \g3[3][49] , \g3[3][48] , \g3[3][47] , \g3[3][46] , 
        \g3[3][45] , \g3[3][44] , \g3[3][43] , \g3[3][42] , \g3[3][41] , 
        \g3[3][40] , \g3[3][39] , \g3[3][38] , \g3[3][37] , \g3[3][36] , 
        \g3[3][35] , \g3[3][34] , \g3[3][33] , \g3[3][32] , \g3[3][31] , 
        \g3[3][30] , \g3[3][29] , \g3[3][28] , \g3[3][27] , \g3[3][26] , 
        \g3[3][25] , \g3[3][24] , \g3[3][23] , \g3[3][22] , \g3[3][21] , 
        \g3[3][20] , \g3[3][19] , \g3[3][18] , \g3[3][17] , \g3[3][16] , 
        \g3[3][15] , \g3[3][14] , \g3[3][13] , \g3[3][12] , \g3[3][11] , 
        \g3[3][10] , \g3[3][9] , \g3[3][8] , \g3[3][7] , \g3[3][6] , 
        \g3[3][5] , \g3[3][4] , \g3[3][3] , \g3[3][2] , \g3[3][1] , \g3[3][0] }), .b({\g3[4][63] , \g3[4][62] , \g3[4][61] , \g3[4][60] , \g3[4][59] , 
        \g3[4][58] , \g3[4][57] , \g3[4][56] , \g3[4][55] , \g3[4][54] , 
        \g3[4][53] , \g3[4][52] , \g3[4][51] , \g3[4][50] , \g3[4][49] , 
        \g3[4][48] , \g3[4][47] , \g3[4][46] , \g3[4][45] , \g3[4][44] , 
        \g3[4][43] , \g3[4][42] , \g3[4][41] , \g3[4][40] , \g3[4][39] , 
        \g3[4][38] , \g3[4][37] , \g3[4][36] , \g3[4][35] , \g3[4][34] , 
        \g3[4][33] , \g3[4][32] , \g3[4][31] , \g3[4][30] , \g3[4][29] , 
        \g3[4][28] , \g3[4][27] , \g3[4][26] , \g3[4][25] , \g3[4][24] , 
        \g3[4][23] , \g3[4][22] , \g3[4][21] , \g3[4][20] , \g3[4][19] , 
        \g3[4][18] , \g3[4][17] , \g3[4][16] , \g3[4][15] , \g3[4][14] , 
        \g3[4][13] , \g3[4][12] , \g3[4][11] , \g3[4][10] , \g3[4][9] , 
        \g3[4][8] , \g3[4][7] , \g3[4][6] , \g3[4][5] , \g3[4][4] , \g3[4][3] , 
        \g3[4][2] , \g3[4][1] , \g3[4][0] }), .cin({\g3[5][63] , \g3[5][62] , 
        \g3[5][61] , \g3[5][60] , \g3[5][59] , \g3[5][58] , \g3[5][57] , 
        \g3[5][56] , \g3[5][55] , \g3[5][54] , \g3[5][53] , \g3[5][52] , 
        \g3[5][51] , \g3[5][50] , \g3[5][49] , \g3[5][48] , \g3[5][47] , 
        \g3[5][46] , \g3[5][45] , \g3[5][44] , \g3[5][43] , \g3[5][42] , 
        \g3[5][41] , \g3[5][40] , \g3[5][39] , \g3[5][38] , \g3[5][37] , 
        \g3[5][36] , \g3[5][35] , \g3[5][34] , \g3[5][33] , \g3[5][32] , 
        \g3[5][31] , \g3[5][30] , \g3[5][29] , \g3[5][28] , \g3[5][27] , 
        \g3[5][26] , \g3[5][25] , \g3[5][24] , \g3[5][23] , \g3[5][22] , 
        \g3[5][21] , \g3[5][20] , \g3[5][19] , \g3[5][18] , \g3[5][17] , 
        \g3[5][16] , \g3[5][15] , \g3[5][14] , \g3[5][13] , \g3[5][12] , 
        \g3[5][11] , \g3[5][10] , \g3[5][9] , \g3[5][8] , \g3[5][7] , 
        \g3[5][6] , \g3[5][5] , \g3[5][4] , \g3[5][3] , \g3[5][2] , \g3[5][1] , 
        \g3[5][0] }), .sum({\g4[1][63] , \g4[1][62] , \g4[1][61] , \g4[1][60] , 
        \g4[1][59] , \g4[1][58] , \g4[1][57] , \g4[1][56] , \g4[1][55] , 
        \g4[1][54] , \g4[1][53] , \g4[1][52] , \g4[1][51] , \g4[1][50] , 
        \g4[1][49] , \g4[1][48] , \g4[1][47] , \g4[1][46] , \g4[1][45] , 
        \g4[1][44] , \g4[1][43] , \g4[1][42] , \g4[1][41] , \g4[1][40] , 
        \g4[1][39] , \g4[1][38] , \g4[1][37] , \g4[1][36] , \g4[1][35] , 
        \g4[1][34] , \g4[1][33] , \g4[1][32] , \g4[1][31] , \g4[1][30] , 
        \g4[1][29] , \g4[1][28] , \g4[1][27] , \g4[1][26] , \g4[1][25] , 
        \g4[1][24] , \g4[1][23] , \g4[1][22] , \g4[1][21] , \g4[1][20] , 
        \g4[1][19] , \g4[1][18] , \g4[1][17] , \g4[1][16] , \g4[1][15] , 
        \g4[1][14] , \g4[1][13] , \g4[1][12] , \g4[1][11] , \g4[1][10] , 
        \g4[1][9] , \g4[1][8] , \g4[1][7] , \g4[1][6] , \g4[1][5] , \g4[1][4] , 
        \g4[1][3] , \g4[1][2] , \g4[1][1] , \g4[1][0] }), .cout({\g4[7][63] , 
        \g4[7][62] , \g4[7][61] , \g4[7][60] , \g4[7][59] , \g4[7][58] , 
        \g4[7][57] , \g4[7][56] , \g4[7][55] , \g4[7][54] , \g4[7][53] , 
        \g4[7][52] , \g4[7][51] , \g4[7][50] , \g4[7][49] , \g4[7][48] , 
        \g4[7][47] , \g4[7][46] , \g4[7][45] , \g4[7][44] , \g4[7][43] , 
        \g4[7][42] , \g4[7][41] , \g4[7][40] , \g4[7][39] , \g4[7][38] , 
        \g4[7][37] , \g4[7][36] , \g4[7][35] , \g4[7][34] , \g4[7][33] , 
        \g4[7][32] , \g4[7][31] , \g4[7][30] , \g4[7][29] , \g4[7][28] , 
        \g4[7][27] , \g4[7][26] , \g4[7][25] , \g4[7][24] , \g4[7][23] , 
        \g4[7][22] , \g4[7][21] , \g4[7][20] , \g4[7][19] , \g4[7][18] , 
        \g4[7][17] , \g4[7][16] , \g4[7][15] , \g4[7][14] , \g4[7][13] , 
        \g4[7][12] , \g4[7][11] , \g4[7][10] , \g4[7][9] , \g4[7][8] , 
        \g4[7][7] , \g4[7][6] , \g4[7][5] , \g4[7][4] , \g4[7][3] , \g4[7][2] , 
        \g4[7][1] , SYNOPSYS_UNCONNECTED__45}) );
  FullAdder \level4[2].x1  ( .a({\g3[6][63] , \g3[6][62] , \g3[6][61] , 
        \g3[6][60] , \g3[6][59] , \g3[6][58] , \g3[6][57] , \g3[6][56] , 
        \g3[6][55] , \g3[6][54] , \g3[6][53] , \g3[6][52] , \g3[6][51] , 
        \g3[6][50] , \g3[6][49] , \g3[6][48] , \g3[6][47] , \g3[6][46] , 
        \g3[6][45] , \g3[6][44] , \g3[6][43] , \g3[6][42] , \g3[6][41] , 
        \g3[6][40] , \g3[6][39] , \g3[6][38] , \g3[6][37] , \g3[6][36] , 
        \g3[6][35] , \g3[6][34] , \g3[6][33] , \g3[6][32] , \g3[6][31] , 
        \g3[6][30] , \g3[6][29] , \g3[6][28] , \g3[6][27] , \g3[6][26] , 
        \g3[6][25] , \g3[6][24] , \g3[6][23] , \g3[6][22] , \g3[6][21] , 
        \g3[6][20] , \g3[6][19] , \g3[6][18] , \g3[6][17] , \g3[6][16] , 
        \g3[6][15] , \g3[6][14] , \g3[6][13] , \g3[6][12] , \g3[6][11] , 
        \g3[6][10] , \g3[6][9] , \g3[6][8] , \g3[6][7] , \g3[6][6] , 
        \g3[6][5] , \g3[6][4] , \g3[6][3] , \g3[6][2] , \g3[6][1] , \g3[6][0] }), .b({\g3[7][63] , \g3[7][62] , \g3[7][61] , \g3[7][60] , \g3[7][59] , 
        \g3[7][58] , \g3[7][57] , \g3[7][56] , \g3[7][55] , \g3[7][54] , 
        \g3[7][53] , \g3[7][52] , \g3[7][51] , \g3[7][50] , \g3[7][49] , 
        \g3[7][48] , \g3[7][47] , \g3[7][46] , \g3[7][45] , \g3[7][44] , 
        \g3[7][43] , \g3[7][42] , \g3[7][41] , \g3[7][40] , \g3[7][39] , 
        \g3[7][38] , \g3[7][37] , \g3[7][36] , \g3[7][35] , \g3[7][34] , 
        \g3[7][33] , \g3[7][32] , \g3[7][31] , \g3[7][30] , \g3[7][29] , 
        \g3[7][28] , \g3[7][27] , \g3[7][26] , \g3[7][25] , \g3[7][24] , 
        \g3[7][23] , \g3[7][22] , \g3[7][21] , \g3[7][20] , \g3[7][19] , 
        \g3[7][18] , \g3[7][17] , \g3[7][16] , \g3[7][15] , \g3[7][14] , 
        \g3[7][13] , \g3[7][12] , \g3[7][11] , \g3[7][10] , \g3[7][9] , 
        \g3[7][8] , \g3[7][7] , \g3[7][6] , \g3[7][5] , \g3[7][4] , \g3[7][3] , 
        \g3[7][2] , \g3[7][1] , \g3[7][0] }), .cin({\g3[8][63] , \g3[8][62] , 
        \g3[8][61] , \g3[8][60] , \g3[8][59] , \g3[8][58] , \g3[8][57] , 
        \g3[8][56] , \g3[8][55] , \g3[8][54] , \g3[8][53] , \g3[8][52] , 
        \g3[8][51] , \g3[8][50] , \g3[8][49] , \g3[8][48] , \g3[8][47] , 
        \g3[8][46] , \g3[8][45] , \g3[8][44] , \g3[8][43] , \g3[8][42] , 
        \g3[8][41] , \g3[8][40] , \g3[8][39] , \g3[8][38] , \g3[8][37] , 
        \g3[8][36] , \g3[8][35] , \g3[8][34] , \g3[8][33] , \g3[8][32] , 
        \g3[8][31] , \g3[8][30] , \g3[8][29] , \g3[8][28] , \g3[8][27] , 
        \g3[8][26] , \g3[8][25] , \g3[8][24] , \g3[8][23] , \g3[8][22] , 
        \g3[8][21] , \g3[8][20] , \g3[8][19] , \g3[8][18] , \g3[8][17] , 
        \g3[8][16] , \g3[8][15] , \g3[8][14] , \g3[8][13] , \g3[8][12] , 
        \g3[8][11] , \g3[8][10] , \g3[8][9] , \g3[8][8] , \g3[8][7] , 
        \g3[8][6] , \g3[8][5] , \g3[8][4] , \g3[8][3] , \g3[8][2] , \g3[8][1] , 
        \g3[8][0] }), .sum({\g4[2][63] , \g4[2][62] , \g4[2][61] , \g4[2][60] , 
        \g4[2][59] , \g4[2][58] , \g4[2][57] , \g4[2][56] , \g4[2][55] , 
        \g4[2][54] , \g4[2][53] , \g4[2][52] , \g4[2][51] , \g4[2][50] , 
        \g4[2][49] , \g4[2][48] , \g4[2][47] , \g4[2][46] , \g4[2][45] , 
        \g4[2][44] , \g4[2][43] , \g4[2][42] , \g4[2][41] , \g4[2][40] , 
        \g4[2][39] , \g4[2][38] , \g4[2][37] , \g4[2][36] , \g4[2][35] , 
        \g4[2][34] , \g4[2][33] , \g4[2][32] , \g4[2][31] , \g4[2][30] , 
        \g4[2][29] , \g4[2][28] , \g4[2][27] , \g4[2][26] , \g4[2][25] , 
        \g4[2][24] , \g4[2][23] , \g4[2][22] , \g4[2][21] , \g4[2][20] , 
        \g4[2][19] , \g4[2][18] , \g4[2][17] , \g4[2][16] , \g4[2][15] , 
        \g4[2][14] , \g4[2][13] , \g4[2][12] , \g4[2][11] , \g4[2][10] , 
        \g4[2][9] , \g4[2][8] , \g4[2][7] , \g4[2][6] , \g4[2][5] , \g4[2][4] , 
        \g4[2][3] , \g4[2][2] , \g4[2][1] , \g4[2][0] }), .cout({\g4[8][63] , 
        \g4[8][62] , \g4[8][61] , \g4[8][60] , \g4[8][59] , \g4[8][58] , 
        \g4[8][57] , \g4[8][56] , \g4[8][55] , \g4[8][54] , \g4[8][53] , 
        \g4[8][52] , \g4[8][51] , \g4[8][50] , \g4[8][49] , \g4[8][48] , 
        \g4[8][47] , \g4[8][46] , \g4[8][45] , \g4[8][44] , \g4[8][43] , 
        \g4[8][42] , \g4[8][41] , \g4[8][40] , \g4[8][39] , \g4[8][38] , 
        \g4[8][37] , \g4[8][36] , \g4[8][35] , \g4[8][34] , \g4[8][33] , 
        \g4[8][32] , \g4[8][31] , \g4[8][30] , \g4[8][29] , \g4[8][28] , 
        \g4[8][27] , \g4[8][26] , \g4[8][25] , \g4[8][24] , \g4[8][23] , 
        \g4[8][22] , \g4[8][21] , \g4[8][20] , \g4[8][19] , \g4[8][18] , 
        \g4[8][17] , \g4[8][16] , \g4[8][15] , \g4[8][14] , \g4[8][13] , 
        \g4[8][12] , \g4[8][11] , \g4[8][10] , \g4[8][9] , \g4[8][8] , 
        \g4[8][7] , \g4[8][6] , \g4[8][5] , \g4[8][4] , \g4[8][3] , \g4[8][2] , 
        \g4[8][1] , SYNOPSYS_UNCONNECTED__46}) );
  FullAdder \level4[3].x1  ( .a({\g3[9][63] , \g3[9][62] , \g3[9][61] , 
        \g3[9][60] , \g3[9][59] , \g3[9][58] , \g3[9][57] , \g3[9][56] , 
        \g3[9][55] , \g3[9][54] , \g3[9][53] , \g3[9][52] , \g3[9][51] , 
        \g3[9][50] , \g3[9][49] , \g3[9][48] , \g3[9][47] , \g3[9][46] , 
        \g3[9][45] , \g3[9][44] , \g3[9][43] , \g3[9][42] , \g3[9][41] , 
        \g3[9][40] , \g3[9][39] , \g3[9][38] , \g3[9][37] , \g3[9][36] , 
        \g3[9][35] , \g3[9][34] , \g3[9][33] , \g3[9][32] , \g3[9][31] , 
        \g3[9][30] , \g3[9][29] , \g3[9][28] , \g3[9][27] , \g3[9][26] , 
        \g3[9][25] , \g3[9][24] , \g3[9][23] , \g3[9][22] , \g3[9][21] , 
        \g3[9][20] , \g3[9][19] , \g3[9][18] , \g3[9][17] , \g3[9][16] , 
        \g3[9][15] , \g3[9][14] , \g3[9][13] , \g3[9][12] , \g3[9][11] , 
        \g3[9][10] , \g3[9][9] , \g3[9][8] , \g3[9][7] , \g3[9][6] , 
        \g3[9][5] , \g3[9][4] , \g3[9][3] , \g3[9][2] , \g3[9][1] , 1'b0}), 
        .b({\g3[10][63] , \g3[10][62] , \g3[10][61] , \g3[10][60] , 
        \g3[10][59] , \g3[10][58] , \g3[10][57] , \g3[10][56] , \g3[10][55] , 
        \g3[10][54] , \g3[10][53] , \g3[10][52] , \g3[10][51] , \g3[10][50] , 
        \g3[10][49] , \g3[10][48] , \g3[10][47] , \g3[10][46] , \g3[10][45] , 
        \g3[10][44] , \g3[10][43] , \g3[10][42] , \g3[10][41] , \g3[10][40] , 
        \g3[10][39] , \g3[10][38] , \g3[10][37] , \g3[10][36] , \g3[10][35] , 
        \g3[10][34] , \g3[10][33] , \g3[10][32] , \g3[10][31] , \g3[10][30] , 
        \g3[10][29] , \g3[10][28] , \g3[10][27] , \g3[10][26] , \g3[10][25] , 
        \g3[10][24] , \g3[10][23] , \g3[10][22] , \g3[10][21] , \g3[10][20] , 
        \g3[10][19] , \g3[10][18] , \g3[10][17] , \g3[10][16] , \g3[10][15] , 
        \g3[10][14] , \g3[10][13] , \g3[10][12] , \g3[10][11] , \g3[10][10] , 
        \g3[10][9] , \g3[10][8] , \g3[10][7] , \g3[10][6] , \g3[10][5] , 
        \g3[10][4] , \g3[10][3] , \g3[10][2] , \g3[10][1] , 1'b0}), .cin({
        \g3[11][63] , \g3[11][62] , \g3[11][61] , \g3[11][60] , \g3[11][59] , 
        \g3[11][58] , \g3[11][57] , \g3[11][56] , \g3[11][55] , \g3[11][54] , 
        \g3[11][53] , \g3[11][52] , \g3[11][51] , \g3[11][50] , \g3[11][49] , 
        \g3[11][48] , \g3[11][47] , \g3[11][46] , \g3[11][45] , \g3[11][44] , 
        \g3[11][43] , \g3[11][42] , \g3[11][41] , \g3[11][40] , \g3[11][39] , 
        \g3[11][38] , \g3[11][37] , \g3[11][36] , \g3[11][35] , \g3[11][34] , 
        \g3[11][33] , \g3[11][32] , \g3[11][31] , \g3[11][30] , \g3[11][29] , 
        \g3[11][28] , \g3[11][27] , \g3[11][26] , \g3[11][25] , \g3[11][24] , 
        \g3[11][23] , \g3[11][22] , \g3[11][21] , \g3[11][20] , \g3[11][19] , 
        \g3[11][18] , \g3[11][17] , \g3[11][16] , \g3[11][15] , \g3[11][14] , 
        \g3[11][13] , \g3[11][12] , \g3[11][11] , \g3[11][10] , \g3[11][9] , 
        \g3[11][8] , \g3[11][7] , \g3[11][6] , \g3[11][5] , \g3[11][4] , 
        \g3[11][3] , \g3[11][2] , \g3[11][1] , 1'b0}), .sum({\g4[3][63] , 
        \g4[3][62] , \g4[3][61] , \g4[3][60] , \g4[3][59] , \g4[3][58] , 
        \g4[3][57] , \g4[3][56] , \g4[3][55] , \g4[3][54] , \g4[3][53] , 
        \g4[3][52] , \g4[3][51] , \g4[3][50] , \g4[3][49] , \g4[3][48] , 
        \g4[3][47] , \g4[3][46] , \g4[3][45] , \g4[3][44] , \g4[3][43] , 
        \g4[3][42] , \g4[3][41] , \g4[3][40] , \g4[3][39] , \g4[3][38] , 
        \g4[3][37] , \g4[3][36] , \g4[3][35] , \g4[3][34] , \g4[3][33] , 
        \g4[3][32] , \g4[3][31] , \g4[3][30] , \g4[3][29] , \g4[3][28] , 
        \g4[3][27] , \g4[3][26] , \g4[3][25] , \g4[3][24] , \g4[3][23] , 
        \g4[3][22] , \g4[3][21] , \g4[3][20] , \g4[3][19] , \g4[3][18] , 
        \g4[3][17] , \g4[3][16] , \g4[3][15] , \g4[3][14] , \g4[3][13] , 
        \g4[3][12] , \g4[3][11] , \g4[3][10] , \g4[3][9] , \g4[3][8] , 
        \g4[3][7] , \g4[3][6] , \g4[3][5] , \g4[3][4] , \g4[3][3] , \g4[3][2] , 
        \g4[3][1] , \g4[3][0] }), .cout({\g4[9][63] , \g4[9][62] , \g4[9][61] , 
        \g4[9][60] , \g4[9][59] , \g4[9][58] , \g4[9][57] , \g4[9][56] , 
        \g4[9][55] , \g4[9][54] , \g4[9][53] , \g4[9][52] , \g4[9][51] , 
        \g4[9][50] , \g4[9][49] , \g4[9][48] , \g4[9][47] , \g4[9][46] , 
        \g4[9][45] , \g4[9][44] , \g4[9][43] , \g4[9][42] , \g4[9][41] , 
        \g4[9][40] , \g4[9][39] , \g4[9][38] , \g4[9][37] , \g4[9][36] , 
        \g4[9][35] , \g4[9][34] , \g4[9][33] , \g4[9][32] , \g4[9][31] , 
        \g4[9][30] , \g4[9][29] , \g4[9][28] , \g4[9][27] , \g4[9][26] , 
        \g4[9][25] , \g4[9][24] , \g4[9][23] , \g4[9][22] , \g4[9][21] , 
        \g4[9][20] , \g4[9][19] , \g4[9][18] , \g4[9][17] , \g4[9][16] , 
        \g4[9][15] , \g4[9][14] , \g4[9][13] , \g4[9][12] , \g4[9][11] , 
        \g4[9][10] , \g4[9][9] , \g4[9][8] , \g4[9][7] , \g4[9][6] , 
        \g4[9][5] , \g4[9][4] , \g4[9][3] , \g4[9][2] , \g4[9][1] , 
        SYNOPSYS_UNCONNECTED__47}) );
  FullAdder \level4[4].x1  ( .a({\g3[12][63] , \g3[12][62] , \g3[12][61] , 
        \g3[12][60] , \g3[12][59] , \g3[12][58] , \g3[12][57] , \g3[12][56] , 
        \g3[12][55] , \g3[12][54] , \g3[12][53] , \g3[12][52] , \g3[12][51] , 
        \g3[12][50] , \g3[12][49] , \g3[12][48] , \g3[12][47] , \g3[12][46] , 
        \g3[12][45] , \g3[12][44] , \g3[12][43] , \g3[12][42] , \g3[12][41] , 
        \g3[12][40] , \g3[12][39] , \g3[12][38] , \g3[12][37] , \g3[12][36] , 
        \g3[12][35] , \g3[12][34] , \g3[12][33] , \g3[12][32] , \g3[12][31] , 
        \g3[12][30] , \g3[12][29] , \g3[12][28] , \g3[12][27] , \g3[12][26] , 
        \g3[12][25] , \g3[12][24] , \g3[12][23] , \g3[12][22] , \g3[12][21] , 
        \g3[12][20] , \g3[12][19] , \g3[12][18] , \g3[12][17] , \g3[12][16] , 
        \g3[12][15] , \g3[12][14] , \g3[12][13] , \g3[12][12] , \g3[12][11] , 
        \g3[12][10] , \g3[12][9] , \g3[12][8] , \g3[12][7] , \g3[12][6] , 
        \g3[12][5] , \g3[12][4] , \g3[12][3] , \g3[12][2] , \g3[12][1] , 1'b0}), .b({\g3[13][63] , \g3[13][62] , \g3[13][61] , \g3[13][60] , \g3[13][59] , 
        \g3[13][58] , \g3[13][57] , \g3[13][56] , \g3[13][55] , \g3[13][54] , 
        \g3[13][53] , \g3[13][52] , \g3[13][51] , \g3[13][50] , \g3[13][49] , 
        \g3[13][48] , \g3[13][47] , \g3[13][46] , \g3[13][45] , \g3[13][44] , 
        \g3[13][43] , \g3[13][42] , \g3[13][41] , \g3[13][40] , \g3[13][39] , 
        \g3[13][38] , \g3[13][37] , \g3[13][36] , \g3[13][35] , \g3[13][34] , 
        \g3[13][33] , \g3[13][32] , \g3[13][31] , \g3[13][30] , \g3[13][29] , 
        \g3[13][28] , \g3[13][27] , \g3[13][26] , \g3[13][25] , \g3[13][24] , 
        \g3[13][23] , \g3[13][22] , \g3[13][21] , \g3[13][20] , \g3[13][19] , 
        \g3[13][18] , \g3[13][17] , \g3[13][16] , \g3[13][15] , \g3[13][14] , 
        \g3[13][13] , \g3[13][12] , \g3[13][11] , \g3[13][10] , \g3[13][9] , 
        \g3[13][8] , \g3[13][7] , \g3[13][6] , \g3[13][5] , \g3[13][4] , 
        \g3[13][3] , \g3[13][2] , \g3[13][1] , 1'b0}), .cin({\g3[14][63] , 
        \g3[14][62] , \g3[14][61] , \g3[14][60] , \g3[14][59] , \g3[14][58] , 
        \g3[14][57] , \g3[14][56] , \g3[14][55] , \g3[14][54] , \g3[14][53] , 
        \g3[14][52] , \g3[14][51] , \g3[14][50] , \g3[14][49] , \g3[14][48] , 
        \g3[14][47] , \g3[14][46] , \g3[14][45] , \g3[14][44] , \g3[14][43] , 
        \g3[14][42] , \g3[14][41] , \g3[14][40] , \g3[14][39] , \g3[14][38] , 
        \g3[14][37] , \g3[14][36] , \g3[14][35] , \g3[14][34] , \g3[14][33] , 
        \g3[14][32] , \g3[14][31] , \g3[14][30] , \g3[14][29] , \g3[14][28] , 
        \g3[14][27] , \g3[14][26] , \g3[14][25] , \g3[14][24] , \g3[14][23] , 
        \g3[14][22] , \g3[14][21] , \g3[14][20] , \g3[14][19] , \g3[14][18] , 
        \g3[14][17] , \g3[14][16] , \g3[14][15] , \g3[14][14] , \g3[14][13] , 
        \g3[14][12] , \g3[14][11] , \g3[14][10] , \g3[14][9] , \g3[14][8] , 
        \g3[14][7] , \g3[14][6] , \g3[14][5] , \g3[14][4] , \g3[14][3] , 
        \g3[14][2] , \g3[14][1] , 1'b0}), .sum({\g4[4][63] , \g4[4][62] , 
        \g4[4][61] , \g4[4][60] , \g4[4][59] , \g4[4][58] , \g4[4][57] , 
        \g4[4][56] , \g4[4][55] , \g4[4][54] , \g4[4][53] , \g4[4][52] , 
        \g4[4][51] , \g4[4][50] , \g4[4][49] , \g4[4][48] , \g4[4][47] , 
        \g4[4][46] , \g4[4][45] , \g4[4][44] , \g4[4][43] , \g4[4][42] , 
        \g4[4][41] , \g4[4][40] , \g4[4][39] , \g4[4][38] , \g4[4][37] , 
        \g4[4][36] , \g4[4][35] , \g4[4][34] , \g4[4][33] , \g4[4][32] , 
        \g4[4][31] , \g4[4][30] , \g4[4][29] , \g4[4][28] , \g4[4][27] , 
        \g4[4][26] , \g4[4][25] , \g4[4][24] , \g4[4][23] , \g4[4][22] , 
        \g4[4][21] , \g4[4][20] , \g4[4][19] , \g4[4][18] , \g4[4][17] , 
        \g4[4][16] , \g4[4][15] , \g4[4][14] , \g4[4][13] , \g4[4][12] , 
        \g4[4][11] , \g4[4][10] , \g4[4][9] , \g4[4][8] , \g4[4][7] , 
        \g4[4][6] , \g4[4][5] , \g4[4][4] , \g4[4][3] , \g4[4][2] , \g4[4][1] , 
        \g4[4][0] }), .cout({\g4[10][63] , \g4[10][62] , \g4[10][61] , 
        \g4[10][60] , \g4[10][59] , \g4[10][58] , \g4[10][57] , \g4[10][56] , 
        \g4[10][55] , \g4[10][54] , \g4[10][53] , \g4[10][52] , \g4[10][51] , 
        \g4[10][50] , \g4[10][49] , \g4[10][48] , \g4[10][47] , \g4[10][46] , 
        \g4[10][45] , \g4[10][44] , \g4[10][43] , \g4[10][42] , \g4[10][41] , 
        \g4[10][40] , \g4[10][39] , \g4[10][38] , \g4[10][37] , \g4[10][36] , 
        \g4[10][35] , \g4[10][34] , \g4[10][33] , \g4[10][32] , \g4[10][31] , 
        \g4[10][30] , \g4[10][29] , \g4[10][28] , \g4[10][27] , \g4[10][26] , 
        \g4[10][25] , \g4[10][24] , \g4[10][23] , \g4[10][22] , \g4[10][21] , 
        \g4[10][20] , \g4[10][19] , \g4[10][18] , \g4[10][17] , \g4[10][16] , 
        \g4[10][15] , \g4[10][14] , \g4[10][13] , \g4[10][12] , \g4[10][11] , 
        \g4[10][10] , \g4[10][9] , \g4[10][8] , \g4[10][7] , \g4[10][6] , 
        \g4[10][5] , \g4[10][4] , \g4[10][3] , \g4[10][2] , \g4[10][1] , 
        SYNOPSYS_UNCONNECTED__48}) );
  FullAdder \level4[5].x1  ( .a({\g3[15][63] , \g3[15][62] , \g3[15][61] , 
        \g3[15][60] , \g3[15][59] , \g3[15][58] , \g3[15][57] , \g3[15][56] , 
        \g3[15][55] , \g3[15][54] , \g3[15][53] , \g3[15][52] , \g3[15][51] , 
        \g3[15][50] , \g3[15][49] , \g3[15][48] , \g3[15][47] , \g3[15][46] , 
        \g3[15][45] , \g3[15][44] , \g3[15][43] , \g3[15][42] , \g3[15][41] , 
        \g3[15][40] , \g3[15][39] , \g3[15][38] , \g3[15][37] , \g3[15][36] , 
        \g3[15][35] , \g3[15][34] , \g3[15][33] , \g3[15][32] , \g3[15][31] , 
        \g3[15][30] , \g3[15][29] , \g3[15][28] , \g3[15][27] , \g3[15][26] , 
        \g3[15][25] , \g3[15][24] , \g3[15][23] , \g3[15][22] , \g3[15][21] , 
        \g3[15][20] , \g3[15][19] , \g3[15][18] , \g3[15][17] , \g3[15][16] , 
        \g3[15][15] , \g3[15][14] , \g3[15][13] , \g3[15][12] , \g3[15][11] , 
        \g3[15][10] , \g3[15][9] , \g3[15][8] , \g3[15][7] , \g3[15][6] , 
        \g3[15][5] , \g3[15][4] , \g3[15][3] , \g3[15][2] , \g3[15][1] , 1'b0}), .b({\g3[16][63] , \g3[16][62] , \g3[16][61] , \g3[16][60] , \g3[16][59] , 
        \g3[16][58] , \g3[16][57] , \g3[16][56] , \g3[16][55] , \g3[16][54] , 
        \g3[16][53] , \g3[16][52] , \g3[16][51] , \g3[16][50] , \g3[16][49] , 
        \g3[16][48] , \g3[16][47] , \g3[16][46] , \g3[16][45] , \g3[16][44] , 
        \g3[16][43] , \g3[16][42] , \g3[16][41] , \g3[16][40] , \g3[16][39] , 
        \g3[16][38] , \g3[16][37] , \g3[16][36] , \g3[16][35] , \g3[16][34] , 
        \g3[16][33] , \g3[16][32] , \g3[16][31] , \g3[16][30] , \g3[16][29] , 
        \g3[16][28] , \g3[16][27] , \g3[16][26] , \g3[16][25] , \g3[16][24] , 
        \g3[16][23] , \g3[16][22] , \g3[16][21] , \g3[16][20] , \g3[16][19] , 
        \g3[16][18] , \g3[16][17] , \g3[16][16] , \g3[16][15] , \g3[16][14] , 
        \g3[16][13] , \g3[16][12] , \g3[16][11] , \g3[16][10] , \g3[16][9] , 
        \g3[16][8] , \g3[16][7] , \g3[16][6] , \g3[16][5] , \g3[16][4] , 
        \g3[16][3] , \g3[16][2] , \g3[16][1] , 1'b0}), .cin({\g3[17][63] , 
        \g3[17][62] , \g3[17][61] , \g3[17][60] , \g3[17][59] , \g3[17][58] , 
        \g3[17][57] , \g3[17][56] , \g3[17][55] , \g3[17][54] , \g3[17][53] , 
        \g3[17][52] , \g3[17][51] , \g3[17][50] , \g3[17][49] , \g3[17][48] , 
        \g3[17][47] , \g3[17][46] , \g3[17][45] , \g3[17][44] , \g3[17][43] , 
        \g3[17][42] , \g3[17][41] , \g3[17][40] , \g3[17][39] , \g3[17][38] , 
        \g3[17][37] , \g3[17][36] , \g3[17][35] , \g3[17][34] , \g3[17][33] , 
        \g3[17][32] , \g3[17][31] , \g3[17][30] , \g3[17][29] , \g3[17][28] , 
        \g3[17][27] , \g3[17][26] , \g3[17][25] , \g3[17][24] , \g3[17][23] , 
        \g3[17][22] , \g3[17][21] , \g3[17][20] , \g3[17][19] , \g3[17][18] , 
        \g3[17][17] , \g3[17][16] , \g3[17][15] , \g3[17][14] , \g3[17][13] , 
        \g3[17][12] , \g3[17][11] , \g3[17][10] , \g3[17][9] , \g3[17][8] , 
        \g3[17][7] , \g3[17][6] , \g3[17][5] , \g3[17][4] , \g3[17][3] , 
        \g3[17][2] , \g3[17][1] , 1'b0}), .sum({\g4[5][63] , \g4[5][62] , 
        \g4[5][61] , \g4[5][60] , \g4[5][59] , \g4[5][58] , \g4[5][57] , 
        \g4[5][56] , \g4[5][55] , \g4[5][54] , \g4[5][53] , \g4[5][52] , 
        \g4[5][51] , \g4[5][50] , \g4[5][49] , \g4[5][48] , \g4[5][47] , 
        \g4[5][46] , \g4[5][45] , \g4[5][44] , \g4[5][43] , \g4[5][42] , 
        \g4[5][41] , \g4[5][40] , \g4[5][39] , \g4[5][38] , \g4[5][37] , 
        \g4[5][36] , \g4[5][35] , \g4[5][34] , \g4[5][33] , \g4[5][32] , 
        \g4[5][31] , \g4[5][30] , \g4[5][29] , \g4[5][28] , \g4[5][27] , 
        \g4[5][26] , \g4[5][25] , \g4[5][24] , \g4[5][23] , \g4[5][22] , 
        \g4[5][21] , \g4[5][20] , \g4[5][19] , \g4[5][18] , \g4[5][17] , 
        \g4[5][16] , \g4[5][15] , \g4[5][14] , \g4[5][13] , \g4[5][12] , 
        \g4[5][11] , \g4[5][10] , \g4[5][9] , \g4[5][8] , \g4[5][7] , 
        \g4[5][6] , \g4[5][5] , \g4[5][4] , \g4[5][3] , \g4[5][2] , \g4[5][1] , 
        \g4[5][0] }), .cout({\g4[11][63] , \g4[11][62] , \g4[11][61] , 
        \g4[11][60] , \g4[11][59] , \g4[11][58] , \g4[11][57] , \g4[11][56] , 
        \g4[11][55] , \g4[11][54] , \g4[11][53] , \g4[11][52] , \g4[11][51] , 
        \g4[11][50] , \g4[11][49] , \g4[11][48] , \g4[11][47] , \g4[11][46] , 
        \g4[11][45] , \g4[11][44] , \g4[11][43] , \g4[11][42] , \g4[11][41] , 
        \g4[11][40] , \g4[11][39] , \g4[11][38] , \g4[11][37] , \g4[11][36] , 
        \g4[11][35] , \g4[11][34] , \g4[11][33] , \g4[11][32] , \g4[11][31] , 
        \g4[11][30] , \g4[11][29] , \g4[11][28] , \g4[11][27] , \g4[11][26] , 
        \g4[11][25] , \g4[11][24] , \g4[11][23] , \g4[11][22] , \g4[11][21] , 
        \g4[11][20] , \g4[11][19] , \g4[11][18] , \g4[11][17] , \g4[11][16] , 
        \g4[11][15] , \g4[11][14] , \g4[11][13] , \g4[11][12] , \g4[11][11] , 
        \g4[11][10] , \g4[11][9] , \g4[11][8] , \g4[11][7] , \g4[11][6] , 
        \g4[11][5] , \g4[11][4] , \g4[11][3] , \g4[11][2] , \g4[11][1] , 
        SYNOPSYS_UNCONNECTED__49}) );
  FullAdder \level5[0].x2  ( .a({\g4[0][63] , \g4[0][62] , \g4[0][61] , 
        \g4[0][60] , \g4[0][59] , \g4[0][58] , \g4[0][57] , \g4[0][56] , 
        \g4[0][55] , \g4[0][54] , \g4[0][53] , \g4[0][52] , \g4[0][51] , 
        \g4[0][50] , \g4[0][49] , \g4[0][48] , \g4[0][47] , \g4[0][46] , 
        \g4[0][45] , \g4[0][44] , \g4[0][43] , \g4[0][42] , \g4[0][41] , 
        \g4[0][40] , \g4[0][39] , \g4[0][38] , \g4[0][37] , \g4[0][36] , 
        \g4[0][35] , \g4[0][34] , \g4[0][33] , \g4[0][32] , \g4[0][31] , 
        \g4[0][30] , \g4[0][29] , \g4[0][28] , \g4[0][27] , \g4[0][26] , 
        \g4[0][25] , \g4[0][24] , \g4[0][23] , \g4[0][22] , \g4[0][21] , 
        \g4[0][20] , \g4[0][19] , \g4[0][18] , \g4[0][17] , \g4[0][16] , 
        \g4[0][15] , \g4[0][14] , \g4[0][13] , \g4[0][12] , \g4[0][11] , 
        \g4[0][10] , \g4[0][9] , \g4[0][8] , \g4[0][7] , \g4[0][6] , 
        \g4[0][5] , \g4[0][4] , \g4[0][3] , \g4[0][2] , \g4[0][1] , \g4[0][0] }), .b({\g4[1][63] , \g4[1][62] , \g4[1][61] , \g4[1][60] , \g4[1][59] , 
        \g4[1][58] , \g4[1][57] , \g4[1][56] , \g4[1][55] , \g4[1][54] , 
        \g4[1][53] , \g4[1][52] , \g4[1][51] , \g4[1][50] , \g4[1][49] , 
        \g4[1][48] , \g4[1][47] , \g4[1][46] , \g4[1][45] , \g4[1][44] , 
        \g4[1][43] , \g4[1][42] , \g4[1][41] , \g4[1][40] , \g4[1][39] , 
        \g4[1][38] , \g4[1][37] , \g4[1][36] , \g4[1][35] , \g4[1][34] , 
        \g4[1][33] , \g4[1][32] , \g4[1][31] , \g4[1][30] , \g4[1][29] , 
        \g4[1][28] , \g4[1][27] , \g4[1][26] , \g4[1][25] , \g4[1][24] , 
        \g4[1][23] , \g4[1][22] , \g4[1][21] , \g4[1][20] , \g4[1][19] , 
        \g4[1][18] , \g4[1][17] , \g4[1][16] , \g4[1][15] , \g4[1][14] , 
        \g4[1][13] , \g4[1][12] , \g4[1][11] , \g4[1][10] , \g4[1][9] , 
        \g4[1][8] , \g4[1][7] , \g4[1][6] , \g4[1][5] , \g4[1][4] , \g4[1][3] , 
        \g4[1][2] , \g4[1][1] , \g4[1][0] }), .cin({\g4[2][63] , \g4[2][62] , 
        \g4[2][61] , \g4[2][60] , \g4[2][59] , \g4[2][58] , \g4[2][57] , 
        \g4[2][56] , \g4[2][55] , \g4[2][54] , \g4[2][53] , \g4[2][52] , 
        \g4[2][51] , \g4[2][50] , \g4[2][49] , \g4[2][48] , \g4[2][47] , 
        \g4[2][46] , \g4[2][45] , \g4[2][44] , \g4[2][43] , \g4[2][42] , 
        \g4[2][41] , \g4[2][40] , \g4[2][39] , \g4[2][38] , \g4[2][37] , 
        \g4[2][36] , \g4[2][35] , \g4[2][34] , \g4[2][33] , \g4[2][32] , 
        \g4[2][31] , \g4[2][30] , \g4[2][29] , \g4[2][28] , \g4[2][27] , 
        \g4[2][26] , \g4[2][25] , \g4[2][24] , \g4[2][23] , \g4[2][22] , 
        \g4[2][21] , \g4[2][20] , \g4[2][19] , \g4[2][18] , \g4[2][17] , 
        \g4[2][16] , \g4[2][15] , \g4[2][14] , \g4[2][13] , \g4[2][12] , 
        \g4[2][11] , \g4[2][10] , \g4[2][9] , \g4[2][8] , \g4[2][7] , 
        \g4[2][6] , \g4[2][5] , \g4[2][4] , \g4[2][3] , \g4[2][2] , \g4[2][1] , 
        \g4[2][0] }), .sum({\g5[0][63] , \g5[0][62] , \g5[0][61] , \g5[0][60] , 
        \g5[0][59] , \g5[0][58] , \g5[0][57] , \g5[0][56] , \g5[0][55] , 
        \g5[0][54] , \g5[0][53] , \g5[0][52] , \g5[0][51] , \g5[0][50] , 
        \g5[0][49] , \g5[0][48] , \g5[0][47] , \g5[0][46] , \g5[0][45] , 
        \g5[0][44] , \g5[0][43] , \g5[0][42] , \g5[0][41] , \g5[0][40] , 
        \g5[0][39] , \g5[0][38] , \g5[0][37] , \g5[0][36] , \g5[0][35] , 
        \g5[0][34] , \g5[0][33] , \g5[0][32] , \g5[0][31] , \g5[0][30] , 
        \g5[0][29] , \g5[0][28] , \g5[0][27] , \g5[0][26] , \g5[0][25] , 
        \g5[0][24] , \g5[0][23] , \g5[0][22] , \g5[0][21] , \g5[0][20] , 
        \g5[0][19] , \g5[0][18] , \g5[0][17] , \g5[0][16] , \g5[0][15] , 
        \g5[0][14] , \g5[0][13] , \g5[0][12] , \g5[0][11] , \g5[0][10] , 
        \g5[0][9] , \g5[0][8] , \g5[0][7] , \g5[0][6] , \g5[0][5] , \g5[0][4] , 
        \g5[0][3] , \g5[0][2] , \g5[0][1] , \g5[0][0] }), .cout({\g5[4][63] , 
        \g5[4][62] , \g5[4][61] , \g5[4][60] , \g5[4][59] , \g5[4][58] , 
        \g5[4][57] , \g5[4][56] , \g5[4][55] , \g5[4][54] , \g5[4][53] , 
        \g5[4][52] , \g5[4][51] , \g5[4][50] , \g5[4][49] , \g5[4][48] , 
        \g5[4][47] , \g5[4][46] , \g5[4][45] , \g5[4][44] , \g5[4][43] , 
        \g5[4][42] , \g5[4][41] , \g5[4][40] , \g5[4][39] , \g5[4][38] , 
        \g5[4][37] , \g5[4][36] , \g5[4][35] , \g5[4][34] , \g5[4][33] , 
        \g5[4][32] , \g5[4][31] , \g5[4][30] , \g5[4][29] , \g5[4][28] , 
        \g5[4][27] , \g5[4][26] , \g5[4][25] , \g5[4][24] , \g5[4][23] , 
        \g5[4][22] , \g5[4][21] , \g5[4][20] , \g5[4][19] , \g5[4][18] , 
        \g5[4][17] , \g5[4][16] , \g5[4][15] , \g5[4][14] , \g5[4][13] , 
        \g5[4][12] , \g5[4][11] , \g5[4][10] , \g5[4][9] , \g5[4][8] , 
        \g5[4][7] , \g5[4][6] , \g5[4][5] , \g5[4][4] , \g5[4][3] , \g5[4][2] , 
        \g5[4][1] , SYNOPSYS_UNCONNECTED__50}) );
  FullAdder \level5[1].x2  ( .a({\g4[3][63] , \g4[3][62] , \g4[3][61] , 
        \g4[3][60] , \g4[3][59] , \g4[3][58] , \g4[3][57] , \g4[3][56] , 
        \g4[3][55] , \g4[3][54] , \g4[3][53] , \g4[3][52] , \g4[3][51] , 
        \g4[3][50] , \g4[3][49] , \g4[3][48] , \g4[3][47] , \g4[3][46] , 
        \g4[3][45] , \g4[3][44] , \g4[3][43] , \g4[3][42] , \g4[3][41] , 
        \g4[3][40] , \g4[3][39] , \g4[3][38] , \g4[3][37] , \g4[3][36] , 
        \g4[3][35] , \g4[3][34] , \g4[3][33] , \g4[3][32] , \g4[3][31] , 
        \g4[3][30] , \g4[3][29] , \g4[3][28] , \g4[3][27] , \g4[3][26] , 
        \g4[3][25] , \g4[3][24] , \g4[3][23] , \g4[3][22] , \g4[3][21] , 
        \g4[3][20] , \g4[3][19] , \g4[3][18] , \g4[3][17] , \g4[3][16] , 
        \g4[3][15] , \g4[3][14] , \g4[3][13] , \g4[3][12] , \g4[3][11] , 
        \g4[3][10] , \g4[3][9] , \g4[3][8] , \g4[3][7] , \g4[3][6] , 
        \g4[3][5] , \g4[3][4] , \g4[3][3] , \g4[3][2] , \g4[3][1] , \g4[3][0] }), .b({\g4[4][63] , \g4[4][62] , \g4[4][61] , \g4[4][60] , \g4[4][59] , 
        \g4[4][58] , \g4[4][57] , \g4[4][56] , \g4[4][55] , \g4[4][54] , 
        \g4[4][53] , \g4[4][52] , \g4[4][51] , \g4[4][50] , \g4[4][49] , 
        \g4[4][48] , \g4[4][47] , \g4[4][46] , \g4[4][45] , \g4[4][44] , 
        \g4[4][43] , \g4[4][42] , \g4[4][41] , \g4[4][40] , \g4[4][39] , 
        \g4[4][38] , \g4[4][37] , \g4[4][36] , \g4[4][35] , \g4[4][34] , 
        \g4[4][33] , \g4[4][32] , \g4[4][31] , \g4[4][30] , \g4[4][29] , 
        \g4[4][28] , \g4[4][27] , \g4[4][26] , \g4[4][25] , \g4[4][24] , 
        \g4[4][23] , \g4[4][22] , \g4[4][21] , \g4[4][20] , \g4[4][19] , 
        \g4[4][18] , \g4[4][17] , \g4[4][16] , \g4[4][15] , \g4[4][14] , 
        \g4[4][13] , \g4[4][12] , \g4[4][11] , \g4[4][10] , \g4[4][9] , 
        \g4[4][8] , \g4[4][7] , \g4[4][6] , \g4[4][5] , \g4[4][4] , \g4[4][3] , 
        \g4[4][2] , \g4[4][1] , \g4[4][0] }), .cin({\g4[5][63] , \g4[5][62] , 
        \g4[5][61] , \g4[5][60] , \g4[5][59] , \g4[5][58] , \g4[5][57] , 
        \g4[5][56] , \g4[5][55] , \g4[5][54] , \g4[5][53] , \g4[5][52] , 
        \g4[5][51] , \g4[5][50] , \g4[5][49] , \g4[5][48] , \g4[5][47] , 
        \g4[5][46] , \g4[5][45] , \g4[5][44] , \g4[5][43] , \g4[5][42] , 
        \g4[5][41] , \g4[5][40] , \g4[5][39] , \g4[5][38] , \g4[5][37] , 
        \g4[5][36] , \g4[5][35] , \g4[5][34] , \g4[5][33] , \g4[5][32] , 
        \g4[5][31] , \g4[5][30] , \g4[5][29] , \g4[5][28] , \g4[5][27] , 
        \g4[5][26] , \g4[5][25] , \g4[5][24] , \g4[5][23] , \g4[5][22] , 
        \g4[5][21] , \g4[5][20] , \g4[5][19] , \g4[5][18] , \g4[5][17] , 
        \g4[5][16] , \g4[5][15] , \g4[5][14] , \g4[5][13] , \g4[5][12] , 
        \g4[5][11] , \g4[5][10] , \g4[5][9] , \g4[5][8] , \g4[5][7] , 
        \g4[5][6] , \g4[5][5] , \g4[5][4] , \g4[5][3] , \g4[5][2] , \g4[5][1] , 
        \g4[5][0] }), .sum({\g5[1][63] , \g5[1][62] , \g5[1][61] , \g5[1][60] , 
        \g5[1][59] , \g5[1][58] , \g5[1][57] , \g5[1][56] , \g5[1][55] , 
        \g5[1][54] , \g5[1][53] , \g5[1][52] , \g5[1][51] , \g5[1][50] , 
        \g5[1][49] , \g5[1][48] , \g5[1][47] , \g5[1][46] , \g5[1][45] , 
        \g5[1][44] , \g5[1][43] , \g5[1][42] , \g5[1][41] , \g5[1][40] , 
        \g5[1][39] , \g5[1][38] , \g5[1][37] , \g5[1][36] , \g5[1][35] , 
        \g5[1][34] , \g5[1][33] , \g5[1][32] , \g5[1][31] , \g5[1][30] , 
        \g5[1][29] , \g5[1][28] , \g5[1][27] , \g5[1][26] , \g5[1][25] , 
        \g5[1][24] , \g5[1][23] , \g5[1][22] , \g5[1][21] , \g5[1][20] , 
        \g5[1][19] , \g5[1][18] , \g5[1][17] , \g5[1][16] , \g5[1][15] , 
        \g5[1][14] , \g5[1][13] , \g5[1][12] , \g5[1][11] , \g5[1][10] , 
        \g5[1][9] , \g5[1][8] , \g5[1][7] , \g5[1][6] , \g5[1][5] , \g5[1][4] , 
        \g5[1][3] , \g5[1][2] , \g5[1][1] , \g5[1][0] }), .cout({\g5[5][63] , 
        \g5[5][62] , \g5[5][61] , \g5[5][60] , \g5[5][59] , \g5[5][58] , 
        \g5[5][57] , \g5[5][56] , \g5[5][55] , \g5[5][54] , \g5[5][53] , 
        \g5[5][52] , \g5[5][51] , \g5[5][50] , \g5[5][49] , \g5[5][48] , 
        \g5[5][47] , \g5[5][46] , \g5[5][45] , \g5[5][44] , \g5[5][43] , 
        \g5[5][42] , \g5[5][41] , \g5[5][40] , \g5[5][39] , \g5[5][38] , 
        \g5[5][37] , \g5[5][36] , \g5[5][35] , \g5[5][34] , \g5[5][33] , 
        \g5[5][32] , \g5[5][31] , \g5[5][30] , \g5[5][29] , \g5[5][28] , 
        \g5[5][27] , \g5[5][26] , \g5[5][25] , \g5[5][24] , \g5[5][23] , 
        \g5[5][22] , \g5[5][21] , \g5[5][20] , \g5[5][19] , \g5[5][18] , 
        \g5[5][17] , \g5[5][16] , \g5[5][15] , \g5[5][14] , \g5[5][13] , 
        \g5[5][12] , \g5[5][11] , \g5[5][10] , \g5[5][9] , \g5[5][8] , 
        \g5[5][7] , \g5[5][6] , \g5[5][5] , \g5[5][4] , \g5[5][3] , \g5[5][2] , 
        \g5[5][1] , SYNOPSYS_UNCONNECTED__51}) );
  FullAdder \level5[2].x2  ( .a({\g4[6][63] , \g4[6][62] , \g4[6][61] , 
        \g4[6][60] , \g4[6][59] , \g4[6][58] , \g4[6][57] , \g4[6][56] , 
        \g4[6][55] , \g4[6][54] , \g4[6][53] , \g4[6][52] , \g4[6][51] , 
        \g4[6][50] , \g4[6][49] , \g4[6][48] , \g4[6][47] , \g4[6][46] , 
        \g4[6][45] , \g4[6][44] , \g4[6][43] , \g4[6][42] , \g4[6][41] , 
        \g4[6][40] , \g4[6][39] , \g4[6][38] , \g4[6][37] , \g4[6][36] , 
        \g4[6][35] , \g4[6][34] , \g4[6][33] , \g4[6][32] , \g4[6][31] , 
        \g4[6][30] , \g4[6][29] , \g4[6][28] , \g4[6][27] , \g4[6][26] , 
        \g4[6][25] , \g4[6][24] , \g4[6][23] , \g4[6][22] , \g4[6][21] , 
        \g4[6][20] , \g4[6][19] , \g4[6][18] , \g4[6][17] , \g4[6][16] , 
        \g4[6][15] , \g4[6][14] , \g4[6][13] , \g4[6][12] , \g4[6][11] , 
        \g4[6][10] , \g4[6][9] , \g4[6][8] , \g4[6][7] , \g4[6][6] , 
        \g4[6][5] , \g4[6][4] , \g4[6][3] , \g4[6][2] , \g4[6][1] , 1'b0}), 
        .b({\g4[7][63] , \g4[7][62] , \g4[7][61] , \g4[7][60] , \g4[7][59] , 
        \g4[7][58] , \g4[7][57] , \g4[7][56] , \g4[7][55] , \g4[7][54] , 
        \g4[7][53] , \g4[7][52] , \g4[7][51] , \g4[7][50] , \g4[7][49] , 
        \g4[7][48] , \g4[7][47] , \g4[7][46] , \g4[7][45] , \g4[7][44] , 
        \g4[7][43] , \g4[7][42] , \g4[7][41] , \g4[7][40] , \g4[7][39] , 
        \g4[7][38] , \g4[7][37] , \g4[7][36] , \g4[7][35] , \g4[7][34] , 
        \g4[7][33] , \g4[7][32] , \g4[7][31] , \g4[7][30] , \g4[7][29] , 
        \g4[7][28] , \g4[7][27] , \g4[7][26] , \g4[7][25] , \g4[7][24] , 
        \g4[7][23] , \g4[7][22] , \g4[7][21] , \g4[7][20] , \g4[7][19] , 
        \g4[7][18] , \g4[7][17] , \g4[7][16] , \g4[7][15] , \g4[7][14] , 
        \g4[7][13] , \g4[7][12] , \g4[7][11] , \g4[7][10] , \g4[7][9] , 
        \g4[7][8] , \g4[7][7] , \g4[7][6] , \g4[7][5] , \g4[7][4] , \g4[7][3] , 
        \g4[7][2] , \g4[7][1] , 1'b0}), .cin({\g4[8][63] , \g4[8][62] , 
        \g4[8][61] , \g4[8][60] , \g4[8][59] , \g4[8][58] , \g4[8][57] , 
        \g4[8][56] , \g4[8][55] , \g4[8][54] , \g4[8][53] , \g4[8][52] , 
        \g4[8][51] , \g4[8][50] , \g4[8][49] , \g4[8][48] , \g4[8][47] , 
        \g4[8][46] , \g4[8][45] , \g4[8][44] , \g4[8][43] , \g4[8][42] , 
        \g4[8][41] , \g4[8][40] , \g4[8][39] , \g4[8][38] , \g4[8][37] , 
        \g4[8][36] , \g4[8][35] , \g4[8][34] , \g4[8][33] , \g4[8][32] , 
        \g4[8][31] , \g4[8][30] , \g4[8][29] , \g4[8][28] , \g4[8][27] , 
        \g4[8][26] , \g4[8][25] , \g4[8][24] , \g4[8][23] , \g4[8][22] , 
        \g4[8][21] , \g4[8][20] , \g4[8][19] , \g4[8][18] , \g4[8][17] , 
        \g4[8][16] , \g4[8][15] , \g4[8][14] , \g4[8][13] , \g4[8][12] , 
        \g4[8][11] , \g4[8][10] , \g4[8][9] , \g4[8][8] , \g4[8][7] , 
        \g4[8][6] , \g4[8][5] , \g4[8][4] , \g4[8][3] , \g4[8][2] , \g4[8][1] , 
        1'b0}), .sum({\g5[2][63] , \g5[2][62] , \g5[2][61] , \g5[2][60] , 
        \g5[2][59] , \g5[2][58] , \g5[2][57] , \g5[2][56] , \g5[2][55] , 
        \g5[2][54] , \g5[2][53] , \g5[2][52] , \g5[2][51] , \g5[2][50] , 
        \g5[2][49] , \g5[2][48] , \g5[2][47] , \g5[2][46] , \g5[2][45] , 
        \g5[2][44] , \g5[2][43] , \g5[2][42] , \g5[2][41] , \g5[2][40] , 
        \g5[2][39] , \g5[2][38] , \g5[2][37] , \g5[2][36] , \g5[2][35] , 
        \g5[2][34] , \g5[2][33] , \g5[2][32] , \g5[2][31] , \g5[2][30] , 
        \g5[2][29] , \g5[2][28] , \g5[2][27] , \g5[2][26] , \g5[2][25] , 
        \g5[2][24] , \g5[2][23] , \g5[2][22] , \g5[2][21] , \g5[2][20] , 
        \g5[2][19] , \g5[2][18] , \g5[2][17] , \g5[2][16] , \g5[2][15] , 
        \g5[2][14] , \g5[2][13] , \g5[2][12] , \g5[2][11] , \g5[2][10] , 
        \g5[2][9] , \g5[2][8] , \g5[2][7] , \g5[2][6] , \g5[2][5] , \g5[2][4] , 
        \g5[2][3] , \g5[2][2] , \g5[2][1] , \g5[2][0] }), .cout({\g5[6][63] , 
        \g5[6][62] , \g5[6][61] , \g5[6][60] , \g5[6][59] , \g5[6][58] , 
        \g5[6][57] , \g5[6][56] , \g5[6][55] , \g5[6][54] , \g5[6][53] , 
        \g5[6][52] , \g5[6][51] , \g5[6][50] , \g5[6][49] , \g5[6][48] , 
        \g5[6][47] , \g5[6][46] , \g5[6][45] , \g5[6][44] , \g5[6][43] , 
        \g5[6][42] , \g5[6][41] , \g5[6][40] , \g5[6][39] , \g5[6][38] , 
        \g5[6][37] , \g5[6][36] , \g5[6][35] , \g5[6][34] , \g5[6][33] , 
        \g5[6][32] , \g5[6][31] , \g5[6][30] , \g5[6][29] , \g5[6][28] , 
        \g5[6][27] , \g5[6][26] , \g5[6][25] , \g5[6][24] , \g5[6][23] , 
        \g5[6][22] , \g5[6][21] , \g5[6][20] , \g5[6][19] , \g5[6][18] , 
        \g5[6][17] , \g5[6][16] , \g5[6][15] , \g5[6][14] , \g5[6][13] , 
        \g5[6][12] , \g5[6][11] , \g5[6][10] , \g5[6][9] , \g5[6][8] , 
        \g5[6][7] , \g5[6][6] , \g5[6][5] , \g5[6][4] , \g5[6][3] , \g5[6][2] , 
        \g5[6][1] , SYNOPSYS_UNCONNECTED__52}) );
  FullAdder \level5[3].x2  ( .a({\g4[9][63] , \g4[9][62] , \g4[9][61] , 
        \g4[9][60] , \g4[9][59] , \g4[9][58] , \g4[9][57] , \g4[9][56] , 
        \g4[9][55] , \g4[9][54] , \g4[9][53] , \g4[9][52] , \g4[9][51] , 
        \g4[9][50] , \g4[9][49] , \g4[9][48] , \g4[9][47] , \g4[9][46] , 
        \g4[9][45] , \g4[9][44] , \g4[9][43] , \g4[9][42] , \g4[9][41] , 
        \g4[9][40] , \g4[9][39] , \g4[9][38] , \g4[9][37] , \g4[9][36] , 
        \g4[9][35] , \g4[9][34] , \g4[9][33] , \g4[9][32] , \g4[9][31] , 
        \g4[9][30] , \g4[9][29] , \g4[9][28] , \g4[9][27] , \g4[9][26] , 
        \g4[9][25] , \g4[9][24] , \g4[9][23] , \g4[9][22] , \g4[9][21] , 
        \g4[9][20] , \g4[9][19] , \g4[9][18] , \g4[9][17] , \g4[9][16] , 
        \g4[9][15] , \g4[9][14] , \g4[9][13] , \g4[9][12] , \g4[9][11] , 
        \g4[9][10] , \g4[9][9] , \g4[9][8] , \g4[9][7] , \g4[9][6] , 
        \g4[9][5] , \g4[9][4] , \g4[9][3] , \g4[9][2] , \g4[9][1] , 1'b0}), 
        .b({\g4[10][63] , \g4[10][62] , \g4[10][61] , \g4[10][60] , 
        \g4[10][59] , \g4[10][58] , \g4[10][57] , \g4[10][56] , \g4[10][55] , 
        \g4[10][54] , \g4[10][53] , \g4[10][52] , \g4[10][51] , \g4[10][50] , 
        \g4[10][49] , \g4[10][48] , \g4[10][47] , \g4[10][46] , \g4[10][45] , 
        \g4[10][44] , \g4[10][43] , \g4[10][42] , \g4[10][41] , \g4[10][40] , 
        \g4[10][39] , \g4[10][38] , \g4[10][37] , \g4[10][36] , \g4[10][35] , 
        \g4[10][34] , \g4[10][33] , \g4[10][32] , \g4[10][31] , \g4[10][30] , 
        \g4[10][29] , \g4[10][28] , \g4[10][27] , \g4[10][26] , \g4[10][25] , 
        \g4[10][24] , \g4[10][23] , \g4[10][22] , \g4[10][21] , \g4[10][20] , 
        \g4[10][19] , \g4[10][18] , \g4[10][17] , \g4[10][16] , \g4[10][15] , 
        \g4[10][14] , \g4[10][13] , \g4[10][12] , \g4[10][11] , \g4[10][10] , 
        \g4[10][9] , \g4[10][8] , \g4[10][7] , \g4[10][6] , \g4[10][5] , 
        \g4[10][4] , \g4[10][3] , \g4[10][2] , \g4[10][1] , 1'b0}), .cin({
        \g4[11][63] , \g4[11][62] , \g4[11][61] , \g4[11][60] , \g4[11][59] , 
        \g4[11][58] , \g4[11][57] , \g4[11][56] , \g4[11][55] , \g4[11][54] , 
        \g4[11][53] , \g4[11][52] , \g4[11][51] , \g4[11][50] , \g4[11][49] , 
        \g4[11][48] , \g4[11][47] , \g4[11][46] , \g4[11][45] , \g4[11][44] , 
        \g4[11][43] , \g4[11][42] , \g4[11][41] , \g4[11][40] , \g4[11][39] , 
        \g4[11][38] , \g4[11][37] , \g4[11][36] , \g4[11][35] , \g4[11][34] , 
        \g4[11][33] , \g4[11][32] , \g4[11][31] , \g4[11][30] , \g4[11][29] , 
        \g4[11][28] , \g4[11][27] , \g4[11][26] , \g4[11][25] , \g4[11][24] , 
        \g4[11][23] , \g4[11][22] , \g4[11][21] , \g4[11][20] , \g4[11][19] , 
        \g4[11][18] , \g4[11][17] , \g4[11][16] , \g4[11][15] , \g4[11][14] , 
        \g4[11][13] , \g4[11][12] , \g4[11][11] , \g4[11][10] , \g4[11][9] , 
        \g4[11][8] , \g4[11][7] , \g4[11][6] , \g4[11][5] , \g4[11][4] , 
        \g4[11][3] , \g4[11][2] , \g4[11][1] , 1'b0}), .sum({\g5[3][63] , 
        \g5[3][62] , \g5[3][61] , \g5[3][60] , \g5[3][59] , \g5[3][58] , 
        \g5[3][57] , \g5[3][56] , \g5[3][55] , \g5[3][54] , \g5[3][53] , 
        \g5[3][52] , \g5[3][51] , \g5[3][50] , \g5[3][49] , \g5[3][48] , 
        \g5[3][47] , \g5[3][46] , \g5[3][45] , \g5[3][44] , \g5[3][43] , 
        \g5[3][42] , \g5[3][41] , \g5[3][40] , \g5[3][39] , \g5[3][38] , 
        \g5[3][37] , \g5[3][36] , \g5[3][35] , \g5[3][34] , \g5[3][33] , 
        \g5[3][32] , \g5[3][31] , \g5[3][30] , \g5[3][29] , \g5[3][28] , 
        \g5[3][27] , \g5[3][26] , \g5[3][25] , \g5[3][24] , \g5[3][23] , 
        \g5[3][22] , \g5[3][21] , \g5[3][20] , \g5[3][19] , \g5[3][18] , 
        \g5[3][17] , \g5[3][16] , \g5[3][15] , \g5[3][14] , \g5[3][13] , 
        \g5[3][12] , \g5[3][11] , \g5[3][10] , \g5[3][9] , \g5[3][8] , 
        \g5[3][7] , \g5[3][6] , \g5[3][5] , \g5[3][4] , \g5[3][3] , \g5[3][2] , 
        \g5[3][1] , \g5[3][0] }), .cout({\g5[7][63] , \g5[7][62] , \g5[7][61] , 
        \g5[7][60] , \g5[7][59] , \g5[7][58] , \g5[7][57] , \g5[7][56] , 
        \g5[7][55] , \g5[7][54] , \g5[7][53] , \g5[7][52] , \g5[7][51] , 
        \g5[7][50] , \g5[7][49] , \g5[7][48] , \g5[7][47] , \g5[7][46] , 
        \g5[7][45] , \g5[7][44] , \g5[7][43] , \g5[7][42] , \g5[7][41] , 
        \g5[7][40] , \g5[7][39] , \g5[7][38] , \g5[7][37] , \g5[7][36] , 
        \g5[7][35] , \g5[7][34] , \g5[7][33] , \g5[7][32] , \g5[7][31] , 
        \g5[7][30] , \g5[7][29] , \g5[7][28] , \g5[7][27] , \g5[7][26] , 
        \g5[7][25] , \g5[7][24] , \g5[7][23] , \g5[7][22] , \g5[7][21] , 
        \g5[7][20] , \g5[7][19] , \g5[7][18] , \g5[7][17] , \g5[7][16] , 
        \g5[7][15] , \g5[7][14] , \g5[7][13] , \g5[7][12] , \g5[7][11] , 
        \g5[7][10] , \g5[7][9] , \g5[7][8] , \g5[7][7] , \g5[7][6] , 
        \g5[7][5] , \g5[7][4] , \g5[7][3] , \g5[7][2] , \g5[7][1] , 
        SYNOPSYS_UNCONNECTED__53}) );
  FullAdder F0 ( .a({\g5[0][63] , \g5[0][62] , \g5[0][61] , \g5[0][60] , 
        \g5[0][59] , \g5[0][58] , \g5[0][57] , \g5[0][56] , \g5[0][55] , 
        \g5[0][54] , \g5[0][53] , \g5[0][52] , \g5[0][51] , \g5[0][50] , 
        \g5[0][49] , \g5[0][48] , \g5[0][47] , \g5[0][46] , \g5[0][45] , 
        \g5[0][44] , \g5[0][43] , \g5[0][42] , \g5[0][41] , \g5[0][40] , 
        \g5[0][39] , \g5[0][38] , \g5[0][37] , \g5[0][36] , \g5[0][35] , 
        \g5[0][34] , \g5[0][33] , \g5[0][32] , \g5[0][31] , \g5[0][30] , 
        \g5[0][29] , \g5[0][28] , \g5[0][27] , \g5[0][26] , \g5[0][25] , 
        \g5[0][24] , \g5[0][23] , \g5[0][22] , \g5[0][21] , \g5[0][20] , 
        \g5[0][19] , \g5[0][18] , \g5[0][17] , \g5[0][16] , \g5[0][15] , 
        \g5[0][14] , \g5[0][13] , \g5[0][12] , \g5[0][11] , \g5[0][10] , 
        \g5[0][9] , \g5[0][8] , \g5[0][7] , \g5[0][6] , \g5[0][5] , \g5[0][4] , 
        \g5[0][3] , \g5[0][2] , \g5[0][1] , \g5[0][0] }), .b({\g5[1][63] , 
        \g5[1][62] , \g5[1][61] , \g5[1][60] , \g5[1][59] , \g5[1][58] , 
        \g5[1][57] , \g5[1][56] , \g5[1][55] , \g5[1][54] , \g5[1][53] , 
        \g5[1][52] , \g5[1][51] , \g5[1][50] , \g5[1][49] , \g5[1][48] , 
        \g5[1][47] , \g5[1][46] , \g5[1][45] , \g5[1][44] , \g5[1][43] , 
        \g5[1][42] , \g5[1][41] , \g5[1][40] , \g5[1][39] , \g5[1][38] , 
        \g5[1][37] , \g5[1][36] , \g5[1][35] , \g5[1][34] , \g5[1][33] , 
        \g5[1][32] , \g5[1][31] , \g5[1][30] , \g5[1][29] , \g5[1][28] , 
        \g5[1][27] , \g5[1][26] , \g5[1][25] , \g5[1][24] , \g5[1][23] , 
        \g5[1][22] , \g5[1][21] , \g5[1][20] , \g5[1][19] , \g5[1][18] , 
        \g5[1][17] , \g5[1][16] , \g5[1][15] , \g5[1][14] , \g5[1][13] , 
        \g5[1][12] , \g5[1][11] , \g5[1][10] , \g5[1][9] , \g5[1][8] , 
        \g5[1][7] , \g5[1][6] , \g5[1][5] , \g5[1][4] , \g5[1][3] , \g5[1][2] , 
        \g5[1][1] , \g5[1][0] }), .cin({\g5[2][63] , \g5[2][62] , \g5[2][61] , 
        \g5[2][60] , \g5[2][59] , \g5[2][58] , \g5[2][57] , \g5[2][56] , 
        \g5[2][55] , \g5[2][54] , \g5[2][53] , \g5[2][52] , \g5[2][51] , 
        \g5[2][50] , \g5[2][49] , \g5[2][48] , \g5[2][47] , \g5[2][46] , 
        \g5[2][45] , \g5[2][44] , \g5[2][43] , \g5[2][42] , \g5[2][41] , 
        \g5[2][40] , \g5[2][39] , \g5[2][38] , \g5[2][37] , \g5[2][36] , 
        \g5[2][35] , \g5[2][34] , \g5[2][33] , \g5[2][32] , \g5[2][31] , 
        \g5[2][30] , \g5[2][29] , \g5[2][28] , \g5[2][27] , \g5[2][26] , 
        \g5[2][25] , \g5[2][24] , \g5[2][23] , \g5[2][22] , \g5[2][21] , 
        \g5[2][20] , \g5[2][19] , \g5[2][18] , \g5[2][17] , \g5[2][16] , 
        \g5[2][15] , \g5[2][14] , \g5[2][13] , \g5[2][12] , \g5[2][11] , 
        \g5[2][10] , \g5[2][9] , \g5[2][8] , \g5[2][7] , \g5[2][6] , 
        \g5[2][5] , \g5[2][4] , \g5[2][3] , \g5[2][2] , \g5[2][1] , \g5[2][0] }), .sum({\g6[0][63] , \g6[0][62] , \g6[0][61] , \g6[0][60] , \g6[0][59] , 
        \g6[0][58] , \g6[0][57] , \g6[0][56] , \g6[0][55] , \g6[0][54] , 
        \g6[0][53] , \g6[0][52] , \g6[0][51] , \g6[0][50] , \g6[0][49] , 
        \g6[0][48] , \g6[0][47] , \g6[0][46] , \g6[0][45] , \g6[0][44] , 
        \g6[0][43] , \g6[0][42] , \g6[0][41] , \g6[0][40] , \g6[0][39] , 
        \g6[0][38] , \g6[0][37] , \g6[0][36] , \g6[0][35] , \g6[0][34] , 
        \g6[0][33] , \g6[0][32] , \g6[0][31] , \g6[0][30] , \g6[0][29] , 
        \g6[0][28] , \g6[0][27] , \g6[0][26] , \g6[0][25] , \g6[0][24] , 
        \g6[0][23] , \g6[0][22] , \g6[0][21] , \g6[0][20] , \g6[0][19] , 
        \g6[0][18] , \g6[0][17] , \g6[0][16] , \g6[0][15] , \g6[0][14] , 
        \g6[0][13] , \g6[0][12] , \g6[0][11] , \g6[0][10] , \g6[0][9] , 
        \g6[0][8] , \g6[0][7] , \g6[0][6] , \g6[0][5] , \g6[0][4] , \g6[0][3] , 
        \g6[0][2] , \g6[0][1] , \g6[0][0] }), .cout({\g6[1][63] , \g6[1][62] , 
        \g6[1][61] , \g6[1][60] , \g6[1][59] , \g6[1][58] , \g6[1][57] , 
        \g6[1][56] , \g6[1][55] , \g6[1][54] , \g6[1][53] , \g6[1][52] , 
        \g6[1][51] , \g6[1][50] , \g6[1][49] , \g6[1][48] , \g6[1][47] , 
        \g6[1][46] , \g6[1][45] , \g6[1][44] , \g6[1][43] , \g6[1][42] , 
        \g6[1][41] , \g6[1][40] , \g6[1][39] , \g6[1][38] , \g6[1][37] , 
        \g6[1][36] , \g6[1][35] , \g6[1][34] , \g6[1][33] , \g6[1][32] , 
        \g6[1][31] , \g6[1][30] , \g6[1][29] , \g6[1][28] , \g6[1][27] , 
        \g6[1][26] , \g6[1][25] , \g6[1][24] , \g6[1][23] , \g6[1][22] , 
        \g6[1][21] , \g6[1][20] , \g6[1][19] , \g6[1][18] , \g6[1][17] , 
        \g6[1][16] , \g6[1][15] , \g6[1][14] , \g6[1][13] , \g6[1][12] , 
        \g6[1][11] , \g6[1][10] , \g6[1][9] , \g6[1][8] , \g6[1][7] , 
        \g6[1][6] , \g6[1][5] , \g6[1][4] , \g6[1][3] , \g6[1][2] , \g6[1][1] , 
        SYNOPSYS_UNCONNECTED__54}) );
  FullAdder F1 ( .a({\g5[3][63] , \g5[3][62] , \g5[3][61] , \g5[3][60] , 
        \g5[3][59] , \g5[3][58] , \g5[3][57] , \g5[3][56] , \g5[3][55] , 
        \g5[3][54] , \g5[3][53] , \g5[3][52] , \g5[3][51] , \g5[3][50] , 
        \g5[3][49] , \g5[3][48] , \g5[3][47] , \g5[3][46] , \g5[3][45] , 
        \g5[3][44] , \g5[3][43] , \g5[3][42] , \g5[3][41] , \g5[3][40] , 
        \g5[3][39] , \g5[3][38] , \g5[3][37] , \g5[3][36] , \g5[3][35] , 
        \g5[3][34] , \g5[3][33] , \g5[3][32] , \g5[3][31] , \g5[3][30] , 
        \g5[3][29] , \g5[3][28] , \g5[3][27] , \g5[3][26] , \g5[3][25] , 
        \g5[3][24] , \g5[3][23] , \g5[3][22] , \g5[3][21] , \g5[3][20] , 
        \g5[3][19] , \g5[3][18] , \g5[3][17] , \g5[3][16] , \g5[3][15] , 
        \g5[3][14] , \g5[3][13] , \g5[3][12] , \g5[3][11] , \g5[3][10] , 
        \g5[3][9] , \g5[3][8] , \g5[3][7] , \g5[3][6] , \g5[3][5] , \g5[3][4] , 
        \g5[3][3] , \g5[3][2] , \g5[3][1] , \g5[3][0] }), .b({\g5[4][63] , 
        \g5[4][62] , \g5[4][61] , \g5[4][60] , \g5[4][59] , \g5[4][58] , 
        \g5[4][57] , \g5[4][56] , \g5[4][55] , \g5[4][54] , \g5[4][53] , 
        \g5[4][52] , \g5[4][51] , \g5[4][50] , \g5[4][49] , \g5[4][48] , 
        \g5[4][47] , \g5[4][46] , \g5[4][45] , \g5[4][44] , \g5[4][43] , 
        \g5[4][42] , \g5[4][41] , \g5[4][40] , \g5[4][39] , \g5[4][38] , 
        \g5[4][37] , \g5[4][36] , \g5[4][35] , \g5[4][34] , \g5[4][33] , 
        \g5[4][32] , \g5[4][31] , \g5[4][30] , \g5[4][29] , \g5[4][28] , 
        \g5[4][27] , \g5[4][26] , \g5[4][25] , \g5[4][24] , \g5[4][23] , 
        \g5[4][22] , \g5[4][21] , \g5[4][20] , \g5[4][19] , \g5[4][18] , 
        \g5[4][17] , \g5[4][16] , \g5[4][15] , \g5[4][14] , \g5[4][13] , 
        \g5[4][12] , \g5[4][11] , \g5[4][10] , \g5[4][9] , \g5[4][8] , 
        \g5[4][7] , \g5[4][6] , \g5[4][5] , \g5[4][4] , \g5[4][3] , \g5[4][2] , 
        \g5[4][1] , 1'b0}), .cin({\g5[5][63] , \g5[5][62] , \g5[5][61] , 
        \g5[5][60] , \g5[5][59] , \g5[5][58] , \g5[5][57] , \g5[5][56] , 
        \g5[5][55] , \g5[5][54] , \g5[5][53] , \g5[5][52] , \g5[5][51] , 
        \g5[5][50] , \g5[5][49] , \g5[5][48] , \g5[5][47] , \g5[5][46] , 
        \g5[5][45] , \g5[5][44] , \g5[5][43] , \g5[5][42] , \g5[5][41] , 
        \g5[5][40] , \g5[5][39] , \g5[5][38] , \g5[5][37] , \g5[5][36] , 
        \g5[5][35] , \g5[5][34] , \g5[5][33] , \g5[5][32] , \g5[5][31] , 
        \g5[5][30] , \g5[5][29] , \g5[5][28] , \g5[5][27] , \g5[5][26] , 
        \g5[5][25] , \g5[5][24] , \g5[5][23] , \g5[5][22] , \g5[5][21] , 
        \g5[5][20] , \g5[5][19] , \g5[5][18] , \g5[5][17] , \g5[5][16] , 
        \g5[5][15] , \g5[5][14] , \g5[5][13] , \g5[5][12] , \g5[5][11] , 
        \g5[5][10] , \g5[5][9] , \g5[5][8] , \g5[5][7] , \g5[5][6] , 
        \g5[5][5] , \g5[5][4] , \g5[5][3] , \g5[5][2] , \g5[5][1] , 1'b0}), 
        .sum({\g6[2][63] , \g6[2][62] , \g6[2][61] , \g6[2][60] , \g6[2][59] , 
        \g6[2][58] , \g6[2][57] , \g6[2][56] , \g6[2][55] , \g6[2][54] , 
        \g6[2][53] , \g6[2][52] , \g6[2][51] , \g6[2][50] , \g6[2][49] , 
        \g6[2][48] , \g6[2][47] , \g6[2][46] , \g6[2][45] , \g6[2][44] , 
        \g6[2][43] , \g6[2][42] , \g6[2][41] , \g6[2][40] , \g6[2][39] , 
        \g6[2][38] , \g6[2][37] , \g6[2][36] , \g6[2][35] , \g6[2][34] , 
        \g6[2][33] , \g6[2][32] , \g6[2][31] , \g6[2][30] , \g6[2][29] , 
        \g6[2][28] , \g6[2][27] , \g6[2][26] , \g6[2][25] , \g6[2][24] , 
        \g6[2][23] , \g6[2][22] , \g6[2][21] , \g6[2][20] , \g6[2][19] , 
        \g6[2][18] , \g6[2][17] , \g6[2][16] , \g6[2][15] , \g6[2][14] , 
        \g6[2][13] , \g6[2][12] , \g6[2][11] , \g6[2][10] , \g6[2][9] , 
        \g6[2][8] , \g6[2][7] , \g6[2][6] , \g6[2][5] , \g6[2][4] , \g6[2][3] , 
        \g6[2][2] , \g6[2][1] , \g6[2][0] }), .cout({\g6[3][63] , \g6[3][62] , 
        \g6[3][61] , \g6[3][60] , \g6[3][59] , \g6[3][58] , \g6[3][57] , 
        \g6[3][56] , \g6[3][55] , \g6[3][54] , \g6[3][53] , \g6[3][52] , 
        \g6[3][51] , \g6[3][50] , \g6[3][49] , \g6[3][48] , \g6[3][47] , 
        \g6[3][46] , \g6[3][45] , \g6[3][44] , \g6[3][43] , \g6[3][42] , 
        \g6[3][41] , \g6[3][40] , \g6[3][39] , \g6[3][38] , \g6[3][37] , 
        \g6[3][36] , \g6[3][35] , \g6[3][34] , \g6[3][33] , \g6[3][32] , 
        \g6[3][31] , \g6[3][30] , \g6[3][29] , \g6[3][28] , \g6[3][27] , 
        \g6[3][26] , \g6[3][25] , \g6[3][24] , \g6[3][23] , \g6[3][22] , 
        \g6[3][21] , \g6[3][20] , \g6[3][19] , \g6[3][18] , \g6[3][17] , 
        \g6[3][16] , \g6[3][15] , \g6[3][14] , \g6[3][13] , \g6[3][12] , 
        \g6[3][11] , \g6[3][10] , \g6[3][9] , \g6[3][8] , \g6[3][7] , 
        \g6[3][6] , \g6[3][5] , \g6[3][4] , \g6[3][3] , \g6[3][2] , \g6[3][1] , 
        SYNOPSYS_UNCONNECTED__55}) );
  FullAdder F2 ( .a({\g5[6][63] , \g5[6][62] , \g5[6][61] , \g5[6][60] , 
        \g5[6][59] , \g5[6][58] , \g5[6][57] , \g5[6][56] , \g5[6][55] , 
        \g5[6][54] , \g5[6][53] , \g5[6][52] , \g5[6][51] , \g5[6][50] , 
        \g5[6][49] , \g5[6][48] , \g5[6][47] , \g5[6][46] , \g5[6][45] , 
        \g5[6][44] , \g5[6][43] , \g5[6][42] , \g5[6][41] , \g5[6][40] , 
        \g5[6][39] , \g5[6][38] , \g5[6][37] , \g5[6][36] , \g5[6][35] , 
        \g5[6][34] , \g5[6][33] , \g5[6][32] , \g5[6][31] , \g5[6][30] , 
        \g5[6][29] , \g5[6][28] , \g5[6][27] , \g5[6][26] , \g5[6][25] , 
        \g5[6][24] , \g5[6][23] , \g5[6][22] , \g5[6][21] , \g5[6][20] , 
        \g5[6][19] , \g5[6][18] , \g5[6][17] , \g5[6][16] , \g5[6][15] , 
        \g5[6][14] , \g5[6][13] , \g5[6][12] , \g5[6][11] , \g5[6][10] , 
        \g5[6][9] , \g5[6][8] , \g5[6][7] , \g5[6][6] , \g5[6][5] , \g5[6][4] , 
        \g5[6][3] , \g5[6][2] , \g5[6][1] , 1'b0}), .b({\g5[7][63] , 
        \g5[7][62] , \g5[7][61] , \g5[7][60] , \g5[7][59] , \g5[7][58] , 
        \g5[7][57] , \g5[7][56] , \g5[7][55] , \g5[7][54] , \g5[7][53] , 
        \g5[7][52] , \g5[7][51] , \g5[7][50] , \g5[7][49] , \g5[7][48] , 
        \g5[7][47] , \g5[7][46] , \g5[7][45] , \g5[7][44] , \g5[7][43] , 
        \g5[7][42] , \g5[7][41] , \g5[7][40] , \g5[7][39] , \g5[7][38] , 
        \g5[7][37] , \g5[7][36] , \g5[7][35] , \g5[7][34] , \g5[7][33] , 
        \g5[7][32] , \g5[7][31] , \g5[7][30] , \g5[7][29] , \g5[7][28] , 
        \g5[7][27] , \g5[7][26] , \g5[7][25] , \g5[7][24] , \g5[7][23] , 
        \g5[7][22] , \g5[7][21] , \g5[7][20] , \g5[7][19] , \g5[7][18] , 
        \g5[7][17] , \g5[7][16] , \g5[7][15] , \g5[7][14] , \g5[7][13] , 
        \g5[7][12] , \g5[7][11] , \g5[7][10] , \g5[7][9] , \g5[7][8] , 
        \g5[7][7] , \g5[7][6] , \g5[7][5] , \g5[7][4] , \g5[7][3] , \g5[7][2] , 
        \g5[7][1] , 1'b0}), .cin({\g2[27][63] , \g2[27][62] , \g2[27][61] , 
        \g2[27][60] , \g2[27][59] , \g2[27][58] , \g2[27][57] , \g2[27][56] , 
        \g2[27][55] , \g2[27][54] , \g2[27][53] , \g2[27][52] , \g2[27][51] , 
        \g2[27][50] , \g2[27][49] , \g2[27][48] , \g2[27][47] , \g2[27][46] , 
        \g2[27][45] , \g2[27][44] , \g2[27][43] , \g2[27][42] , \g2[27][41] , 
        \g2[27][40] , \g2[27][39] , \g2[27][38] , \g2[27][37] , \g2[27][36] , 
        \g2[27][35] , \g2[27][34] , \g2[27][33] , \g2[27][32] , \g2[27][31] , 
        \g2[27][30] , \g2[27][29] , \g2[27][28] , \g2[27][27] , \g2[27][26] , 
        \g2[27][25] , \g2[27][24] , \g2[27][23] , \g2[27][22] , \g2[27][21] , 
        \g2[27][20] , \g2[27][19] , \g2[27][18] , \g2[27][17] , \g2[27][16] , 
        \g2[27][15] , \g2[27][14] , \g2[27][13] , \g2[27][12] , \g2[27][11] , 
        \g2[27][10] , \g2[27][9] , \g2[27][8] , \g2[27][7] , \g2[27][6] , 
        \g2[27][5] , \g2[27][4] , \g2[27][3] , \g2[27][2] , \g2[27][1] , 1'b0}), .sum({\g6[4][63] , \g6[4][62] , \g6[4][61] , \g6[4][60] , \g6[4][59] , 
        \g6[4][58] , \g6[4][57] , \g6[4][56] , \g6[4][55] , \g6[4][54] , 
        \g6[4][53] , \g6[4][52] , \g6[4][51] , \g6[4][50] , \g6[4][49] , 
        \g6[4][48] , \g6[4][47] , \g6[4][46] , \g6[4][45] , \g6[4][44] , 
        \g6[4][43] , \g6[4][42] , \g6[4][41] , \g6[4][40] , \g6[4][39] , 
        \g6[4][38] , \g6[4][37] , \g6[4][36] , \g6[4][35] , \g6[4][34] , 
        \g6[4][33] , \g6[4][32] , \g6[4][31] , \g6[4][30] , \g6[4][29] , 
        \g6[4][28] , \g6[4][27] , \g6[4][26] , \g6[4][25] , \g6[4][24] , 
        \g6[4][23] , \g6[4][22] , \g6[4][21] , \g6[4][20] , \g6[4][19] , 
        \g6[4][18] , \g6[4][17] , \g6[4][16] , \g6[4][15] , \g6[4][14] , 
        \g6[4][13] , \g6[4][12] , \g6[4][11] , \g6[4][10] , \g6[4][9] , 
        \g6[4][8] , \g6[4][7] , \g6[4][6] , \g6[4][5] , \g6[4][4] , \g6[4][3] , 
        \g6[4][2] , \g6[4][1] , \g6[4][0] }), .cout({\g6[5][63] , \g6[5][62] , 
        \g6[5][61] , \g6[5][60] , \g6[5][59] , \g6[5][58] , \g6[5][57] , 
        \g6[5][56] , \g6[5][55] , \g6[5][54] , \g6[5][53] , \g6[5][52] , 
        \g6[5][51] , \g6[5][50] , \g6[5][49] , \g6[5][48] , \g6[5][47] , 
        \g6[5][46] , \g6[5][45] , \g6[5][44] , \g6[5][43] , \g6[5][42] , 
        \g6[5][41] , \g6[5][40] , \g6[5][39] , \g6[5][38] , \g6[5][37] , 
        \g6[5][36] , \g6[5][35] , \g6[5][34] , \g6[5][33] , \g6[5][32] , 
        \g6[5][31] , \g6[5][30] , \g6[5][29] , \g6[5][28] , \g6[5][27] , 
        \g6[5][26] , \g6[5][25] , \g6[5][24] , \g6[5][23] , \g6[5][22] , 
        \g6[5][21] , \g6[5][20] , \g6[5][19] , \g6[5][18] , \g6[5][17] , 
        \g6[5][16] , \g6[5][15] , \g6[5][14] , \g6[5][13] , \g6[5][12] , 
        \g6[5][11] , \g6[5][10] , \g6[5][9] , \g6[5][8] , \g6[5][7] , 
        \g6[5][6] , \g6[5][5] , \g6[5][4] , \g6[5][3] , \g6[5][2] , \g6[5][1] , 
        SYNOPSYS_UNCONNECTED__56}) );
  FullAdder F3 ( .a({\g6[0][63] , \g6[0][62] , \g6[0][61] , \g6[0][60] , 
        \g6[0][59] , \g6[0][58] , \g6[0][57] , \g6[0][56] , \g6[0][55] , 
        \g6[0][54] , \g6[0][53] , \g6[0][52] , \g6[0][51] , \g6[0][50] , 
        \g6[0][49] , \g6[0][48] , \g6[0][47] , \g6[0][46] , \g6[0][45] , 
        \g6[0][44] , \g6[0][43] , \g6[0][42] , \g6[0][41] , \g6[0][40] , 
        \g6[0][39] , \g6[0][38] , \g6[0][37] , \g6[0][36] , \g6[0][35] , 
        \g6[0][34] , \g6[0][33] , \g6[0][32] , \g6[0][31] , \g6[0][30] , 
        \g6[0][29] , \g6[0][28] , \g6[0][27] , \g6[0][26] , \g6[0][25] , 
        \g6[0][24] , \g6[0][23] , \g6[0][22] , \g6[0][21] , \g6[0][20] , 
        \g6[0][19] , \g6[0][18] , \g6[0][17] , \g6[0][16] , \g6[0][15] , 
        \g6[0][14] , \g6[0][13] , \g6[0][12] , \g6[0][11] , \g6[0][10] , 
        \g6[0][9] , \g6[0][8] , \g6[0][7] , \g6[0][6] , \g6[0][5] , \g6[0][4] , 
        \g6[0][3] , \g6[0][2] , \g6[0][1] , \g6[0][0] }), .b({\g6[1][63] , 
        \g6[1][62] , \g6[1][61] , \g6[1][60] , \g6[1][59] , \g6[1][58] , 
        \g6[1][57] , \g6[1][56] , \g6[1][55] , \g6[1][54] , \g6[1][53] , 
        \g6[1][52] , \g6[1][51] , \g6[1][50] , \g6[1][49] , \g6[1][48] , 
        \g6[1][47] , \g6[1][46] , \g6[1][45] , \g6[1][44] , \g6[1][43] , 
        \g6[1][42] , \g6[1][41] , \g6[1][40] , \g6[1][39] , \g6[1][38] , 
        \g6[1][37] , \g6[1][36] , \g6[1][35] , \g6[1][34] , \g6[1][33] , 
        \g6[1][32] , \g6[1][31] , \g6[1][30] , \g6[1][29] , \g6[1][28] , 
        \g6[1][27] , \g6[1][26] , \g6[1][25] , \g6[1][24] , \g6[1][23] , 
        \g6[1][22] , \g6[1][21] , \g6[1][20] , \g6[1][19] , \g6[1][18] , 
        \g6[1][17] , \g6[1][16] , \g6[1][15] , \g6[1][14] , \g6[1][13] , 
        \g6[1][12] , \g6[1][11] , \g6[1][10] , \g6[1][9] , \g6[1][8] , 
        \g6[1][7] , \g6[1][6] , \g6[1][5] , \g6[1][4] , \g6[1][3] , \g6[1][2] , 
        \g6[1][1] , 1'b0}), .cin({\g6[2][63] , \g6[2][62] , \g6[2][61] , 
        \g6[2][60] , \g6[2][59] , \g6[2][58] , \g6[2][57] , \g6[2][56] , 
        \g6[2][55] , \g6[2][54] , \g6[2][53] , \g6[2][52] , \g6[2][51] , 
        \g6[2][50] , \g6[2][49] , \g6[2][48] , \g6[2][47] , \g6[2][46] , 
        \g6[2][45] , \g6[2][44] , \g6[2][43] , \g6[2][42] , \g6[2][41] , 
        \g6[2][40] , \g6[2][39] , \g6[2][38] , \g6[2][37] , \g6[2][36] , 
        \g6[2][35] , \g6[2][34] , \g6[2][33] , \g6[2][32] , \g6[2][31] , 
        \g6[2][30] , \g6[2][29] , \g6[2][28] , \g6[2][27] , \g6[2][26] , 
        \g6[2][25] , \g6[2][24] , \g6[2][23] , \g6[2][22] , \g6[2][21] , 
        \g6[2][20] , \g6[2][19] , \g6[2][18] , \g6[2][17] , \g6[2][16] , 
        \g6[2][15] , \g6[2][14] , \g6[2][13] , \g6[2][12] , \g6[2][11] , 
        \g6[2][10] , \g6[2][9] , \g6[2][8] , \g6[2][7] , \g6[2][6] , 
        \g6[2][5] , \g6[2][4] , \g6[2][3] , \g6[2][2] , \g6[2][1] , \g6[2][0] }), .sum({\g7[0][63] , \g7[0][62] , \g7[0][61] , \g7[0][60] , \g7[0][59] , 
        \g7[0][58] , \g7[0][57] , \g7[0][56] , \g7[0][55] , \g7[0][54] , 
        \g7[0][53] , \g7[0][52] , \g7[0][51] , \g7[0][50] , \g7[0][49] , 
        \g7[0][48] , \g7[0][47] , \g7[0][46] , \g7[0][45] , \g7[0][44] , 
        \g7[0][43] , \g7[0][42] , \g7[0][41] , \g7[0][40] , \g7[0][39] , 
        \g7[0][38] , \g7[0][37] , \g7[0][36] , \g7[0][35] , \g7[0][34] , 
        \g7[0][33] , \g7[0][32] , \g7[0][31] , \g7[0][30] , \g7[0][29] , 
        \g7[0][28] , \g7[0][27] , \g7[0][26] , \g7[0][25] , \g7[0][24] , 
        \g7[0][23] , \g7[0][22] , \g7[0][21] , \g7[0][20] , \g7[0][19] , 
        \g7[0][18] , \g7[0][17] , \g7[0][16] , \g7[0][15] , \g7[0][14] , 
        \g7[0][13] , \g7[0][12] , \g7[0][11] , \g7[0][10] , \g7[0][9] , 
        \g7[0][8] , \g7[0][7] , \g7[0][6] , \g7[0][5] , \g7[0][4] , \g7[0][3] , 
        \g7[0][2] , \g7[0][1] , \g7[0][0] }), .cout({\g7[1][63] , \g7[1][62] , 
        \g7[1][61] , \g7[1][60] , \g7[1][59] , \g7[1][58] , \g7[1][57] , 
        \g7[1][56] , \g7[1][55] , \g7[1][54] , \g7[1][53] , \g7[1][52] , 
        \g7[1][51] , \g7[1][50] , \g7[1][49] , \g7[1][48] , \g7[1][47] , 
        \g7[1][46] , \g7[1][45] , \g7[1][44] , \g7[1][43] , \g7[1][42] , 
        \g7[1][41] , \g7[1][40] , \g7[1][39] , \g7[1][38] , \g7[1][37] , 
        \g7[1][36] , \g7[1][35] , \g7[1][34] , \g7[1][33] , \g7[1][32] , 
        \g7[1][31] , \g7[1][30] , \g7[1][29] , \g7[1][28] , \g7[1][27] , 
        \g7[1][26] , \g7[1][25] , \g7[1][24] , \g7[1][23] , \g7[1][22] , 
        \g7[1][21] , \g7[1][20] , \g7[1][19] , \g7[1][18] , \g7[1][17] , 
        \g7[1][16] , \g7[1][15] , \g7[1][14] , \g7[1][13] , \g7[1][12] , 
        \g7[1][11] , \g7[1][10] , \g7[1][9] , \g7[1][8] , \g7[1][7] , 
        \g7[1][6] , \g7[1][5] , \g7[1][4] , \g7[1][3] , \g7[1][2] , \g7[1][1] , 
        SYNOPSYS_UNCONNECTED__57}) );
  FullAdder F4 ( .a({\g6[3][63] , \g6[3][62] , \g6[3][61] , \g6[3][60] , 
        \g6[3][59] , \g6[3][58] , \g6[3][57] , \g6[3][56] , \g6[3][55] , 
        \g6[3][54] , \g6[3][53] , \g6[3][52] , \g6[3][51] , \g6[3][50] , 
        \g6[3][49] , \g6[3][48] , \g6[3][47] , \g6[3][46] , \g6[3][45] , 
        \g6[3][44] , \g6[3][43] , \g6[3][42] , \g6[3][41] , \g6[3][40] , 
        \g6[3][39] , \g6[3][38] , \g6[3][37] , \g6[3][36] , \g6[3][35] , 
        \g6[3][34] , \g6[3][33] , \g6[3][32] , \g6[3][31] , \g6[3][30] , 
        \g6[3][29] , \g6[3][28] , \g6[3][27] , \g6[3][26] , \g6[3][25] , 
        \g6[3][24] , \g6[3][23] , \g6[3][22] , \g6[3][21] , \g6[3][20] , 
        \g6[3][19] , \g6[3][18] , \g6[3][17] , \g6[3][16] , \g6[3][15] , 
        \g6[3][14] , \g6[3][13] , \g6[3][12] , \g6[3][11] , \g6[3][10] , 
        \g6[3][9] , \g6[3][8] , \g6[3][7] , \g6[3][6] , \g6[3][5] , \g6[3][4] , 
        \g6[3][3] , \g6[3][2] , \g6[3][1] , 1'b0}), .b({\g6[4][63] , 
        \g6[4][62] , \g6[4][61] , \g6[4][60] , \g6[4][59] , \g6[4][58] , 
        \g6[4][57] , \g6[4][56] , \g6[4][55] , \g6[4][54] , \g6[4][53] , 
        \g6[4][52] , \g6[4][51] , \g6[4][50] , \g6[4][49] , \g6[4][48] , 
        \g6[4][47] , \g6[4][46] , \g6[4][45] , \g6[4][44] , \g6[4][43] , 
        \g6[4][42] , \g6[4][41] , \g6[4][40] , \g6[4][39] , \g6[4][38] , 
        \g6[4][37] , \g6[4][36] , \g6[4][35] , \g6[4][34] , \g6[4][33] , 
        \g6[4][32] , \g6[4][31] , \g6[4][30] , \g6[4][29] , \g6[4][28] , 
        \g6[4][27] , \g6[4][26] , \g6[4][25] , \g6[4][24] , \g6[4][23] , 
        \g6[4][22] , \g6[4][21] , \g6[4][20] , \g6[4][19] , \g6[4][18] , 
        \g6[4][17] , \g6[4][16] , \g6[4][15] , \g6[4][14] , \g6[4][13] , 
        \g6[4][12] , \g6[4][11] , \g6[4][10] , \g6[4][9] , \g6[4][8] , 
        \g6[4][7] , \g6[4][6] , \g6[4][5] , \g6[4][4] , \g6[4][3] , \g6[4][2] , 
        \g6[4][1] , \g6[4][0] }), .cin({\g6[5][63] , \g6[5][62] , \g6[5][61] , 
        \g6[5][60] , \g6[5][59] , \g6[5][58] , \g6[5][57] , \g6[5][56] , 
        \g6[5][55] , \g6[5][54] , \g6[5][53] , \g6[5][52] , \g6[5][51] , 
        \g6[5][50] , \g6[5][49] , \g6[5][48] , \g6[5][47] , \g6[5][46] , 
        \g6[5][45] , \g6[5][44] , \g6[5][43] , \g6[5][42] , \g6[5][41] , 
        \g6[5][40] , \g6[5][39] , \g6[5][38] , \g6[5][37] , \g6[5][36] , 
        \g6[5][35] , \g6[5][34] , \g6[5][33] , \g6[5][32] , \g6[5][31] , 
        \g6[5][30] , \g6[5][29] , \g6[5][28] , \g6[5][27] , \g6[5][26] , 
        \g6[5][25] , \g6[5][24] , \g6[5][23] , \g6[5][22] , \g6[5][21] , 
        \g6[5][20] , \g6[5][19] , \g6[5][18] , \g6[5][17] , \g6[5][16] , 
        \g6[5][15] , \g6[5][14] , \g6[5][13] , \g6[5][12] , \g6[5][11] , 
        \g6[5][10] , \g6[5][9] , \g6[5][8] , \g6[5][7] , \g6[5][6] , 
        \g6[5][5] , \g6[5][4] , \g6[5][3] , \g6[5][2] , \g6[5][1] , 1'b0}), 
        .sum({\g7[2][63] , \g7[2][62] , \g7[2][61] , \g7[2][60] , \g7[2][59] , 
        \g7[2][58] , \g7[2][57] , \g7[2][56] , \g7[2][55] , \g7[2][54] , 
        \g7[2][53] , \g7[2][52] , \g7[2][51] , \g7[2][50] , \g7[2][49] , 
        \g7[2][48] , \g7[2][47] , \g7[2][46] , \g7[2][45] , \g7[2][44] , 
        \g7[2][43] , \g7[2][42] , \g7[2][41] , \g7[2][40] , \g7[2][39] , 
        \g7[2][38] , \g7[2][37] , \g7[2][36] , \g7[2][35] , \g7[2][34] , 
        \g7[2][33] , \g7[2][32] , \g7[2][31] , \g7[2][30] , \g7[2][29] , 
        \g7[2][28] , \g7[2][27] , \g7[2][26] , \g7[2][25] , \g7[2][24] , 
        \g7[2][23] , \g7[2][22] , \g7[2][21] , \g7[2][20] , \g7[2][19] , 
        \g7[2][18] , \g7[2][17] , \g7[2][16] , \g7[2][15] , \g7[2][14] , 
        \g7[2][13] , \g7[2][12] , \g7[2][11] , \g7[2][10] , \g7[2][9] , 
        \g7[2][8] , \g7[2][7] , \g7[2][6] , \g7[2][5] , \g7[2][4] , \g7[2][3] , 
        \g7[2][2] , \g7[2][1] , \g7[2][0] }), .cout({\g7[3][63] , \g7[3][62] , 
        \g7[3][61] , \g7[3][60] , \g7[3][59] , \g7[3][58] , \g7[3][57] , 
        \g7[3][56] , \g7[3][55] , \g7[3][54] , \g7[3][53] , \g7[3][52] , 
        \g7[3][51] , \g7[3][50] , \g7[3][49] , \g7[3][48] , \g7[3][47] , 
        \g7[3][46] , \g7[3][45] , \g7[3][44] , \g7[3][43] , \g7[3][42] , 
        \g7[3][41] , \g7[3][40] , \g7[3][39] , \g7[3][38] , \g7[3][37] , 
        \g7[3][36] , \g7[3][35] , \g7[3][34] , \g7[3][33] , \g7[3][32] , 
        \g7[3][31] , \g7[3][30] , \g7[3][29] , \g7[3][28] , \g7[3][27] , 
        \g7[3][26] , \g7[3][25] , \g7[3][24] , \g7[3][23] , \g7[3][22] , 
        \g7[3][21] , \g7[3][20] , \g7[3][19] , \g7[3][18] , \g7[3][17] , 
        \g7[3][16] , \g7[3][15] , \g7[3][14] , \g7[3][13] , \g7[3][12] , 
        \g7[3][11] , \g7[3][10] , \g7[3][9] , \g7[3][8] , \g7[3][7] , 
        \g7[3][6] , \g7[3][5] , \g7[3][4] , \g7[3][3] , \g7[3][2] , \g7[3][1] , 
        SYNOPSYS_UNCONNECTED__58}) );
  FullAdder F5 ( .a({\g7[0][63] , \g7[0][62] , \g7[0][61] , \g7[0][60] , 
        \g7[0][59] , \g7[0][58] , \g7[0][57] , \g7[0][56] , \g7[0][55] , 
        \g7[0][54] , \g7[0][53] , \g7[0][52] , \g7[0][51] , \g7[0][50] , 
        \g7[0][49] , \g7[0][48] , \g7[0][47] , \g7[0][46] , \g7[0][45] , 
        \g7[0][44] , \g7[0][43] , \g7[0][42] , \g7[0][41] , \g7[0][40] , 
        \g7[0][39] , \g7[0][38] , \g7[0][37] , \g7[0][36] , \g7[0][35] , 
        \g7[0][34] , \g7[0][33] , \g7[0][32] , \g7[0][31] , \g7[0][30] , 
        \g7[0][29] , \g7[0][28] , \g7[0][27] , \g7[0][26] , \g7[0][25] , 
        \g7[0][24] , \g7[0][23] , \g7[0][22] , \g7[0][21] , \g7[0][20] , 
        \g7[0][19] , \g7[0][18] , \g7[0][17] , \g7[0][16] , \g7[0][15] , 
        \g7[0][14] , \g7[0][13] , \g7[0][12] , \g7[0][11] , \g7[0][10] , 
        \g7[0][9] , \g7[0][8] , \g7[0][7] , \g7[0][6] , \g7[0][5] , \g7[0][4] , 
        \g7[0][3] , \g7[0][2] , \g7[0][1] , \g7[0][0] }), .b({\g7[1][63] , 
        \g7[1][62] , \g7[1][61] , \g7[1][60] , \g7[1][59] , \g7[1][58] , 
        \g7[1][57] , \g7[1][56] , \g7[1][55] , \g7[1][54] , \g7[1][53] , 
        \g7[1][52] , \g7[1][51] , \g7[1][50] , \g7[1][49] , \g7[1][48] , 
        \g7[1][47] , \g7[1][46] , \g7[1][45] , \g7[1][44] , \g7[1][43] , 
        \g7[1][42] , \g7[1][41] , \g7[1][40] , \g7[1][39] , \g7[1][38] , 
        \g7[1][37] , \g7[1][36] , \g7[1][35] , \g7[1][34] , \g7[1][33] , 
        \g7[1][32] , \g7[1][31] , \g7[1][30] , \g7[1][29] , \g7[1][28] , 
        \g7[1][27] , \g7[1][26] , \g7[1][25] , \g7[1][24] , \g7[1][23] , 
        \g7[1][22] , \g7[1][21] , \g7[1][20] , \g7[1][19] , \g7[1][18] , 
        \g7[1][17] , \g7[1][16] , \g7[1][15] , \g7[1][14] , \g7[1][13] , 
        \g7[1][12] , \g7[1][11] , \g7[1][10] , \g7[1][9] , \g7[1][8] , 
        \g7[1][7] , \g7[1][6] , \g7[1][5] , \g7[1][4] , \g7[1][3] , \g7[1][2] , 
        \g7[1][1] , 1'b0}), .cin({\g7[2][63] , \g7[2][62] , \g7[2][61] , 
        \g7[2][60] , \g7[2][59] , \g7[2][58] , \g7[2][57] , \g7[2][56] , 
        \g7[2][55] , \g7[2][54] , \g7[2][53] , \g7[2][52] , \g7[2][51] , 
        \g7[2][50] , \g7[2][49] , \g7[2][48] , \g7[2][47] , \g7[2][46] , 
        \g7[2][45] , \g7[2][44] , \g7[2][43] , \g7[2][42] , \g7[2][41] , 
        \g7[2][40] , \g7[2][39] , \g7[2][38] , \g7[2][37] , \g7[2][36] , 
        \g7[2][35] , \g7[2][34] , \g7[2][33] , \g7[2][32] , \g7[2][31] , 
        \g7[2][30] , \g7[2][29] , \g7[2][28] , \g7[2][27] , \g7[2][26] , 
        \g7[2][25] , \g7[2][24] , \g7[2][23] , \g7[2][22] , \g7[2][21] , 
        \g7[2][20] , \g7[2][19] , \g7[2][18] , \g7[2][17] , \g7[2][16] , 
        \g7[2][15] , \g7[2][14] , \g7[2][13] , \g7[2][12] , \g7[2][11] , 
        \g7[2][10] , \g7[2][9] , \g7[2][8] , \g7[2][7] , \g7[2][6] , 
        \g7[2][5] , \g7[2][4] , \g7[2][3] , \g7[2][2] , \g7[2][1] , \g7[2][0] }), .sum({\g8[0][63] , \g8[0][62] , \g8[0][61] , \g8[0][60] , \g8[0][59] , 
        \g8[0][58] , \g8[0][57] , \g8[0][56] , \g8[0][55] , \g8[0][54] , 
        \g8[0][53] , \g8[0][52] , \g8[0][51] , \g8[0][50] , \g8[0][49] , 
        \g8[0][48] , \g8[0][47] , \g8[0][46] , \g8[0][45] , \g8[0][44] , 
        \g8[0][43] , \g8[0][42] , \g8[0][41] , \g8[0][40] , \g8[0][39] , 
        \g8[0][38] , \g8[0][37] , \g8[0][36] , \g8[0][35] , \g8[0][34] , 
        \g8[0][33] , \g8[0][32] , \g8[0][31] , \g8[0][30] , \g8[0][29] , 
        \g8[0][28] , \g8[0][27] , \g8[0][26] , \g8[0][25] , \g8[0][24] , 
        \g8[0][23] , \g8[0][22] , \g8[0][21] , \g8[0][20] , \g8[0][19] , 
        \g8[0][18] , \g8[0][17] , \g8[0][16] , \g8[0][15] , \g8[0][14] , 
        \g8[0][13] , \g8[0][12] , \g8[0][11] , \g8[0][10] , \g8[0][9] , 
        \g8[0][8] , \g8[0][7] , \g8[0][6] , \g8[0][5] , \g8[0][4] , \g8[0][3] , 
        \g8[0][2] , \g8[0][1] , \g8[0][0] }), .cout({\g8[1][63] , \g8[1][62] , 
        \g8[1][61] , \g8[1][60] , \g8[1][59] , \g8[1][58] , \g8[1][57] , 
        \g8[1][56] , \g8[1][55] , \g8[1][54] , \g8[1][53] , \g8[1][52] , 
        \g8[1][51] , \g8[1][50] , \g8[1][49] , \g8[1][48] , \g8[1][47] , 
        \g8[1][46] , \g8[1][45] , \g8[1][44] , \g8[1][43] , \g8[1][42] , 
        \g8[1][41] , \g8[1][40] , \g8[1][39] , \g8[1][38] , \g8[1][37] , 
        \g8[1][36] , \g8[1][35] , \g8[1][34] , \g8[1][33] , \g8[1][32] , 
        \g8[1][31] , \g8[1][30] , \g8[1][29] , \g8[1][28] , \g8[1][27] , 
        \g8[1][26] , \g8[1][25] , \g8[1][24] , \g8[1][23] , \g8[1][22] , 
        \g8[1][21] , \g8[1][20] , \g8[1][19] , \g8[1][18] , \g8[1][17] , 
        \g8[1][16] , \g8[1][15] , \g8[1][14] , \g8[1][13] , \g8[1][12] , 
        \g8[1][11] , \g8[1][10] , \g8[1][9] , \g8[1][8] , \g8[1][7] , 
        \g8[1][6] , \g8[1][5] , \g8[1][4] , \g8[1][3] , \g8[1][2] , \g8[1][1] , 
        SYNOPSYS_UNCONNECTED__59}) );
  FullAdder F6 ( .a({\g8[0][63] , \g8[0][62] , \g8[0][61] , \g8[0][60] , 
        \g8[0][59] , \g8[0][58] , \g8[0][57] , \g8[0][56] , \g8[0][55] , 
        \g8[0][54] , \g8[0][53] , \g8[0][52] , \g8[0][51] , \g8[0][50] , 
        \g8[0][49] , \g8[0][48] , \g8[0][47] , \g8[0][46] , \g8[0][45] , 
        \g8[0][44] , \g8[0][43] , \g8[0][42] , \g8[0][41] , \g8[0][40] , 
        \g8[0][39] , \g8[0][38] , \g8[0][37] , \g8[0][36] , \g8[0][35] , 
        \g8[0][34] , \g8[0][33] , \g8[0][32] , \g8[0][31] , \g8[0][30] , 
        \g8[0][29] , \g8[0][28] , \g8[0][27] , \g8[0][26] , \g8[0][25] , 
        \g8[0][24] , \g8[0][23] , \g8[0][22] , \g8[0][21] , \g8[0][20] , 
        \g8[0][19] , \g8[0][18] , \g8[0][17] , \g8[0][16] , \g8[0][15] , 
        \g8[0][14] , \g8[0][13] , \g8[0][12] , \g8[0][11] , \g8[0][10] , 
        \g8[0][9] , \g8[0][8] , \g8[0][7] , \g8[0][6] , \g8[0][5] , \g8[0][4] , 
        \g8[0][3] , \g8[0][2] , \g8[0][1] , \g8[0][0] }), .b({\g8[1][63] , 
        \g8[1][62] , \g8[1][61] , \g8[1][60] , \g8[1][59] , \g8[1][58] , 
        \g8[1][57] , \g8[1][56] , \g8[1][55] , \g8[1][54] , \g8[1][53] , 
        \g8[1][52] , \g8[1][51] , \g8[1][50] , \g8[1][49] , \g8[1][48] , 
        \g8[1][47] , \g8[1][46] , \g8[1][45] , \g8[1][44] , \g8[1][43] , 
        \g8[1][42] , \g8[1][41] , \g8[1][40] , \g8[1][39] , \g8[1][38] , 
        \g8[1][37] , \g8[1][36] , \g8[1][35] , \g8[1][34] , \g8[1][33] , 
        \g8[1][32] , \g8[1][31] , \g8[1][30] , \g8[1][29] , \g8[1][28] , 
        \g8[1][27] , \g8[1][26] , \g8[1][25] , \g8[1][24] , \g8[1][23] , 
        \g8[1][22] , \g8[1][21] , \g8[1][20] , \g8[1][19] , \g8[1][18] , 
        \g8[1][17] , \g8[1][16] , \g8[1][15] , \g8[1][14] , \g8[1][13] , 
        \g8[1][12] , \g8[1][11] , \g8[1][10] , \g8[1][9] , \g8[1][8] , 
        \g8[1][7] , \g8[1][6] , \g8[1][5] , \g8[1][4] , \g8[1][3] , \g8[1][2] , 
        \g8[1][1] , 1'b0}), .cin({\g7[3][63] , \g7[3][62] , \g7[3][61] , 
        \g7[3][60] , \g7[3][59] , \g7[3][58] , \g7[3][57] , \g7[3][56] , 
        \g7[3][55] , \g7[3][54] , \g7[3][53] , \g7[3][52] , \g7[3][51] , 
        \g7[3][50] , \g7[3][49] , \g7[3][48] , \g7[3][47] , \g7[3][46] , 
        \g7[3][45] , \g7[3][44] , \g7[3][43] , \g7[3][42] , \g7[3][41] , 
        \g7[3][40] , \g7[3][39] , \g7[3][38] , \g7[3][37] , \g7[3][36] , 
        \g7[3][35] , \g7[3][34] , \g7[3][33] , \g7[3][32] , \g7[3][31] , 
        \g7[3][30] , \g7[3][29] , \g7[3][28] , \g7[3][27] , \g7[3][26] , 
        \g7[3][25] , \g7[3][24] , \g7[3][23] , \g7[3][22] , \g7[3][21] , 
        \g7[3][20] , \g7[3][19] , \g7[3][18] , \g7[3][17] , \g7[3][16] , 
        \g7[3][15] , \g7[3][14] , \g7[3][13] , \g7[3][12] , \g7[3][11] , 
        \g7[3][10] , \g7[3][9] , \g7[3][8] , \g7[3][7] , \g7[3][6] , 
        \g7[3][5] , \g7[3][4] , \g7[3][3] , \g7[3][2] , \g7[3][1] , 1'b0}), 
        .sum({\g9[0][63] , \g9[0][62] , \g9[0][61] , \g9[0][60] , \g9[0][59] , 
        \g9[0][58] , \g9[0][57] , \g9[0][56] , \g9[0][55] , \g9[0][54] , 
        \g9[0][53] , \g9[0][52] , \g9[0][51] , \g9[0][50] , \g9[0][49] , 
        \g9[0][48] , \g9[0][47] , \g9[0][46] , \g9[0][45] , \g9[0][44] , 
        \g9[0][43] , \g9[0][42] , \g9[0][41] , \g9[0][40] , \g9[0][39] , 
        \g9[0][38] , \g9[0][37] , \g9[0][36] , \g9[0][35] , \g9[0][34] , 
        \g9[0][33] , \g9[0][32] , \g9[0][31] , \g9[0][30] , \g9[0][29] , 
        \g9[0][28] , \g9[0][27] , \g9[0][26] , \g9[0][25] , \g9[0][24] , 
        \g9[0][23] , \g9[0][22] , \g9[0][21] , \g9[0][20] , \g9[0][19] , 
        \g9[0][18] , \g9[0][17] , \g9[0][16] , \g9[0][15] , \g9[0][14] , 
        \g9[0][13] , \g9[0][12] , \g9[0][11] , \g9[0][10] , \g9[0][9] , 
        \g9[0][8] , \g9[0][7] , \g9[0][6] , \g9[0][5] , \g9[0][4] , \g9[0][3] , 
        \g9[0][2] , \g9[0][1] , \g9[0][0] }), .cout({\g9[1][63] , \g9[1][62] , 
        \g9[1][61] , \g9[1][60] , \g9[1][59] , \g9[1][58] , \g9[1][57] , 
        \g9[1][56] , \g9[1][55] , \g9[1][54] , \g9[1][53] , \g9[1][52] , 
        \g9[1][51] , \g9[1][50] , \g9[1][49] , \g9[1][48] , \g9[1][47] , 
        \g9[1][46] , \g9[1][45] , \g9[1][44] , \g9[1][43] , \g9[1][42] , 
        \g9[1][41] , \g9[1][40] , \g9[1][39] , \g9[1][38] , \g9[1][37] , 
        \g9[1][36] , \g9[1][35] , \g9[1][34] , \g9[1][33] , \g9[1][32] , 
        \g9[1][31] , \g9[1][30] , \g9[1][29] , \g9[1][28] , \g9[1][27] , 
        \g9[1][26] , \g9[1][25] , \g9[1][24] , \g9[1][23] , \g9[1][22] , 
        \g9[1][21] , \g9[1][20] , \g9[1][19] , \g9[1][18] , \g9[1][17] , 
        \g9[1][16] , \g9[1][15] , \g9[1][14] , \g9[1][13] , \g9[1][12] , 
        \g9[1][11] , \g9[1][10] , \g9[1][9] , \g9[1][8] , \g9[1][7] , 
        \g9[1][6] , \g9[1][5] , \g9[1][4] , \g9[1][3] , \g9[1][2] , \g9[1][1] , 
        SYNOPSYS_UNCONNECTED__60}) );
  FullAdder F7 ( .a({\g9[0][63] , \g9[0][62] , \g9[0][61] , \g9[0][60] , 
        \g9[0][59] , \g9[0][58] , \g9[0][57] , \g9[0][56] , \g9[0][55] , 
        \g9[0][54] , \g9[0][53] , \g9[0][52] , \g9[0][51] , \g9[0][50] , 
        \g9[0][49] , \g9[0][48] , \g9[0][47] , \g9[0][46] , \g9[0][45] , 
        \g9[0][44] , \g9[0][43] , \g9[0][42] , \g9[0][41] , \g9[0][40] , 
        \g9[0][39] , \g9[0][38] , \g9[0][37] , \g9[0][36] , \g9[0][35] , 
        \g9[0][34] , \g9[0][33] , \g9[0][32] , \g9[0][31] , \g9[0][30] , 
        \g9[0][29] , \g9[0][28] , \g9[0][27] , \g9[0][26] , \g9[0][25] , 
        \g9[0][24] , \g9[0][23] , \g9[0][22] , \g9[0][21] , \g9[0][20] , 
        \g9[0][19] , \g9[0][18] , \g9[0][17] , \g9[0][16] , \g9[0][15] , 
        \g9[0][14] , \g9[0][13] , \g9[0][12] , \g9[0][11] , \g9[0][10] , 
        \g9[0][9] , \g9[0][8] , \g9[0][7] , \g9[0][6] , \g9[0][5] , \g9[0][4] , 
        \g9[0][3] , \g9[0][2] , \g9[0][1] , \g9[0][0] }), .b({\g9[1][63] , 
        \g9[1][62] , \g9[1][61] , \g9[1][60] , \g9[1][59] , \g9[1][58] , 
        \g9[1][57] , \g9[1][56] , \g9[1][55] , \g9[1][54] , \g9[1][53] , 
        \g9[1][52] , \g9[1][51] , \g9[1][50] , \g9[1][49] , \g9[1][48] , 
        \g9[1][47] , \g9[1][46] , \g9[1][45] , \g9[1][44] , \g9[1][43] , 
        \g9[1][42] , \g9[1][41] , \g9[1][40] , \g9[1][39] , \g9[1][38] , 
        \g9[1][37] , \g9[1][36] , \g9[1][35] , \g9[1][34] , \g9[1][33] , 
        \g9[1][32] , \g9[1][31] , \g9[1][30] , \g9[1][29] , \g9[1][28] , 
        \g9[1][27] , \g9[1][26] , \g9[1][25] , \g9[1][24] , \g9[1][23] , 
        \g9[1][22] , \g9[1][21] , \g9[1][20] , \g9[1][19] , \g9[1][18] , 
        \g9[1][17] , \g9[1][16] , \g9[1][15] , \g9[1][14] , \g9[1][13] , 
        \g9[1][12] , \g9[1][11] , \g9[1][10] , \g9[1][9] , \g9[1][8] , 
        \g9[1][7] , \g9[1][6] , \g9[1][5] , \g9[1][4] , \g9[1][3] , \g9[1][2] , 
        \g9[1][1] , 1'b0}), .cin({n407, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({
        \g10[0][63] , \g10[0][62] , \g10[0][61] , \g10[0][60] , \g10[0][59] , 
        \g10[0][58] , \g10[0][57] , \g10[0][56] , \g10[0][55] , \g10[0][54] , 
        \g10[0][53] , \g10[0][52] , \g10[0][51] , \g10[0][50] , \g10[0][49] , 
        \g10[0][48] , \g10[0][47] , \g10[0][46] , \g10[0][45] , \g10[0][44] , 
        \g10[0][43] , \g10[0][42] , \g10[0][41] , \g10[0][40] , \g10[0][39] , 
        \g10[0][38] , \g10[0][37] , \g10[0][36] , \g10[0][35] , \g10[0][34] , 
        \g10[0][33] , \g10[0][32] , \g10[0][31] , \g10[0][30] , \g10[0][29] , 
        \g10[0][28] , \g10[0][27] , \g10[0][26] , \g10[0][25] , \g10[0][24] , 
        \g10[0][23] , \g10[0][22] , \g10[0][21] , \g10[0][20] , \g10[0][19] , 
        \g10[0][18] , \g10[0][17] , \g10[0][16] , \g10[0][15] , \g10[0][14] , 
        \g10[0][13] , \g10[0][12] , \g10[0][11] , \g10[0][10] , \g10[0][9] , 
        \g10[0][8] , \g10[0][7] , \g10[0][6] , \g10[0][5] , \g10[0][4] , 
        \g10[0][3] , \g10[0][2] , \g10[0][1] , \g10[0][0] }), .cout({
        \g10[1][63] , \g10[1][62] , \g10[1][61] , \g10[1][60] , \g10[1][59] , 
        \g10[1][58] , \g10[1][57] , \g10[1][56] , \g10[1][55] , \g10[1][54] , 
        \g10[1][53] , \g10[1][52] , \g10[1][51] , \g10[1][50] , \g10[1][49] , 
        \g10[1][48] , \g10[1][47] , \g10[1][46] , \g10[1][45] , \g10[1][44] , 
        \g10[1][43] , \g10[1][42] , \g10[1][41] , \g10[1][40] , \g10[1][39] , 
        \g10[1][38] , \g10[1][37] , \g10[1][36] , \g10[1][35] , \g10[1][34] , 
        \g10[1][33] , \g10[1][32] , \g10[1][31] , \g10[1][30] , \g10[1][29] , 
        \g10[1][28] , \g10[1][27] , \g10[1][26] , \g10[1][25] , \g10[1][24] , 
        \g10[1][23] , \g10[1][22] , \g10[1][21] , \g10[1][20] , \g10[1][19] , 
        \g10[1][18] , \g10[1][17] , \g10[1][16] , \g10[1][15] , \g10[1][14] , 
        \g10[1][13] , \g10[1][12] , \g10[1][11] , \g10[1][10] , \g10[1][9] , 
        \g10[1][8] , \g10[1][7] , \g10[1][6] , \g10[1][5] , \g10[1][4] , 
        \g10[1][3] , \g10[1][2] , \g10[1][1] , SYNOPSYS_UNCONNECTED__61}) );
  WallaceTreeMultiplier_DW01_add_0 add_110 ( .A({\g10[1][63] , \g10[1][62] , 
        \g10[1][61] , \g10[1][60] , \g10[1][59] , \g10[1][58] , \g10[1][57] , 
        \g10[1][56] , \g10[1][55] , \g10[1][54] , \g10[1][53] , \g10[1][52] , 
        \g10[1][51] , \g10[1][50] , \g10[1][49] , \g10[1][48] , \g10[1][47] , 
        \g10[1][46] , \g10[1][45] , \g10[1][44] , \g10[1][43] , \g10[1][42] , 
        \g10[1][41] , \g10[1][40] , \g10[1][39] , \g10[1][38] , \g10[1][37] , 
        \g10[1][36] , \g10[1][35] , \g10[1][34] , \g10[1][33] , \g10[1][32] , 
        \g10[1][31] , \g10[1][30] , \g10[1][29] , \g10[1][28] , \g10[1][27] , 
        \g10[1][26] , \g10[1][25] , \g10[1][24] , \g10[1][23] , \g10[1][22] , 
        \g10[1][21] , \g10[1][20] , \g10[1][19] , \g10[1][18] , \g10[1][17] , 
        \g10[1][16] , \g10[1][15] , \g10[1][14] , \g10[1][13] , \g10[1][12] , 
        \g10[1][11] , \g10[1][10] , \g10[1][9] , \g10[1][8] , \g10[1][7] , 
        \g10[1][6] , \g10[1][5] , \g10[1][4] , \g10[1][3] , \g10[1][2] , 
        \g10[1][1] , 1'b0}), .B({\g10[0][63] , \g10[0][62] , \g10[0][61] , 
        \g10[0][60] , \g10[0][59] , \g10[0][58] , \g10[0][57] , \g10[0][56] , 
        \g10[0][55] , \g10[0][54] , \g10[0][53] , \g10[0][52] , \g10[0][51] , 
        \g10[0][50] , \g10[0][49] , \g10[0][48] , \g10[0][47] , \g10[0][46] , 
        \g10[0][45] , \g10[0][44] , \g10[0][43] , \g10[0][42] , \g10[0][41] , 
        \g10[0][40] , \g10[0][39] , \g10[0][38] , \g10[0][37] , \g10[0][36] , 
        \g10[0][35] , \g10[0][34] , \g10[0][33] , \g10[0][32] , \g10[0][31] , 
        \g10[0][30] , \g10[0][29] , \g10[0][28] , \g10[0][27] , \g10[0][26] , 
        \g10[0][25] , \g10[0][24] , \g10[0][23] , \g10[0][22] , \g10[0][21] , 
        \g10[0][20] , \g10[0][19] , \g10[0][18] , \g10[0][17] , \g10[0][16] , 
        \g10[0][15] , \g10[0][14] , \g10[0][13] , \g10[0][12] , \g10[0][11] , 
        \g10[0][10] , \g10[0][9] , \g10[0][8] , \g10[0][7] , \g10[0][6] , 
        \g10[0][5] , \g10[0][4] , \g10[0][3] , \g10[0][2] , \g10[0][1] , 
        \g10[0][0] }), .CI(1'b0), .SUM({N194, N193, N192, N191, N190, N189, 
        N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, 
        N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, 
        N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, 
        N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, 
        N140, N139, N138, N137, N136, N135, N134, N133, N132, N131}) );
  DFF_X1 \out_reg[63]  ( .D(N258), .CK(clk), .Q(out[63]) );
  BUF_X2 U1219 ( .A(n132), .Z(n316) );
  BUF_X2 U1220 ( .A(n66), .Z(n214) );
  AND2_X1 U1221 ( .A1(N132), .A2(n142), .ZN(N196) );
  BUF_X1 U1222 ( .A(n125), .Z(n127) );
  INV_X1 U1223 ( .A(A_reg[1]), .ZN(n442) );
  CLKBUF_X1 U1224 ( .A(A_reg[3]), .Z(n109) );
  AND2_X1 U1225 ( .A1(A_reg[6]), .A2(B_reg[0]), .ZN(\p[0][6] ) );
  BUF_X2 U1226 ( .A(n132), .Z(n317) );
  INV_X2 U1227 ( .A(A_reg[2]), .ZN(n441) );
  INV_X1 U1228 ( .A(B_reg[1]), .ZN(n110) );
  AND2_X1 U1229 ( .A1(B_reg[0]), .A2(A_reg[7]), .ZN(\p[0][7] ) );
  BUF_X1 U1230 ( .A(A_reg[5]), .Z(n111) );
  BUF_X2 U1231 ( .A(n66), .Z(n215) );
  BUF_X2 U1232 ( .A(n440), .Z(n226) );
  AND2_X1 U1233 ( .A1(A_reg[3]), .A2(B_reg[3]), .ZN(\p[3][6] ) );
  AND2_X1 U1234 ( .A1(B_reg[3]), .A2(A_reg[5]), .ZN(\p[3][8] ) );
  BUF_X2 U1235 ( .A(n115), .Z(n302) );
  BUF_X2 U1236 ( .A(n133), .Z(n136) );
  BUF_X1 U1237 ( .A(n130), .Z(n113) );
  INV_X1 U1238 ( .A(n132), .ZN(n114) );
  CLKBUF_X1 U1239 ( .A(n67), .Z(n217) );
  BUF_X1 U1240 ( .A(n67), .Z(n218) );
  BUF_X1 U1241 ( .A(n115), .Z(n301) );
  CLKBUF_X1 U1242 ( .A(n122), .Z(n308) );
  BUF_X2 U1243 ( .A(n441), .Z(n232) );
  CLKBUF_X1 U1244 ( .A(n90), .Z(n207) );
  CLKBUF_X1 U1245 ( .A(n66), .Z(n213) );
  CLKBUF_X1 U1246 ( .A(n91), .Z(n210) );
  CLKBUF_X1 U1247 ( .A(n112), .Z(n299) );
  BUF_X2 U1248 ( .A(n68), .Z(n303) );
  CLKBUF_X1 U1249 ( .A(n118), .Z(n313) );
  CLKBUF_X1 U1250 ( .A(n68), .Z(n304) );
  CLKBUF_X1 U1251 ( .A(n92), .Z(n296) );
  CLKBUF_X1 U1252 ( .A(n93), .Z(n293) );
  BUF_X1 U1253 ( .A(n444), .Z(n311) );
  CLKBUF_X1 U1254 ( .A(n440), .Z(n227) );
  BUF_X1 U1255 ( .A(n442), .Z(n234) );
  CLKBUF_X1 U1256 ( .A(n68), .Z(n305) );
  CLKBUF_X1 U1257 ( .A(n112), .Z(n298) );
  CLKBUF_X1 U1258 ( .A(n92), .Z(n295) );
  CLKBUF_X1 U1259 ( .A(n93), .Z(n292) );
  BUF_X1 U1260 ( .A(\p[54][63] ), .Z(n379) );
  BUF_X1 U1261 ( .A(\p[53][63] ), .Z(n377) );
  BUF_X1 U1262 ( .A(\p[52][63] ), .Z(n375) );
  BUF_X1 U1263 ( .A(\p[9][63] ), .Z(n323) );
  BUF_X1 U1264 ( .A(\p[10][63] ), .Z(n325) );
  BUF_X1 U1265 ( .A(\p[11][63] ), .Z(n327) );
  BUF_X1 U1266 ( .A(n139), .Z(n222) );
  BUF_X1 U1267 ( .A(n140), .Z(n229) );
  NOR2_X1 U1268 ( .A1(n439), .A2(n125), .ZN(\p[6][13] ) );
  NOR2_X1 U1269 ( .A1(n227), .A2(n125), .ZN(\p[6][10] ) );
  AND2_X1 U1270 ( .A1(n433), .A2(A_reg[21]), .ZN(\p[42][63] ) );
  AND2_X1 U1271 ( .A1(B_reg[21]), .A2(n436), .ZN(\p[21][63] ) );
  AND2_X1 U1272 ( .A1(B_reg[22]), .A2(n436), .ZN(\p[22][63] ) );
  AND2_X1 U1273 ( .A1(n433), .A2(A_reg[22]), .ZN(\p[41][63] ) );
  AND2_X1 U1274 ( .A1(n433), .A2(A_reg[23]), .ZN(\p[40][63] ) );
  AND2_X1 U1275 ( .A1(B_reg[23]), .A2(n436), .ZN(\p[23][63] ) );
  NOR2_X1 U1276 ( .A1(n232), .A2(n294), .ZN(\p[12][14] ) );
  NOR2_X1 U1277 ( .A1(n232), .A2(n276), .ZN(\p[18][20] ) );
  NOR2_X1 U1278 ( .A1(n192), .A2(n306), .ZN(\p[7][24] ) );
  NOR2_X1 U1279 ( .A1(n186), .A2(n306), .ZN(\p[7][26] ) );
  NOR2_X1 U1280 ( .A1(n220), .A2(n305), .ZN(\p[8][15] ) );
  NOR2_X1 U1281 ( .A1(n220), .A2(n296), .ZN(\p[11][18] ) );
  NOR2_X1 U1282 ( .A1(n220), .A2(n287), .ZN(\p[14][21] ) );
  NOR2_X1 U1283 ( .A1(n220), .A2(n278), .ZN(\p[17][24] ) );
  NOR2_X1 U1284 ( .A1(n220), .A2(n293), .ZN(\p[12][19] ) );
  NOR2_X1 U1285 ( .A1(n220), .A2(n284), .ZN(\p[15][22] ) );
  NOR2_X1 U1286 ( .A1(n220), .A2(n275), .ZN(\p[18][25] ) );
  NOR2_X1 U1287 ( .A1(n219), .A2(n305), .ZN(\p[8][16] ) );
  NOR2_X1 U1288 ( .A1(n219), .A2(n278), .ZN(\p[17][25] ) );
  NOR2_X1 U1289 ( .A1(n219), .A2(n275), .ZN(\p[18][26] ) );
  NOR2_X1 U1290 ( .A1(n220), .A2(n299), .ZN(\p[10][17] ) );
  NOR2_X1 U1291 ( .A1(n220), .A2(n290), .ZN(\p[13][20] ) );
  NOR2_X1 U1292 ( .A1(n220), .A2(n281), .ZN(\p[16][23] ) );
  NOR2_X1 U1293 ( .A1(n220), .A2(n272), .ZN(\p[19][26] ) );
  NOR2_X1 U1294 ( .A1(n226), .A2(n297), .ZN(\p[11][15] ) );
  NOR2_X1 U1295 ( .A1(n226), .A2(n294), .ZN(\p[12][16] ) );
  NOR2_X1 U1296 ( .A1(n219), .A2(n307), .ZN(\p[7][15] ) );
  NOR2_X1 U1297 ( .A1(n219), .A2(n281), .ZN(\p[16][24] ) );
  NOR2_X1 U1298 ( .A1(n215), .A2(n296), .ZN(\p[11][21] ) );
  NOR2_X1 U1299 ( .A1(n212), .A2(n296), .ZN(\p[11][22] ) );
  NOR2_X1 U1300 ( .A1(n209), .A2(n296), .ZN(\p[11][23] ) );
  NOR2_X1 U1301 ( .A1(n206), .A2(n296), .ZN(\p[11][24] ) );
  NOR2_X1 U1302 ( .A1(n215), .A2(n287), .ZN(\p[14][24] ) );
  NOR2_X1 U1303 ( .A1(n203), .A2(n296), .ZN(\p[11][25] ) );
  NOR2_X1 U1304 ( .A1(n212), .A2(n287), .ZN(\p[14][25] ) );
  NOR2_X1 U1305 ( .A1(n200), .A2(n296), .ZN(\p[11][26] ) );
  NOR2_X1 U1306 ( .A1(n209), .A2(n287), .ZN(\p[14][26] ) );
  NOR2_X1 U1307 ( .A1(n215), .A2(n293), .ZN(\p[12][22] ) );
  NOR2_X1 U1308 ( .A1(n212), .A2(n293), .ZN(\p[12][23] ) );
  NOR2_X1 U1309 ( .A1(n209), .A2(n293), .ZN(\p[12][24] ) );
  NOR2_X1 U1310 ( .A1(n206), .A2(n293), .ZN(\p[12][25] ) );
  NOR2_X1 U1311 ( .A1(n215), .A2(n284), .ZN(\p[15][25] ) );
  NOR2_X1 U1312 ( .A1(n203), .A2(n293), .ZN(\p[12][26] ) );
  NOR2_X1 U1313 ( .A1(n212), .A2(n284), .ZN(\p[15][26] ) );
  NOR2_X1 U1314 ( .A1(n200), .A2(n293), .ZN(\p[12][27] ) );
  NOR2_X1 U1315 ( .A1(n215), .A2(n299), .ZN(\p[10][20] ) );
  NOR2_X1 U1316 ( .A1(n212), .A2(n299), .ZN(\p[10][21] ) );
  NOR2_X1 U1317 ( .A1(n209), .A2(n299), .ZN(\p[10][22] ) );
  NOR2_X1 U1318 ( .A1(n206), .A2(n299), .ZN(\p[10][23] ) );
  NOR2_X1 U1319 ( .A1(n215), .A2(n290), .ZN(\p[13][23] ) );
  NOR2_X1 U1320 ( .A1(n203), .A2(n299), .ZN(\p[10][24] ) );
  NOR2_X1 U1321 ( .A1(n212), .A2(n290), .ZN(\p[13][24] ) );
  NOR2_X1 U1322 ( .A1(n200), .A2(n299), .ZN(\p[10][25] ) );
  NOR2_X1 U1323 ( .A1(n209), .A2(n290), .ZN(\p[13][25] ) );
  NOR2_X1 U1324 ( .A1(n197), .A2(n299), .ZN(\p[10][26] ) );
  NOR2_X1 U1325 ( .A1(n206), .A2(n290), .ZN(\p[13][26] ) );
  NOR2_X1 U1326 ( .A1(n194), .A2(n299), .ZN(\p[10][27] ) );
  NOR2_X1 U1327 ( .A1(n203), .A2(n290), .ZN(\p[13][27] ) );
  NOR2_X1 U1328 ( .A1(n227), .A2(n288), .ZN(\p[14][18] ) );
  NOR2_X1 U1329 ( .A1(n226), .A2(n279), .ZN(\p[17][21] ) );
  NOR2_X1 U1330 ( .A1(n226), .A2(n270), .ZN(\p[20][24] ) );
  NOR2_X1 U1331 ( .A1(n236), .A2(n279), .ZN(\p[17][17] ) );
  NOR2_X1 U1332 ( .A1(n236), .A2(n270), .ZN(\p[20][20] ) );
  NOR2_X1 U1333 ( .A1(n236), .A2(n261), .ZN(\p[23][23] ) );
  NOR2_X1 U1334 ( .A1(n226), .A2(n285), .ZN(\p[15][19] ) );
  NOR2_X1 U1335 ( .A1(n226), .A2(n276), .ZN(\p[18][22] ) );
  NOR2_X1 U1336 ( .A1(n227), .A2(n267), .ZN(\p[21][25] ) );
  NOR2_X1 U1337 ( .A1(n236), .A2(n285), .ZN(\p[15][15] ) );
  NOR2_X1 U1338 ( .A1(n236), .A2(n276), .ZN(\p[18][18] ) );
  NOR2_X1 U1339 ( .A1(n236), .A2(n267), .ZN(\p[21][21] ) );
  NOR2_X1 U1340 ( .A1(n236), .A2(n258), .ZN(\p[24][24] ) );
  NOR2_X1 U1341 ( .A1(n236), .A2(n249), .ZN(\p[27][27] ) );
  NOR2_X1 U1342 ( .A1(n302), .A2(n220), .ZN(\p[9][16] ) );
  NOR2_X1 U1343 ( .A1(n226), .A2(n305), .ZN(\p[8][12] ) );
  NOR2_X1 U1344 ( .A1(n232), .A2(n261), .ZN(\p[23][25] ) );
  NOR2_X1 U1345 ( .A1(n301), .A2(n219), .ZN(\p[9][17] ) );
  NOR2_X1 U1346 ( .A1(n226), .A2(n291), .ZN(\p[13][17] ) );
  NOR2_X1 U1347 ( .A1(n227), .A2(n282), .ZN(\p[16][20] ) );
  NOR2_X1 U1348 ( .A1(n227), .A2(n273), .ZN(\p[19][23] ) );
  NOR2_X1 U1349 ( .A1(n227), .A2(n264), .ZN(\p[22][26] ) );
  NOR2_X1 U1350 ( .A1(n236), .A2(n315), .ZN(\p[1][1] ) );
  NOR2_X1 U1351 ( .A1(n236), .A2(n282), .ZN(\p[16][16] ) );
  NOR2_X1 U1352 ( .A1(n236), .A2(n273), .ZN(\p[19][19] ) );
  NOR2_X1 U1353 ( .A1(n236), .A2(n264), .ZN(\p[22][22] ) );
  NOR2_X1 U1354 ( .A1(n236), .A2(n255), .ZN(\p[25][25] ) );
  NOR2_X1 U1355 ( .A1(n232), .A2(n267), .ZN(\p[21][23] ) );
  NOR2_X1 U1356 ( .A1(n207), .A2(n314), .ZN(\p[2][14] ) );
  NOR2_X1 U1357 ( .A1(n204), .A2(n314), .ZN(\p[2][15] ) );
  NOR2_X1 U1358 ( .A1(n201), .A2(n314), .ZN(\p[2][16] ) );
  NOR2_X1 U1359 ( .A1(n213), .A2(n314), .ZN(\p[2][12] ) );
  NOR2_X1 U1360 ( .A1(n217), .A2(n314), .ZN(\p[2][11] ) );
  NOR2_X1 U1361 ( .A1(n210), .A2(n314), .ZN(\p[2][13] ) );
  NOR2_X1 U1362 ( .A1(n225), .A2(n297), .ZN(\p[11][16] ) );
  NOR2_X1 U1363 ( .A1(n225), .A2(n288), .ZN(\p[14][19] ) );
  NOR2_X1 U1364 ( .A1(n225), .A2(n294), .ZN(\p[12][17] ) );
  NOR2_X1 U1365 ( .A1(n234), .A2(n288), .ZN(\p[14][15] ) );
  NOR2_X1 U1366 ( .A1(n234), .A2(n279), .ZN(\p[17][18] ) );
  NOR2_X1 U1367 ( .A1(n234), .A2(n270), .ZN(\p[20][21] ) );
  NOR2_X1 U1368 ( .A1(n234), .A2(n261), .ZN(\p[23][24] ) );
  NOR2_X1 U1369 ( .A1(n225), .A2(n285), .ZN(\p[15][20] ) );
  NOR2_X1 U1370 ( .A1(n234), .A2(n285), .ZN(\p[15][16] ) );
  NOR2_X1 U1371 ( .A1(n234), .A2(n276), .ZN(\p[18][19] ) );
  NOR2_X1 U1372 ( .A1(n234), .A2(n267), .ZN(\p[21][22] ) );
  NOR2_X1 U1373 ( .A1(n234), .A2(n258), .ZN(\p[24][25] ) );
  NOR2_X1 U1374 ( .A1(n235), .A2(n288), .ZN(\p[14][14] ) );
  NOR2_X1 U1375 ( .A1(n216), .A2(n309), .ZN(\p[5][14] ) );
  NOR2_X1 U1376 ( .A1(n213), .A2(n309), .ZN(\p[5][15] ) );
  NOR2_X1 U1377 ( .A1(n210), .A2(n309), .ZN(\p[5][16] ) );
  NOR2_X1 U1378 ( .A1(n226), .A2(n112), .ZN(\p[10][14] ) );
  NOR2_X1 U1379 ( .A1(n207), .A2(n308), .ZN(\p[5][17] ) );
  NOR2_X1 U1380 ( .A1(n204), .A2(n308), .ZN(\p[5][18] ) );
  NOR2_X1 U1381 ( .A1(n201), .A2(n308), .ZN(\p[5][19] ) );
  NOR2_X1 U1382 ( .A1(n198), .A2(n308), .ZN(\p[5][20] ) );
  NOR2_X1 U1383 ( .A1(n195), .A2(n308), .ZN(\p[5][21] ) );
  NOR2_X1 U1384 ( .A1(n192), .A2(n308), .ZN(\p[5][22] ) );
  NOR2_X1 U1385 ( .A1(n189), .A2(n308), .ZN(\p[5][23] ) );
  NOR2_X1 U1386 ( .A1(n186), .A2(n308), .ZN(\p[5][24] ) );
  NOR2_X1 U1387 ( .A1(n183), .A2(n308), .ZN(\p[5][25] ) );
  NOR2_X1 U1388 ( .A1(n180), .A2(n308), .ZN(\p[5][26] ) );
  NOR2_X1 U1389 ( .A1(n196), .A2(n315), .ZN(\p[1][17] ) );
  NOR2_X1 U1390 ( .A1(n211), .A2(n315), .ZN(\p[1][12] ) );
  NOR2_X1 U1391 ( .A1(n199), .A2(n315), .ZN(\p[1][16] ) );
  NOR2_X1 U1392 ( .A1(n208), .A2(n315), .ZN(\p[1][13] ) );
  NOR2_X1 U1393 ( .A1(n205), .A2(n315), .ZN(\p[1][14] ) );
  NOR2_X1 U1394 ( .A1(n202), .A2(n315), .ZN(\p[1][15] ) );
  NOR2_X1 U1395 ( .A1(n193), .A2(n315), .ZN(\p[1][18] ) );
  NOR2_X1 U1396 ( .A1(n190), .A2(n315), .ZN(\p[1][19] ) );
  NOR2_X1 U1397 ( .A1(n187), .A2(n315), .ZN(\p[1][20] ) );
  NOR2_X1 U1398 ( .A1(n184), .A2(n315), .ZN(\p[1][21] ) );
  NOR2_X1 U1399 ( .A1(n181), .A2(n315), .ZN(\p[1][22] ) );
  NOR2_X1 U1400 ( .A1(n178), .A2(n315), .ZN(\p[1][23] ) );
  NOR2_X1 U1401 ( .A1(n175), .A2(n315), .ZN(\p[1][24] ) );
  NOR2_X1 U1402 ( .A1(n172), .A2(n315), .ZN(\p[1][25] ) );
  NOR2_X1 U1403 ( .A1(n169), .A2(n315), .ZN(\p[1][26] ) );
  NOR2_X1 U1404 ( .A1(n166), .A2(n315), .ZN(\p[1][27] ) );
  NOR2_X1 U1405 ( .A1(n225), .A2(n300), .ZN(\p[10][15] ) );
  NOR2_X1 U1406 ( .A1(n225), .A2(n291), .ZN(\p[13][18] ) );
  NOR2_X1 U1407 ( .A1(n234), .A2(n282), .ZN(\p[16][17] ) );
  NOR2_X1 U1408 ( .A1(n234), .A2(n273), .ZN(\p[19][20] ) );
  NOR2_X1 U1409 ( .A1(n234), .A2(n264), .ZN(\p[22][23] ) );
  NOR2_X1 U1410 ( .A1(n198), .A2(n313), .ZN(\p[2][17] ) );
  NOR2_X1 U1411 ( .A1(n216), .A2(n304), .ZN(\p[8][17] ) );
  NOR2_X1 U1412 ( .A1(n195), .A2(n313), .ZN(\p[2][18] ) );
  NOR2_X1 U1413 ( .A1(n213), .A2(n304), .ZN(\p[8][18] ) );
  NOR2_X1 U1414 ( .A1(n192), .A2(n313), .ZN(\p[2][19] ) );
  NOR2_X1 U1415 ( .A1(n210), .A2(n304), .ZN(\p[8][19] ) );
  NOR2_X1 U1416 ( .A1(n189), .A2(n313), .ZN(\p[2][20] ) );
  NOR2_X1 U1417 ( .A1(n207), .A2(n304), .ZN(\p[8][20] ) );
  NOR2_X1 U1418 ( .A1(n186), .A2(n313), .ZN(\p[2][21] ) );
  NOR2_X1 U1419 ( .A1(n204), .A2(n304), .ZN(\p[8][21] ) );
  NOR2_X1 U1420 ( .A1(n183), .A2(n313), .ZN(\p[2][22] ) );
  NOR2_X1 U1421 ( .A1(n201), .A2(n304), .ZN(\p[8][22] ) );
  NOR2_X1 U1422 ( .A1(n180), .A2(n313), .ZN(\p[2][23] ) );
  NOR2_X1 U1423 ( .A1(n198), .A2(n304), .ZN(\p[8][23] ) );
  NOR2_X1 U1424 ( .A1(n195), .A2(n304), .ZN(\p[8][24] ) );
  NOR2_X1 U1425 ( .A1(n192), .A2(n304), .ZN(\p[8][25] ) );
  NOR2_X1 U1426 ( .A1(n177), .A2(n313), .ZN(\p[2][24] ) );
  NOR2_X1 U1427 ( .A1(n174), .A2(n313), .ZN(\p[2][25] ) );
  NOR2_X1 U1428 ( .A1(n204), .A2(n311), .ZN(\p[4][17] ) );
  NOR2_X1 U1429 ( .A1(n207), .A2(n311), .ZN(\p[4][16] ) );
  NOR2_X1 U1430 ( .A1(n210), .A2(n311), .ZN(\p[4][15] ) );
  NOR2_X1 U1431 ( .A1(n201), .A2(n311), .ZN(\p[4][18] ) );
  NOR2_X1 U1432 ( .A1(n198), .A2(n311), .ZN(\p[4][19] ) );
  NOR2_X1 U1433 ( .A1(n195), .A2(n311), .ZN(\p[4][20] ) );
  NOR2_X1 U1434 ( .A1(n192), .A2(n311), .ZN(\p[4][21] ) );
  NOR2_X1 U1435 ( .A1(n189), .A2(n311), .ZN(\p[4][22] ) );
  NOR2_X1 U1436 ( .A1(n186), .A2(n311), .ZN(\p[4][23] ) );
  NOR2_X1 U1437 ( .A1(n183), .A2(n311), .ZN(\p[4][24] ) );
  NOR2_X1 U1438 ( .A1(n180), .A2(n311), .ZN(\p[4][25] ) );
  NOR2_X1 U1439 ( .A1(n177), .A2(n311), .ZN(\p[4][26] ) );
  NOR2_X1 U1440 ( .A1(n174), .A2(n311), .ZN(\p[4][27] ) );
  NOR2_X1 U1441 ( .A1(n216), .A2(n307), .ZN(\p[7][16] ) );
  NOR2_X1 U1442 ( .A1(n221), .A2(n307), .ZN(\p[7][14] ) );
  NOR2_X1 U1443 ( .A1(n213), .A2(n307), .ZN(\p[7][17] ) );
  NOR2_X1 U1444 ( .A1(n210), .A2(n307), .ZN(\p[7][18] ) );
  NOR2_X1 U1445 ( .A1(n207), .A2(n307), .ZN(\p[7][19] ) );
  NOR2_X1 U1446 ( .A1(n204), .A2(n307), .ZN(\p[7][20] ) );
  NOR2_X1 U1447 ( .A1(n201), .A2(n307), .ZN(\p[7][21] ) );
  NOR2_X1 U1448 ( .A1(n198), .A2(n307), .ZN(\p[7][22] ) );
  NOR2_X1 U1449 ( .A1(n195), .A2(n307), .ZN(\p[7][23] ) );
  NOR2_X1 U1450 ( .A1(n189), .A2(n307), .ZN(\p[7][25] ) );
  NOR2_X1 U1451 ( .A1(n171), .A2(n313), .ZN(\p[2][26] ) );
  NOR2_X1 U1452 ( .A1(n301), .A2(n216), .ZN(\p[9][18] ) );
  NOR2_X1 U1453 ( .A1(n301), .A2(n213), .ZN(\p[9][19] ) );
  NOR2_X1 U1454 ( .A1(n301), .A2(n210), .ZN(\p[9][20] ) );
  NOR2_X1 U1455 ( .A1(n301), .A2(n207), .ZN(\p[9][21] ) );
  NOR2_X1 U1456 ( .A1(n301), .A2(n204), .ZN(\p[9][22] ) );
  NOR2_X1 U1457 ( .A1(n301), .A2(n201), .ZN(\p[9][23] ) );
  NOR2_X1 U1458 ( .A1(n301), .A2(n198), .ZN(\p[9][24] ) );
  NOR2_X1 U1459 ( .A1(n301), .A2(n195), .ZN(\p[9][25] ) );
  NOR2_X1 U1460 ( .A1(n301), .A2(n192), .ZN(\p[9][26] ) );
  NOR2_X1 U1461 ( .A1(n301), .A2(n189), .ZN(\p[9][27] ) );
  NOR2_X1 U1462 ( .A1(n216), .A2(n281), .ZN(\p[16][25] ) );
  NOR2_X1 U1463 ( .A1(n214), .A2(n281), .ZN(\p[16][26] ) );
  BUF_X1 U1464 ( .A(\p[62][63] ), .Z(n404) );
  BUF_X2 U1465 ( .A(\p[63][63] ), .Z(n405) );
  BUF_X2 U1466 ( .A(\p[62][63] ), .Z(n402) );
  BUF_X2 U1467 ( .A(\p[60][63] ), .Z(n396) );
  BUF_X2 U1468 ( .A(\p[58][63] ), .Z(n390) );
  BUF_X2 U1469 ( .A(\p[59][63] ), .Z(n393) );
  BUF_X2 U1470 ( .A(\p[57][63] ), .Z(n387) );
  BUF_X2 U1471 ( .A(\p[56][63] ), .Z(n384) );
  BUF_X2 U1472 ( .A(\p[0][63] ), .Z(n408) );
  BUF_X2 U1473 ( .A(\p[3][63] ), .Z(n417) );
  BUF_X2 U1474 ( .A(\p[6][63] ), .Z(n426) );
  BUF_X2 U1475 ( .A(\p[63][63] ), .Z(n406) );
  BUF_X2 U1476 ( .A(\p[62][63] ), .Z(n403) );
  BUF_X2 U1477 ( .A(\p[60][63] ), .Z(n397) );
  BUF_X2 U1478 ( .A(\p[58][63] ), .Z(n391) );
  BUF_X2 U1479 ( .A(\p[59][63] ), .Z(n394) );
  BUF_X2 U1480 ( .A(\p[57][63] ), .Z(n388) );
  BUF_X2 U1481 ( .A(\p[56][63] ), .Z(n385) );
  BUF_X2 U1482 ( .A(\p[4][63] ), .Z(n420) );
  BUF_X2 U1483 ( .A(\p[1][63] ), .Z(n411) );
  BUF_X1 U1484 ( .A(\p[60][63] ), .Z(n398) );
  BUF_X1 U1485 ( .A(\p[63][63] ), .Z(n407) );
  BUF_X1 U1486 ( .A(\p[59][63] ), .Z(n395) );
  BUF_X1 U1487 ( .A(\p[58][63] ), .Z(n392) );
  NOR2_X1 U1488 ( .A1(n180), .A2(n306), .ZN(\p[7][28] ) );
  NOR2_X1 U1489 ( .A1(n220), .A2(n269), .ZN(\p[20][27] ) );
  NOR2_X1 U1490 ( .A1(n220), .A2(n260), .ZN(\p[23][30] ) );
  NOR2_X1 U1491 ( .A1(n220), .A2(n251), .ZN(\p[26][33] ) );
  NOR2_X1 U1492 ( .A1(n220), .A2(n242), .ZN(\p[29][36] ) );
  NOR2_X1 U1493 ( .A1(n220), .A2(n266), .ZN(\p[21][28] ) );
  NOR2_X1 U1494 ( .A1(n220), .A2(n257), .ZN(\p[24][31] ) );
  NOR2_X1 U1495 ( .A1(n220), .A2(n248), .ZN(\p[27][34] ) );
  NOR2_X1 U1496 ( .A1(n220), .A2(n239), .ZN(\p[30][37] ) );
  NOR2_X1 U1497 ( .A1(n219), .A2(n269), .ZN(\p[20][28] ) );
  NOR2_X1 U1498 ( .A1(n219), .A2(n260), .ZN(\p[23][31] ) );
  NOR2_X1 U1499 ( .A1(n219), .A2(n251), .ZN(\p[26][34] ) );
  NOR2_X1 U1500 ( .A1(n219), .A2(n242), .ZN(\p[29][37] ) );
  NOR2_X1 U1501 ( .A1(n219), .A2(n266), .ZN(\p[21][29] ) );
  NOR2_X1 U1502 ( .A1(n219), .A2(n257), .ZN(\p[24][32] ) );
  NOR2_X1 U1503 ( .A1(n219), .A2(n248), .ZN(\p[27][35] ) );
  NOR2_X1 U1504 ( .A1(n219), .A2(n239), .ZN(\p[30][38] ) );
  NOR2_X1 U1505 ( .A1(n220), .A2(n263), .ZN(\p[22][29] ) );
  NOR2_X1 U1506 ( .A1(n220), .A2(n254), .ZN(\p[25][32] ) );
  NOR2_X1 U1507 ( .A1(n220), .A2(n245), .ZN(\p[28][35] ) );
  NOR2_X1 U1508 ( .A1(n219), .A2(n272), .ZN(\p[19][27] ) );
  NOR2_X1 U1509 ( .A1(n219), .A2(n263), .ZN(\p[22][30] ) );
  NOR2_X1 U1510 ( .A1(n219), .A2(n254), .ZN(\p[25][33] ) );
  NOR2_X1 U1511 ( .A1(n219), .A2(n245), .ZN(\p[28][36] ) );
  NOR2_X1 U1512 ( .A1(n197), .A2(n296), .ZN(\p[11][27] ) );
  NOR2_X1 U1513 ( .A1(n206), .A2(n287), .ZN(\p[14][27] ) );
  NOR2_X1 U1514 ( .A1(n194), .A2(n296), .ZN(\p[11][28] ) );
  NOR2_X1 U1515 ( .A1(n203), .A2(n287), .ZN(\p[14][28] ) );
  NOR2_X1 U1516 ( .A1(n191), .A2(n296), .ZN(\p[11][29] ) );
  NOR2_X1 U1517 ( .A1(n200), .A2(n287), .ZN(\p[14][29] ) );
  NOR2_X1 U1518 ( .A1(n188), .A2(n295), .ZN(\p[11][30] ) );
  NOR2_X1 U1519 ( .A1(n197), .A2(n287), .ZN(\p[14][30] ) );
  NOR2_X1 U1520 ( .A1(n185), .A2(n295), .ZN(\p[11][31] ) );
  NOR2_X1 U1521 ( .A1(n194), .A2(n287), .ZN(\p[14][31] ) );
  NOR2_X1 U1522 ( .A1(n182), .A2(n295), .ZN(\p[11][32] ) );
  NOR2_X1 U1523 ( .A1(n191), .A2(n287), .ZN(\p[14][32] ) );
  NOR2_X1 U1524 ( .A1(n188), .A2(n286), .ZN(\p[14][33] ) );
  NOR2_X1 U1525 ( .A1(n179), .A2(n295), .ZN(\p[11][33] ) );
  NOR2_X1 U1526 ( .A1(n185), .A2(n286), .ZN(\p[14][34] ) );
  NOR2_X1 U1527 ( .A1(n176), .A2(n295), .ZN(\p[11][34] ) );
  NOR2_X1 U1528 ( .A1(n182), .A2(n286), .ZN(\p[14][35] ) );
  NOR2_X1 U1529 ( .A1(n173), .A2(n295), .ZN(\p[11][35] ) );
  NOR2_X1 U1530 ( .A1(n179), .A2(n286), .ZN(\p[14][36] ) );
  NOR2_X1 U1531 ( .A1(n170), .A2(n295), .ZN(\p[11][36] ) );
  NOR2_X1 U1532 ( .A1(n176), .A2(n286), .ZN(\p[14][37] ) );
  NOR2_X1 U1533 ( .A1(n167), .A2(n295), .ZN(\p[11][37] ) );
  NOR2_X1 U1534 ( .A1(n173), .A2(n286), .ZN(\p[14][38] ) );
  NOR2_X1 U1535 ( .A1(n209), .A2(n284), .ZN(\p[15][27] ) );
  NOR2_X1 U1536 ( .A1(n197), .A2(n293), .ZN(\p[12][28] ) );
  NOR2_X1 U1537 ( .A1(n206), .A2(n284), .ZN(\p[15][28] ) );
  NOR2_X1 U1538 ( .A1(n194), .A2(n293), .ZN(\p[12][29] ) );
  NOR2_X1 U1539 ( .A1(n203), .A2(n284), .ZN(\p[15][29] ) );
  NOR2_X1 U1540 ( .A1(n191), .A2(n293), .ZN(\p[12][30] ) );
  NOR2_X1 U1541 ( .A1(n200), .A2(n284), .ZN(\p[15][30] ) );
  NOR2_X1 U1542 ( .A1(n188), .A2(n292), .ZN(\p[12][31] ) );
  NOR2_X1 U1543 ( .A1(n197), .A2(n284), .ZN(\p[15][31] ) );
  NOR2_X1 U1544 ( .A1(n185), .A2(n292), .ZN(\p[12][32] ) );
  NOR2_X1 U1545 ( .A1(n194), .A2(n284), .ZN(\p[15][32] ) );
  NOR2_X1 U1546 ( .A1(n182), .A2(n292), .ZN(\p[12][33] ) );
  NOR2_X1 U1547 ( .A1(n191), .A2(n284), .ZN(\p[15][33] ) );
  NOR2_X1 U1548 ( .A1(n179), .A2(n292), .ZN(\p[12][34] ) );
  NOR2_X1 U1549 ( .A1(n188), .A2(n283), .ZN(\p[15][34] ) );
  NOR2_X1 U1550 ( .A1(n176), .A2(n292), .ZN(\p[12][35] ) );
  NOR2_X1 U1551 ( .A1(n185), .A2(n283), .ZN(\p[15][35] ) );
  NOR2_X1 U1552 ( .A1(n173), .A2(n292), .ZN(\p[12][36] ) );
  NOR2_X1 U1553 ( .A1(n182), .A2(n283), .ZN(\p[15][36] ) );
  NOR2_X1 U1554 ( .A1(n170), .A2(n292), .ZN(\p[12][37] ) );
  NOR2_X1 U1555 ( .A1(n179), .A2(n283), .ZN(\p[15][37] ) );
  NOR2_X1 U1556 ( .A1(n167), .A2(n292), .ZN(\p[12][38] ) );
  NOR2_X1 U1557 ( .A1(n176), .A2(n283), .ZN(\p[15][38] ) );
  NOR2_X1 U1558 ( .A1(n164), .A2(n295), .ZN(\p[11][38] ) );
  NOR2_X1 U1559 ( .A1(n164), .A2(n292), .ZN(\p[12][39] ) );
  NOR2_X1 U1560 ( .A1(n191), .A2(n299), .ZN(\p[10][28] ) );
  NOR2_X1 U1561 ( .A1(n200), .A2(n290), .ZN(\p[13][28] ) );
  NOR2_X1 U1562 ( .A1(n188), .A2(n298), .ZN(\p[10][29] ) );
  NOR2_X1 U1563 ( .A1(n197), .A2(n290), .ZN(\p[13][29] ) );
  NOR2_X1 U1564 ( .A1(n185), .A2(n298), .ZN(\p[10][30] ) );
  NOR2_X1 U1565 ( .A1(n194), .A2(n290), .ZN(\p[13][30] ) );
  NOR2_X1 U1566 ( .A1(n182), .A2(n298), .ZN(\p[10][31] ) );
  NOR2_X1 U1567 ( .A1(n191), .A2(n290), .ZN(\p[13][31] ) );
  NOR2_X1 U1568 ( .A1(n179), .A2(n298), .ZN(\p[10][32] ) );
  NOR2_X1 U1569 ( .A1(n188), .A2(n289), .ZN(\p[13][32] ) );
  NOR2_X1 U1570 ( .A1(n185), .A2(n289), .ZN(\p[13][33] ) );
  NOR2_X1 U1571 ( .A1(n176), .A2(n298), .ZN(\p[10][33] ) );
  NOR2_X1 U1572 ( .A1(n182), .A2(n289), .ZN(\p[13][34] ) );
  NOR2_X1 U1573 ( .A1(n173), .A2(n298), .ZN(\p[10][34] ) );
  NOR2_X1 U1574 ( .A1(n179), .A2(n289), .ZN(\p[13][35] ) );
  NOR2_X1 U1575 ( .A1(n170), .A2(n298), .ZN(\p[10][35] ) );
  NOR2_X1 U1576 ( .A1(n176), .A2(n289), .ZN(\p[13][36] ) );
  NOR2_X1 U1577 ( .A1(n167), .A2(n298), .ZN(\p[10][36] ) );
  NOR2_X1 U1578 ( .A1(n173), .A2(n289), .ZN(\p[13][37] ) );
  NOR2_X1 U1579 ( .A1(n170), .A2(n289), .ZN(\p[13][38] ) );
  NOR2_X1 U1580 ( .A1(n167), .A2(n289), .ZN(\p[13][39] ) );
  NOR2_X1 U1581 ( .A1(n226), .A2(n261), .ZN(\p[23][27] ) );
  NOR2_X1 U1582 ( .A1(n137), .A2(n252), .ZN(\p[26][30] ) );
  NOR2_X1 U1583 ( .A1(n226), .A2(n243), .ZN(\p[29][33] ) );
  NOR2_X1 U1584 ( .A1(n236), .A2(n252), .ZN(\p[26][26] ) );
  NOR2_X1 U1585 ( .A1(n236), .A2(n243), .ZN(\p[29][29] ) );
  NOR2_X1 U1586 ( .A1(n227), .A2(n258), .ZN(\p[24][28] ) );
  NOR2_X1 U1587 ( .A1(n137), .A2(n249), .ZN(\p[27][31] ) );
  NOR2_X1 U1588 ( .A1(n227), .A2(n240), .ZN(\p[30][34] ) );
  NOR2_X1 U1589 ( .A1(n236), .A2(n240), .ZN(\p[30][30] ) );
  NOR2_X1 U1590 ( .A1(n164), .A2(n298), .ZN(\p[10][37] ) );
  NOR2_X1 U1591 ( .A1(n161), .A2(n298), .ZN(\p[10][38] ) );
  NOR2_X1 U1592 ( .A1(n158), .A2(n298), .ZN(\p[10][39] ) );
  NOR2_X1 U1593 ( .A1(n226), .A2(n255), .ZN(\p[25][29] ) );
  NOR2_X1 U1594 ( .A1(n227), .A2(n246), .ZN(\p[28][32] ) );
  NOR2_X1 U1595 ( .A1(n236), .A2(n246), .ZN(\p[28][28] ) );
  NOR2_X1 U1596 ( .A1(n234), .A2(n252), .ZN(\p[26][27] ) );
  NOR2_X1 U1597 ( .A1(n234), .A2(n249), .ZN(\p[27][28] ) );
  NOR2_X1 U1598 ( .A1(n234), .A2(n240), .ZN(\p[30][31] ) );
  NOR2_X1 U1599 ( .A1(n177), .A2(n308), .ZN(\p[5][27] ) );
  NOR2_X1 U1600 ( .A1(n174), .A2(n308), .ZN(\p[5][28] ) );
  NOR2_X1 U1601 ( .A1(n234), .A2(n255), .ZN(\p[25][26] ) );
  NOR2_X1 U1602 ( .A1(n234), .A2(n246), .ZN(\p[28][29] ) );
  NOR2_X1 U1603 ( .A1(n189), .A2(n304), .ZN(\p[8][26] ) );
  NOR2_X1 U1604 ( .A1(n216), .A2(n278), .ZN(\p[17][26] ) );
  NOR2_X1 U1605 ( .A1(n186), .A2(n304), .ZN(\p[8][27] ) );
  NOR2_X1 U1606 ( .A1(n214), .A2(n278), .ZN(\p[17][27] ) );
  NOR2_X1 U1607 ( .A1(n183), .A2(n304), .ZN(\p[8][28] ) );
  NOR2_X1 U1608 ( .A1(n211), .A2(n278), .ZN(\p[17][28] ) );
  NOR2_X1 U1609 ( .A1(n216), .A2(n269), .ZN(\p[20][29] ) );
  NOR2_X1 U1610 ( .A1(n180), .A2(n303), .ZN(\p[8][29] ) );
  NOR2_X1 U1611 ( .A1(n208), .A2(n278), .ZN(\p[17][29] ) );
  NOR2_X1 U1612 ( .A1(n205), .A2(n278), .ZN(\p[17][30] ) );
  NOR2_X1 U1613 ( .A1(n214), .A2(n269), .ZN(\p[20][30] ) );
  NOR2_X1 U1614 ( .A1(n211), .A2(n269), .ZN(\p[20][31] ) );
  NOR2_X1 U1615 ( .A1(n202), .A2(n278), .ZN(\p[17][31] ) );
  NOR2_X1 U1616 ( .A1(n217), .A2(n260), .ZN(\p[23][32] ) );
  NOR2_X1 U1617 ( .A1(n208), .A2(n269), .ZN(\p[20][32] ) );
  NOR2_X1 U1618 ( .A1(n199), .A2(n278), .ZN(\p[17][32] ) );
  NOR2_X1 U1619 ( .A1(n214), .A2(n260), .ZN(\p[23][33] ) );
  NOR2_X1 U1620 ( .A1(n205), .A2(n269), .ZN(\p[20][33] ) );
  NOR2_X1 U1621 ( .A1(n196), .A2(n278), .ZN(\p[17][33] ) );
  NOR2_X1 U1622 ( .A1(n211), .A2(n260), .ZN(\p[23][34] ) );
  NOR2_X1 U1623 ( .A1(n202), .A2(n269), .ZN(\p[20][34] ) );
  NOR2_X1 U1624 ( .A1(n193), .A2(n278), .ZN(\p[17][34] ) );
  NOR2_X1 U1625 ( .A1(n208), .A2(n260), .ZN(\p[23][35] ) );
  NOR2_X1 U1626 ( .A1(n199), .A2(n269), .ZN(\p[20][35] ) );
  NOR2_X1 U1627 ( .A1(n190), .A2(n278), .ZN(\p[17][35] ) );
  NOR2_X1 U1628 ( .A1(n216), .A2(n251), .ZN(\p[26][35] ) );
  NOR2_X1 U1629 ( .A1(n205), .A2(n260), .ZN(\p[23][36] ) );
  NOR2_X1 U1630 ( .A1(n196), .A2(n269), .ZN(\p[20][36] ) );
  NOR2_X1 U1631 ( .A1(n187), .A2(n277), .ZN(\p[17][36] ) );
  NOR2_X1 U1632 ( .A1(n214), .A2(n251), .ZN(\p[26][36] ) );
  NOR2_X1 U1633 ( .A1(n202), .A2(n260), .ZN(\p[23][37] ) );
  NOR2_X1 U1634 ( .A1(n193), .A2(n269), .ZN(\p[20][37] ) );
  NOR2_X1 U1635 ( .A1(n184), .A2(n277), .ZN(\p[17][37] ) );
  NOR2_X1 U1636 ( .A1(n216), .A2(n242), .ZN(\p[29][38] ) );
  NOR2_X1 U1637 ( .A1(n177), .A2(n303), .ZN(\p[8][30] ) );
  NOR2_X1 U1638 ( .A1(n174), .A2(n303), .ZN(\p[8][31] ) );
  NOR2_X1 U1639 ( .A1(n171), .A2(n311), .ZN(\p[4][28] ) );
  NOR2_X1 U1640 ( .A1(n183), .A2(n307), .ZN(\p[7][27] ) );
  NOR2_X1 U1641 ( .A1(n171), .A2(n303), .ZN(\p[8][32] ) );
  NOR2_X1 U1642 ( .A1(n168), .A2(n313), .ZN(\p[2][27] ) );
  NOR2_X1 U1643 ( .A1(n168), .A2(n303), .ZN(\p[8][33] ) );
  NOR2_X1 U1644 ( .A1(n165), .A2(n313), .ZN(\p[2][28] ) );
  NOR2_X1 U1645 ( .A1(n165), .A2(n303), .ZN(\p[8][34] ) );
  NOR2_X1 U1646 ( .A1(n162), .A2(n303), .ZN(\p[8][35] ) );
  NOR2_X1 U1647 ( .A1(n159), .A2(n303), .ZN(\p[8][36] ) );
  NOR2_X1 U1648 ( .A1(n156), .A2(n303), .ZN(\p[8][37] ) );
  NOR2_X1 U1649 ( .A1(n301), .A2(n186), .ZN(\p[9][28] ) );
  NOR2_X1 U1650 ( .A1(n216), .A2(n275), .ZN(\p[18][27] ) );
  NOR2_X1 U1651 ( .A1(n214), .A2(n275), .ZN(\p[18][28] ) );
  NOR2_X1 U1652 ( .A1(n211), .A2(n275), .ZN(\p[18][29] ) );
  NOR2_X1 U1653 ( .A1(n216), .A2(n266), .ZN(\p[21][30] ) );
  NOR2_X1 U1654 ( .A1(n208), .A2(n275), .ZN(\p[18][30] ) );
  NOR2_X1 U1655 ( .A1(n214), .A2(n266), .ZN(\p[21][31] ) );
  NOR2_X1 U1656 ( .A1(n205), .A2(n275), .ZN(\p[18][31] ) );
  NOR2_X1 U1657 ( .A1(n211), .A2(n266), .ZN(\p[21][32] ) );
  NOR2_X1 U1658 ( .A1(n202), .A2(n275), .ZN(\p[18][32] ) );
  NOR2_X1 U1659 ( .A1(n208), .A2(n266), .ZN(\p[21][33] ) );
  NOR2_X1 U1660 ( .A1(n199), .A2(n275), .ZN(\p[18][33] ) );
  NOR2_X1 U1661 ( .A1(n216), .A2(n257), .ZN(\p[24][33] ) );
  NOR2_X1 U1662 ( .A1(n205), .A2(n266), .ZN(\p[21][34] ) );
  NOR2_X1 U1663 ( .A1(n196), .A2(n275), .ZN(\p[18][34] ) );
  NOR2_X1 U1664 ( .A1(n214), .A2(n257), .ZN(\p[24][34] ) );
  NOR2_X1 U1665 ( .A1(n202), .A2(n266), .ZN(\p[21][35] ) );
  NOR2_X1 U1666 ( .A1(n193), .A2(n275), .ZN(\p[18][35] ) );
  NOR2_X1 U1667 ( .A1(n211), .A2(n257), .ZN(\p[24][35] ) );
  NOR2_X1 U1668 ( .A1(n216), .A2(n248), .ZN(\p[27][36] ) );
  NOR2_X1 U1669 ( .A1(n199), .A2(n266), .ZN(\p[21][36] ) );
  NOR2_X1 U1670 ( .A1(n190), .A2(n275), .ZN(\p[18][36] ) );
  NOR2_X1 U1671 ( .A1(n208), .A2(n257), .ZN(\p[24][36] ) );
  NOR2_X1 U1672 ( .A1(n213), .A2(n248), .ZN(\p[27][37] ) );
  NOR2_X1 U1673 ( .A1(n196), .A2(n266), .ZN(\p[21][37] ) );
  NOR2_X1 U1674 ( .A1(n187), .A2(n274), .ZN(\p[18][37] ) );
  NOR2_X1 U1675 ( .A1(n205), .A2(n257), .ZN(\p[24][37] ) );
  NOR2_X1 U1676 ( .A1(n210), .A2(n248), .ZN(\p[27][38] ) );
  NOR2_X1 U1677 ( .A1(n193), .A2(n266), .ZN(\p[21][38] ) );
  NOR2_X1 U1678 ( .A1(n184), .A2(n274), .ZN(\p[18][38] ) );
  NOR2_X1 U1679 ( .A1(n217), .A2(n239), .ZN(\p[30][39] ) );
  NOR2_X1 U1680 ( .A1(n207), .A2(n248), .ZN(\p[27][39] ) );
  NOR2_X1 U1681 ( .A1(n301), .A2(n183), .ZN(\p[9][29] ) );
  NOR2_X1 U1682 ( .A1(n301), .A2(n180), .ZN(\p[9][30] ) );
  NOR2_X1 U1683 ( .A1(n301), .A2(n177), .ZN(\p[9][31] ) );
  NOR2_X1 U1684 ( .A1(n301), .A2(n174), .ZN(\p[9][32] ) );
  NOR2_X1 U1685 ( .A1(n301), .A2(n171), .ZN(\p[9][33] ) );
  NOR2_X1 U1686 ( .A1(n301), .A2(n168), .ZN(\p[9][34] ) );
  NOR2_X1 U1687 ( .A1(n301), .A2(n165), .ZN(\p[9][35] ) );
  NOR2_X1 U1688 ( .A1(n301), .A2(n162), .ZN(\p[9][36] ) );
  NOR2_X1 U1689 ( .A1(n301), .A2(n159), .ZN(\p[9][37] ) );
  NOR2_X1 U1690 ( .A1(n301), .A2(n156), .ZN(\p[9][38] ) );
  NOR2_X1 U1691 ( .A1(n301), .A2(n153), .ZN(\p[9][39] ) );
  NOR2_X1 U1692 ( .A1(n211), .A2(n281), .ZN(\p[16][27] ) );
  NOR2_X1 U1693 ( .A1(n217), .A2(n272), .ZN(\p[19][28] ) );
  NOR2_X1 U1694 ( .A1(n208), .A2(n281), .ZN(\p[16][28] ) );
  NOR2_X1 U1695 ( .A1(n214), .A2(n272), .ZN(\p[19][29] ) );
  NOR2_X1 U1696 ( .A1(n205), .A2(n281), .ZN(\p[16][29] ) );
  NOR2_X1 U1697 ( .A1(n202), .A2(n281), .ZN(\p[16][30] ) );
  NOR2_X1 U1698 ( .A1(n211), .A2(n272), .ZN(\p[19][30] ) );
  NOR2_X1 U1699 ( .A1(n216), .A2(n263), .ZN(\p[22][31] ) );
  NOR2_X1 U1700 ( .A1(n208), .A2(n272), .ZN(\p[19][31] ) );
  NOR2_X1 U1701 ( .A1(n199), .A2(n281), .ZN(\p[16][31] ) );
  NOR2_X1 U1702 ( .A1(n214), .A2(n263), .ZN(\p[22][32] ) );
  NOR2_X1 U1703 ( .A1(n205), .A2(n272), .ZN(\p[19][32] ) );
  NOR2_X1 U1704 ( .A1(n196), .A2(n281), .ZN(\p[16][32] ) );
  NOR2_X1 U1705 ( .A1(n211), .A2(n263), .ZN(\p[22][33] ) );
  NOR2_X1 U1706 ( .A1(n202), .A2(n272), .ZN(\p[19][33] ) );
  NOR2_X1 U1707 ( .A1(n193), .A2(n281), .ZN(\p[16][33] ) );
  NOR2_X1 U1708 ( .A1(n208), .A2(n263), .ZN(\p[22][34] ) );
  NOR2_X1 U1709 ( .A1(n199), .A2(n272), .ZN(\p[19][34] ) );
  NOR2_X1 U1710 ( .A1(n190), .A2(n281), .ZN(\p[16][34] ) );
  NOR2_X1 U1711 ( .A1(n216), .A2(n254), .ZN(\p[25][34] ) );
  NOR2_X1 U1712 ( .A1(n205), .A2(n263), .ZN(\p[22][35] ) );
  NOR2_X1 U1713 ( .A1(n196), .A2(n272), .ZN(\p[19][35] ) );
  NOR2_X1 U1714 ( .A1(n187), .A2(n280), .ZN(\p[16][35] ) );
  NOR2_X1 U1715 ( .A1(n214), .A2(n254), .ZN(\p[25][35] ) );
  NOR2_X1 U1716 ( .A1(n202), .A2(n263), .ZN(\p[22][36] ) );
  NOR2_X1 U1717 ( .A1(n193), .A2(n272), .ZN(\p[19][36] ) );
  NOR2_X1 U1718 ( .A1(n184), .A2(n280), .ZN(\p[16][36] ) );
  NOR2_X1 U1719 ( .A1(n211), .A2(n254), .ZN(\p[25][36] ) );
  NOR2_X1 U1720 ( .A1(n217), .A2(n245), .ZN(\p[28][37] ) );
  NOR2_X1 U1721 ( .A1(n199), .A2(n263), .ZN(\p[22][37] ) );
  NOR2_X1 U1722 ( .A1(n190), .A2(n272), .ZN(\p[19][37] ) );
  NOR2_X1 U1723 ( .A1(n181), .A2(n280), .ZN(\p[16][37] ) );
  NOR2_X1 U1724 ( .A1(n208), .A2(n254), .ZN(\p[25][37] ) );
  NOR2_X1 U1725 ( .A1(n213), .A2(n245), .ZN(\p[28][38] ) );
  NOR2_X1 U1726 ( .A1(n196), .A2(n263), .ZN(\p[22][38] ) );
  NOR2_X1 U1727 ( .A1(n187), .A2(n271), .ZN(\p[19][38] ) );
  NOR2_X1 U1728 ( .A1(n178), .A2(n280), .ZN(\p[16][38] ) );
  NOR2_X1 U1729 ( .A1(n210), .A2(n245), .ZN(\p[28][39] ) );
  BUF_X1 U1730 ( .A(\p[57][63] ), .Z(n389) );
  BUF_X2 U1731 ( .A(\p[0][63] ), .Z(n409) );
  BUF_X2 U1732 ( .A(\p[3][63] ), .Z(n418) );
  BUF_X2 U1733 ( .A(\p[6][63] ), .Z(n427) );
  BUF_X2 U1734 ( .A(\p[4][63] ), .Z(n421) );
  BUF_X2 U1735 ( .A(\p[1][63] ), .Z(n412) );
  NOR2_X1 U1736 ( .A1(n170), .A2(n286), .ZN(\p[14][39] ) );
  NOR2_X1 U1737 ( .A1(n167), .A2(n286), .ZN(\p[14][40] ) );
  NOR2_X1 U1738 ( .A1(n173), .A2(n283), .ZN(\p[15][39] ) );
  NOR2_X1 U1739 ( .A1(n170), .A2(n283), .ZN(\p[15][40] ) );
  NOR2_X1 U1740 ( .A1(n167), .A2(n283), .ZN(\p[15][41] ) );
  NOR2_X1 U1741 ( .A1(n161), .A2(n295), .ZN(\p[11][39] ) );
  NOR2_X1 U1742 ( .A1(n158), .A2(n295), .ZN(\p[11][40] ) );
  NOR2_X1 U1743 ( .A1(n155), .A2(n295), .ZN(\p[11][41] ) );
  NOR2_X1 U1744 ( .A1(n164), .A2(n286), .ZN(\p[14][41] ) );
  NOR2_X1 U1745 ( .A1(n161), .A2(n286), .ZN(\p[14][42] ) );
  NOR2_X1 U1746 ( .A1(n158), .A2(n286), .ZN(\p[14][43] ) );
  NOR2_X1 U1747 ( .A1(n155), .A2(n286), .ZN(\p[14][44] ) );
  NOR2_X1 U1748 ( .A1(n161), .A2(n292), .ZN(\p[12][40] ) );
  NOR2_X1 U1749 ( .A1(n158), .A2(n292), .ZN(\p[12][41] ) );
  NOR2_X1 U1750 ( .A1(n155), .A2(n292), .ZN(\p[12][42] ) );
  NOR2_X1 U1751 ( .A1(n164), .A2(n283), .ZN(\p[15][42] ) );
  NOR2_X1 U1752 ( .A1(n161), .A2(n283), .ZN(\p[15][43] ) );
  NOR2_X1 U1753 ( .A1(n158), .A2(n283), .ZN(\p[15][44] ) );
  NOR2_X1 U1754 ( .A1(n155), .A2(n283), .ZN(\p[15][45] ) );
  NOR2_X1 U1755 ( .A1(n155), .A2(n298), .ZN(\p[10][40] ) );
  NOR2_X1 U1756 ( .A1(n164), .A2(n289), .ZN(\p[13][40] ) );
  NOR2_X1 U1757 ( .A1(n161), .A2(n289), .ZN(\p[13][41] ) );
  NOR2_X1 U1758 ( .A1(n158), .A2(n289), .ZN(\p[13][42] ) );
  NOR2_X1 U1759 ( .A1(n155), .A2(n289), .ZN(\p[13][43] ) );
  NOR2_X1 U1760 ( .A1(n211), .A2(n251), .ZN(\p[26][37] ) );
  NOR2_X1 U1761 ( .A1(n199), .A2(n260), .ZN(\p[23][38] ) );
  NOR2_X1 U1762 ( .A1(n190), .A2(n269), .ZN(\p[20][38] ) );
  NOR2_X1 U1763 ( .A1(n181), .A2(n277), .ZN(\p[17][38] ) );
  NOR2_X1 U1764 ( .A1(n208), .A2(n251), .ZN(\p[26][38] ) );
  NOR2_X1 U1765 ( .A1(n213), .A2(n242), .ZN(\p[29][39] ) );
  NOR2_X1 U1766 ( .A1(n196), .A2(n260), .ZN(\p[23][39] ) );
  NOR2_X1 U1767 ( .A1(n187), .A2(n268), .ZN(\p[20][39] ) );
  NOR2_X1 U1768 ( .A1(n178), .A2(n277), .ZN(\p[17][39] ) );
  NOR2_X1 U1769 ( .A1(n205), .A2(n251), .ZN(\p[26][39] ) );
  NOR2_X1 U1770 ( .A1(n210), .A2(n242), .ZN(\p[29][40] ) );
  NOR2_X1 U1771 ( .A1(n193), .A2(n260), .ZN(\p[23][40] ) );
  NOR2_X1 U1772 ( .A1(n184), .A2(n268), .ZN(\p[20][40] ) );
  NOR2_X1 U1773 ( .A1(n175), .A2(n277), .ZN(\p[17][40] ) );
  NOR2_X1 U1774 ( .A1(n202), .A2(n251), .ZN(\p[26][40] ) );
  NOR2_X1 U1775 ( .A1(n207), .A2(n242), .ZN(\p[29][41] ) );
  NOR2_X1 U1776 ( .A1(n190), .A2(n260), .ZN(\p[23][41] ) );
  NOR2_X1 U1777 ( .A1(n181), .A2(n268), .ZN(\p[20][41] ) );
  NOR2_X1 U1778 ( .A1(n172), .A2(n277), .ZN(\p[17][41] ) );
  NOR2_X1 U1779 ( .A1(n199), .A2(n251), .ZN(\p[26][41] ) );
  NOR2_X1 U1780 ( .A1(n204), .A2(n242), .ZN(\p[29][42] ) );
  NOR2_X1 U1781 ( .A1(n187), .A2(n259), .ZN(\p[23][42] ) );
  NOR2_X1 U1782 ( .A1(n178), .A2(n268), .ZN(\p[20][42] ) );
  NOR2_X1 U1783 ( .A1(n169), .A2(n277), .ZN(\p[17][42] ) );
  NOR2_X1 U1784 ( .A1(n196), .A2(n251), .ZN(\p[26][42] ) );
  NOR2_X1 U1785 ( .A1(n201), .A2(n242), .ZN(\p[29][43] ) );
  NOR2_X1 U1786 ( .A1(n184), .A2(n259), .ZN(\p[23][43] ) );
  NOR2_X1 U1787 ( .A1(n175), .A2(n268), .ZN(\p[20][43] ) );
  NOR2_X1 U1788 ( .A1(n166), .A2(n277), .ZN(\p[17][43] ) );
  NOR2_X1 U1789 ( .A1(n193), .A2(n251), .ZN(\p[26][43] ) );
  NOR2_X1 U1790 ( .A1(n198), .A2(n242), .ZN(\p[29][44] ) );
  NOR2_X1 U1791 ( .A1(n181), .A2(n259), .ZN(\p[23][44] ) );
  NOR2_X1 U1792 ( .A1(n172), .A2(n268), .ZN(\p[20][44] ) );
  NOR2_X1 U1793 ( .A1(n190), .A2(n251), .ZN(\p[26][44] ) );
  NOR2_X1 U1794 ( .A1(n195), .A2(n242), .ZN(\p[29][45] ) );
  NOR2_X1 U1795 ( .A1(n178), .A2(n259), .ZN(\p[23][45] ) );
  NOR2_X1 U1796 ( .A1(n169), .A2(n268), .ZN(\p[20][45] ) );
  NOR2_X1 U1797 ( .A1(n187), .A2(n250), .ZN(\p[26][45] ) );
  NOR2_X1 U1798 ( .A1(n192), .A2(n242), .ZN(\p[29][46] ) );
  NOR2_X1 U1799 ( .A1(n175), .A2(n259), .ZN(\p[23][46] ) );
  NOR2_X1 U1800 ( .A1(n166), .A2(n268), .ZN(\p[20][46] ) );
  NOR2_X1 U1801 ( .A1(n184), .A2(n250), .ZN(\p[26][46] ) );
  NOR2_X1 U1802 ( .A1(n189), .A2(n242), .ZN(\p[29][47] ) );
  NOR2_X1 U1803 ( .A1(n172), .A2(n259), .ZN(\p[23][47] ) );
  NOR2_X1 U1804 ( .A1(n181), .A2(n250), .ZN(\p[26][47] ) );
  NOR2_X1 U1805 ( .A1(n186), .A2(n241), .ZN(\p[29][48] ) );
  NOR2_X1 U1806 ( .A1(n169), .A2(n259), .ZN(\p[23][48] ) );
  NOR2_X1 U1807 ( .A1(n178), .A2(n250), .ZN(\p[26][48] ) );
  NOR2_X1 U1808 ( .A1(n166), .A2(n259), .ZN(\p[23][49] ) );
  NOR2_X1 U1809 ( .A1(n183), .A2(n241), .ZN(\p[29][49] ) );
  NOR2_X1 U1810 ( .A1(n180), .A2(n241), .ZN(\p[29][50] ) );
  NOR2_X1 U1811 ( .A1(n163), .A2(n277), .ZN(\p[17][44] ) );
  NOR2_X1 U1812 ( .A1(n160), .A2(n277), .ZN(\p[17][45] ) );
  NOR2_X1 U1813 ( .A1(n157), .A2(n277), .ZN(\p[17][46] ) );
  NOR2_X1 U1814 ( .A1(n163), .A2(n268), .ZN(\p[20][47] ) );
  NOR2_X1 U1815 ( .A1(n154), .A2(n277), .ZN(\p[17][47] ) );
  NOR2_X1 U1816 ( .A1(n160), .A2(n268), .ZN(\p[20][48] ) );
  NOR2_X1 U1817 ( .A1(n157), .A2(n268), .ZN(\p[20][49] ) );
  NOR2_X1 U1818 ( .A1(n153), .A2(n303), .ZN(\p[8][38] ) );
  NOR2_X1 U1819 ( .A1(n202), .A2(n257), .ZN(\p[24][38] ) );
  NOR2_X1 U1820 ( .A1(n190), .A2(n266), .ZN(\p[21][39] ) );
  NOR2_X1 U1821 ( .A1(n181), .A2(n274), .ZN(\p[18][39] ) );
  NOR2_X1 U1822 ( .A1(n199), .A2(n257), .ZN(\p[24][39] ) );
  NOR2_X1 U1823 ( .A1(n213), .A2(n239), .ZN(\p[30][40] ) );
  NOR2_X1 U1824 ( .A1(n204), .A2(n248), .ZN(\p[27][40] ) );
  NOR2_X1 U1825 ( .A1(n187), .A2(n265), .ZN(\p[21][40] ) );
  NOR2_X1 U1826 ( .A1(n178), .A2(n274), .ZN(\p[18][40] ) );
  NOR2_X1 U1827 ( .A1(n196), .A2(n257), .ZN(\p[24][40] ) );
  NOR2_X1 U1828 ( .A1(n210), .A2(n239), .ZN(\p[30][41] ) );
  NOR2_X1 U1829 ( .A1(n201), .A2(n248), .ZN(\p[27][41] ) );
  NOR2_X1 U1830 ( .A1(n184), .A2(n265), .ZN(\p[21][41] ) );
  NOR2_X1 U1831 ( .A1(n175), .A2(n274), .ZN(\p[18][41] ) );
  NOR2_X1 U1832 ( .A1(n193), .A2(n257), .ZN(\p[24][41] ) );
  NOR2_X1 U1833 ( .A1(n207), .A2(n239), .ZN(\p[30][42] ) );
  NOR2_X1 U1834 ( .A1(n198), .A2(n248), .ZN(\p[27][42] ) );
  NOR2_X1 U1835 ( .A1(n181), .A2(n265), .ZN(\p[21][42] ) );
  NOR2_X1 U1836 ( .A1(n172), .A2(n274), .ZN(\p[18][42] ) );
  NOR2_X1 U1837 ( .A1(n190), .A2(n257), .ZN(\p[24][42] ) );
  NOR2_X1 U1838 ( .A1(n204), .A2(n239), .ZN(\p[30][43] ) );
  NOR2_X1 U1839 ( .A1(n195), .A2(n248), .ZN(\p[27][43] ) );
  NOR2_X1 U1840 ( .A1(n178), .A2(n265), .ZN(\p[21][43] ) );
  NOR2_X1 U1841 ( .A1(n169), .A2(n274), .ZN(\p[18][43] ) );
  NOR2_X1 U1842 ( .A1(n187), .A2(n256), .ZN(\p[24][43] ) );
  NOR2_X1 U1843 ( .A1(n201), .A2(n239), .ZN(\p[30][44] ) );
  NOR2_X1 U1844 ( .A1(n192), .A2(n248), .ZN(\p[27][44] ) );
  NOR2_X1 U1845 ( .A1(n175), .A2(n265), .ZN(\p[21][44] ) );
  NOR2_X1 U1846 ( .A1(n166), .A2(n274), .ZN(\p[18][44] ) );
  NOR2_X1 U1847 ( .A1(n184), .A2(n256), .ZN(\p[24][44] ) );
  NOR2_X1 U1848 ( .A1(n198), .A2(n239), .ZN(\p[30][45] ) );
  NOR2_X1 U1849 ( .A1(n189), .A2(n248), .ZN(\p[27][45] ) );
  NOR2_X1 U1850 ( .A1(n172), .A2(n265), .ZN(\p[21][45] ) );
  NOR2_X1 U1851 ( .A1(n181), .A2(n256), .ZN(\p[24][45] ) );
  NOR2_X1 U1852 ( .A1(n195), .A2(n239), .ZN(\p[30][46] ) );
  NOR2_X1 U1853 ( .A1(n186), .A2(n247), .ZN(\p[27][46] ) );
  NOR2_X1 U1854 ( .A1(n169), .A2(n265), .ZN(\p[21][46] ) );
  NOR2_X1 U1855 ( .A1(n178), .A2(n256), .ZN(\p[24][46] ) );
  NOR2_X1 U1856 ( .A1(n192), .A2(n239), .ZN(\p[30][47] ) );
  NOR2_X1 U1857 ( .A1(n183), .A2(n247), .ZN(\p[27][47] ) );
  NOR2_X1 U1858 ( .A1(n166), .A2(n265), .ZN(\p[21][47] ) );
  NOR2_X1 U1859 ( .A1(n175), .A2(n256), .ZN(\p[24][47] ) );
  NOR2_X1 U1860 ( .A1(n189), .A2(n239), .ZN(\p[30][48] ) );
  NOR2_X1 U1861 ( .A1(n180), .A2(n247), .ZN(\p[27][48] ) );
  NOR2_X1 U1862 ( .A1(n172), .A2(n256), .ZN(\p[24][48] ) );
  NOR2_X1 U1863 ( .A1(n186), .A2(n238), .ZN(\p[30][49] ) );
  NOR2_X1 U1864 ( .A1(n169), .A2(n256), .ZN(\p[24][49] ) );
  NOR2_X1 U1865 ( .A1(n183), .A2(n238), .ZN(\p[30][50] ) );
  NOR2_X1 U1866 ( .A1(n180), .A2(n238), .ZN(\p[30][51] ) );
  NOR2_X1 U1867 ( .A1(n163), .A2(n274), .ZN(\p[18][45] ) );
  NOR2_X1 U1868 ( .A1(n160), .A2(n274), .ZN(\p[18][46] ) );
  NOR2_X1 U1869 ( .A1(n157), .A2(n274), .ZN(\p[18][47] ) );
  NOR2_X1 U1870 ( .A1(n163), .A2(n265), .ZN(\p[21][48] ) );
  NOR2_X1 U1871 ( .A1(n154), .A2(n274), .ZN(\p[18][48] ) );
  NOR2_X1 U1872 ( .A1(n160), .A2(n265), .ZN(\p[21][49] ) );
  NOR2_X1 U1873 ( .A1(n177), .A2(n247), .ZN(\p[27][49] ) );
  NOR2_X1 U1874 ( .A1(n174), .A2(n247), .ZN(\p[27][50] ) );
  NOR2_X1 U1875 ( .A1(n157), .A2(n265), .ZN(\p[21][50] ) );
  NOR2_X1 U1876 ( .A1(n171), .A2(n247), .ZN(\p[27][51] ) );
  NOR2_X1 U1877 ( .A1(n205), .A2(n254), .ZN(\p[25][38] ) );
  NOR2_X1 U1878 ( .A1(n193), .A2(n263), .ZN(\p[22][39] ) );
  NOR2_X1 U1879 ( .A1(n184), .A2(n271), .ZN(\p[19][39] ) );
  NOR2_X1 U1880 ( .A1(n175), .A2(n280), .ZN(\p[16][39] ) );
  NOR2_X1 U1881 ( .A1(n202), .A2(n254), .ZN(\p[25][39] ) );
  NOR2_X1 U1882 ( .A1(n207), .A2(n245), .ZN(\p[28][40] ) );
  NOR2_X1 U1883 ( .A1(n190), .A2(n263), .ZN(\p[22][40] ) );
  NOR2_X1 U1884 ( .A1(n181), .A2(n271), .ZN(\p[19][40] ) );
  NOR2_X1 U1885 ( .A1(n172), .A2(n280), .ZN(\p[16][40] ) );
  NOR2_X1 U1886 ( .A1(n199), .A2(n254), .ZN(\p[25][40] ) );
  NOR2_X1 U1887 ( .A1(n204), .A2(n245), .ZN(\p[28][41] ) );
  NOR2_X1 U1888 ( .A1(n187), .A2(n262), .ZN(\p[22][41] ) );
  NOR2_X1 U1889 ( .A1(n178), .A2(n271), .ZN(\p[19][41] ) );
  NOR2_X1 U1890 ( .A1(n169), .A2(n280), .ZN(\p[16][41] ) );
  NOR2_X1 U1891 ( .A1(n196), .A2(n254), .ZN(\p[25][41] ) );
  NOR2_X1 U1892 ( .A1(n201), .A2(n245), .ZN(\p[28][42] ) );
  NOR2_X1 U1893 ( .A1(n184), .A2(n262), .ZN(\p[22][42] ) );
  NOR2_X1 U1894 ( .A1(n175), .A2(n271), .ZN(\p[19][42] ) );
  NOR2_X1 U1895 ( .A1(n166), .A2(n280), .ZN(\p[16][42] ) );
  NOR2_X1 U1896 ( .A1(n193), .A2(n254), .ZN(\p[25][42] ) );
  NOR2_X1 U1897 ( .A1(n198), .A2(n245), .ZN(\p[28][43] ) );
  NOR2_X1 U1898 ( .A1(n181), .A2(n262), .ZN(\p[22][43] ) );
  NOR2_X1 U1899 ( .A1(n172), .A2(n271), .ZN(\p[19][43] ) );
  NOR2_X1 U1900 ( .A1(n190), .A2(n254), .ZN(\p[25][43] ) );
  NOR2_X1 U1901 ( .A1(n195), .A2(n245), .ZN(\p[28][44] ) );
  NOR2_X1 U1902 ( .A1(n178), .A2(n262), .ZN(\p[22][44] ) );
  NOR2_X1 U1903 ( .A1(n169), .A2(n271), .ZN(\p[19][44] ) );
  NOR2_X1 U1904 ( .A1(n187), .A2(n253), .ZN(\p[25][44] ) );
  NOR2_X1 U1905 ( .A1(n192), .A2(n245), .ZN(\p[28][45] ) );
  NOR2_X1 U1906 ( .A1(n175), .A2(n262), .ZN(\p[22][45] ) );
  NOR2_X1 U1907 ( .A1(n166), .A2(n271), .ZN(\p[19][45] ) );
  NOR2_X1 U1908 ( .A1(n184), .A2(n253), .ZN(\p[25][45] ) );
  NOR2_X1 U1909 ( .A1(n189), .A2(n245), .ZN(\p[28][46] ) );
  NOR2_X1 U1910 ( .A1(n172), .A2(n262), .ZN(\p[22][46] ) );
  NOR2_X1 U1911 ( .A1(n181), .A2(n253), .ZN(\p[25][46] ) );
  NOR2_X1 U1912 ( .A1(n186), .A2(n244), .ZN(\p[28][47] ) );
  NOR2_X1 U1913 ( .A1(n169), .A2(n262), .ZN(\p[22][47] ) );
  NOR2_X1 U1914 ( .A1(n178), .A2(n253), .ZN(\p[25][47] ) );
  NOR2_X1 U1915 ( .A1(n183), .A2(n244), .ZN(\p[28][48] ) );
  NOR2_X1 U1916 ( .A1(n166), .A2(n262), .ZN(\p[22][48] ) );
  NOR2_X1 U1917 ( .A1(n175), .A2(n253), .ZN(\p[25][48] ) );
  NOR2_X1 U1918 ( .A1(n180), .A2(n244), .ZN(\p[28][49] ) );
  NOR2_X1 U1919 ( .A1(n172), .A2(n253), .ZN(\p[25][49] ) );
  NOR2_X1 U1920 ( .A1(n163), .A2(n280), .ZN(\p[16][43] ) );
  NOR2_X1 U1921 ( .A1(n160), .A2(n280), .ZN(\p[16][44] ) );
  NOR2_X1 U1922 ( .A1(n157), .A2(n280), .ZN(\p[16][45] ) );
  NOR2_X1 U1923 ( .A1(n163), .A2(n271), .ZN(\p[19][46] ) );
  NOR2_X1 U1924 ( .A1(n154), .A2(n280), .ZN(\p[16][46] ) );
  NOR2_X1 U1925 ( .A1(n160), .A2(n271), .ZN(\p[19][47] ) );
  NOR2_X1 U1926 ( .A1(n157), .A2(n271), .ZN(\p[19][48] ) );
  NOR2_X1 U1927 ( .A1(n154), .A2(n271), .ZN(\p[19][49] ) );
  NOR2_X1 U1928 ( .A1(n163), .A2(n262), .ZN(\p[22][49] ) );
  NOR2_X1 U1929 ( .A1(n177), .A2(n244), .ZN(\p[28][50] ) );
  NOR2_X1 U1930 ( .A1(n160), .A2(n262), .ZN(\p[22][50] ) );
  NOR2_X1 U1931 ( .A1(n174), .A2(n244), .ZN(\p[28][51] ) );
  BUF_X1 U1932 ( .A(\p[56][63] ), .Z(n386) );
  BUF_X1 U1933 ( .A(\p[1][63] ), .Z(n413) );
  BUF_X1 U1934 ( .A(\p[3][63] ), .Z(n419) );
  BUF_X1 U1935 ( .A(\p[0][63] ), .Z(n410) );
  BUF_X1 U1936 ( .A(\p[4][63] ), .Z(n422) );
  NOR2_X1 U1937 ( .A1(n175), .A2(n250), .ZN(\p[26][49] ) );
  NOR2_X1 U1938 ( .A1(n172), .A2(n250), .ZN(\p[26][50] ) );
  NOR2_X1 U1939 ( .A1(n169), .A2(n250), .ZN(\p[26][51] ) );
  NOR2_X1 U1940 ( .A1(n166), .A2(n250), .ZN(\p[26][52] ) );
  NOR2_X1 U1941 ( .A1(n154), .A2(n268), .ZN(\p[20][50] ) );
  NOR2_X1 U1942 ( .A1(n163), .A2(n259), .ZN(\p[23][50] ) );
  NOR2_X1 U1943 ( .A1(n177), .A2(n241), .ZN(\p[29][51] ) );
  NOR2_X1 U1944 ( .A1(n160), .A2(n259), .ZN(\p[23][51] ) );
  NOR2_X1 U1945 ( .A1(n157), .A2(n259), .ZN(\p[23][52] ) );
  NOR2_X1 U1946 ( .A1(n174), .A2(n241), .ZN(\p[29][52] ) );
  NOR2_X1 U1947 ( .A1(n154), .A2(n259), .ZN(\p[23][53] ) );
  NOR2_X1 U1948 ( .A1(n163), .A2(n250), .ZN(\p[26][53] ) );
  NOR2_X1 U1949 ( .A1(n160), .A2(n250), .ZN(\p[26][54] ) );
  NOR2_X1 U1950 ( .A1(n157), .A2(n250), .ZN(\p[26][55] ) );
  NOR2_X1 U1951 ( .A1(n154), .A2(n250), .ZN(\p[26][56] ) );
  NOR2_X1 U1952 ( .A1(n171), .A2(n241), .ZN(\p[29][53] ) );
  NOR2_X1 U1953 ( .A1(n168), .A2(n241), .ZN(\p[29][54] ) );
  NOR2_X1 U1954 ( .A1(n165), .A2(n241), .ZN(\p[29][55] ) );
  NOR2_X1 U1955 ( .A1(n159), .A2(n241), .ZN(\p[29][57] ) );
  NOR2_X1 U1956 ( .A1(n156), .A2(n241), .ZN(\p[29][58] ) );
  NOR2_X1 U1957 ( .A1(n162), .A2(n241), .ZN(\p[29][56] ) );
  NOR2_X1 U1958 ( .A1(n153), .A2(n241), .ZN(\p[29][59] ) );
  NOR2_X1 U1959 ( .A1(n166), .A2(n256), .ZN(\p[24][50] ) );
  NOR2_X1 U1960 ( .A1(n154), .A2(n265), .ZN(\p[21][51] ) );
  NOR2_X1 U1961 ( .A1(n163), .A2(n256), .ZN(\p[24][51] ) );
  NOR2_X1 U1962 ( .A1(n177), .A2(n238), .ZN(\p[30][52] ) );
  NOR2_X1 U1963 ( .A1(n160), .A2(n256), .ZN(\p[24][52] ) );
  NOR2_X1 U1964 ( .A1(n174), .A2(n238), .ZN(\p[30][53] ) );
  NOR2_X1 U1965 ( .A1(n157), .A2(n256), .ZN(\p[24][53] ) );
  NOR2_X1 U1966 ( .A1(n154), .A2(n256), .ZN(\p[24][54] ) );
  NOR2_X1 U1967 ( .A1(n171), .A2(n238), .ZN(\p[30][54] ) );
  NOR2_X1 U1968 ( .A1(n168), .A2(n247), .ZN(\p[27][52] ) );
  NOR2_X1 U1969 ( .A1(n168), .A2(n238), .ZN(\p[30][55] ) );
  NOR2_X1 U1970 ( .A1(n165), .A2(n247), .ZN(\p[27][53] ) );
  NOR2_X1 U1971 ( .A1(n165), .A2(n238), .ZN(\p[30][56] ) );
  NOR2_X1 U1972 ( .A1(n162), .A2(n247), .ZN(\p[27][54] ) );
  NOR2_X1 U1973 ( .A1(n159), .A2(n247), .ZN(\p[27][55] ) );
  NOR2_X1 U1974 ( .A1(n162), .A2(n238), .ZN(\p[30][57] ) );
  NOR2_X1 U1975 ( .A1(n153), .A2(n247), .ZN(\p[27][57] ) );
  NOR2_X1 U1976 ( .A1(n159), .A2(n238), .ZN(\p[30][58] ) );
  NOR2_X1 U1977 ( .A1(n156), .A2(n247), .ZN(\p[27][56] ) );
  NOR2_X1 U1978 ( .A1(n156), .A2(n238), .ZN(\p[30][59] ) );
  NOR2_X1 U1979 ( .A1(n153), .A2(n238), .ZN(\p[30][60] ) );
  NOR2_X1 U1980 ( .A1(n169), .A2(n253), .ZN(\p[25][50] ) );
  NOR2_X1 U1981 ( .A1(n166), .A2(n253), .ZN(\p[25][51] ) );
  NOR2_X1 U1982 ( .A1(n157), .A2(n262), .ZN(\p[22][51] ) );
  NOR2_X1 U1983 ( .A1(n154), .A2(n262), .ZN(\p[22][52] ) );
  NOR2_X1 U1984 ( .A1(n163), .A2(n253), .ZN(\p[25][52] ) );
  NOR2_X1 U1985 ( .A1(n160), .A2(n253), .ZN(\p[25][53] ) );
  NOR2_X1 U1986 ( .A1(n157), .A2(n253), .ZN(\p[25][54] ) );
  NOR2_X1 U1987 ( .A1(n154), .A2(n253), .ZN(\p[25][55] ) );
  NOR2_X1 U1988 ( .A1(n171), .A2(n244), .ZN(\p[28][52] ) );
  NOR2_X1 U1989 ( .A1(n168), .A2(n244), .ZN(\p[28][53] ) );
  NOR2_X1 U1990 ( .A1(n165), .A2(n244), .ZN(\p[28][54] ) );
  NOR2_X1 U1991 ( .A1(n162), .A2(n244), .ZN(\p[28][55] ) );
  NOR2_X1 U1992 ( .A1(n156), .A2(n244), .ZN(\p[28][57] ) );
  NOR2_X1 U1993 ( .A1(n153), .A2(n244), .ZN(\p[28][58] ) );
  NOR2_X1 U1994 ( .A1(n159), .A2(n244), .ZN(\p[28][56] ) );
  BUF_X1 U1995 ( .A(\p[6][63] ), .Z(n428) );
  BUF_X2 U1996 ( .A(n110), .Z(n315) );
  BUF_X2 U1997 ( .A(n119), .Z(n307) );
  BUF_X2 U1998 ( .A(n443), .Z(n236) );
  BUF_X1 U1999 ( .A(n224), .Z(n225) );
  BUF_X1 U2000 ( .A(n93), .Z(n294) );
  BUF_X1 U2001 ( .A(n112), .Z(n300) );
  BUF_X1 U2002 ( .A(n118), .Z(n314) );
  BUF_X1 U2003 ( .A(n76), .Z(n194) );
  BUF_X1 U2004 ( .A(n73), .Z(n200) );
  BUF_X1 U2005 ( .A(n75), .Z(n197) );
  BUF_X1 U2006 ( .A(n90), .Z(n209) );
  BUF_X1 U2007 ( .A(n91), .Z(n212) );
  BUF_X1 U2008 ( .A(n69), .Z(n206) );
  BUF_X1 U2009 ( .A(n72), .Z(n203) );
  BUF_X1 U2010 ( .A(n70), .Z(n191) );
  BUF_X1 U2011 ( .A(n74), .Z(n188) );
  BUF_X1 U2012 ( .A(n71), .Z(n185) );
  BUF_X1 U2013 ( .A(n77), .Z(n182) );
  BUF_X1 U2014 ( .A(n79), .Z(n179) );
  BUF_X1 U2015 ( .A(n78), .Z(n176) );
  BUF_X1 U2016 ( .A(n94), .Z(n173) );
  BUF_X1 U2017 ( .A(n100), .Z(n170) );
  BUF_X1 U2018 ( .A(n99), .Z(n167) );
  BUF_X1 U2019 ( .A(n122), .Z(n309) );
  BUF_X1 U2020 ( .A(n87), .Z(n285) );
  BUF_X1 U2021 ( .A(n88), .Z(n288) );
  BUF_X1 U2022 ( .A(n92), .Z(n297) );
  BUF_X1 U2023 ( .A(n89), .Z(n291) );
  BUF_X1 U2024 ( .A(n85), .Z(n276) );
  BUF_X1 U2025 ( .A(n82), .Z(n267) );
  BUF_X1 U2026 ( .A(n104), .Z(n261) );
  BUF_X1 U2027 ( .A(n98), .Z(n164) );
  BUF_X1 U2028 ( .A(n86), .Z(n281) );
  BUF_X1 U2029 ( .A(n84), .Z(n278) );
  BUF_X1 U2030 ( .A(n85), .Z(n275) );
  BUF_X1 U2031 ( .A(n83), .Z(n272) );
  BUF_X1 U2032 ( .A(n86), .Z(n282) );
  BUF_X1 U2033 ( .A(n84), .Z(n279) );
  BUF_X1 U2034 ( .A(n83), .Z(n273) );
  BUF_X1 U2035 ( .A(n81), .Z(n270) );
  BUF_X1 U2036 ( .A(n80), .Z(n264) );
  BUF_X1 U2037 ( .A(n103), .Z(n258) );
  BUF_X1 U2038 ( .A(n102), .Z(n255) );
  BUF_X1 U2039 ( .A(n108), .Z(n249) );
  BUF_X2 U2040 ( .A(n67), .Z(n216) );
  BUF_X1 U2041 ( .A(n69), .Z(n204) );
  BUF_X1 U2042 ( .A(n72), .Z(n201) );
  BUF_X1 U2043 ( .A(n73), .Z(n198) );
  BUF_X1 U2044 ( .A(n75), .Z(n195) );
  BUF_X1 U2045 ( .A(n76), .Z(n192) );
  BUF_X1 U2046 ( .A(n70), .Z(n189) );
  BUF_X1 U2047 ( .A(n74), .Z(n186) );
  BUF_X1 U2048 ( .A(n71), .Z(n183) );
  BUF_X1 U2049 ( .A(n77), .Z(n180) );
  BUF_X1 U2050 ( .A(n75), .Z(n196) );
  BUF_X1 U2051 ( .A(n73), .Z(n199) );
  BUF_X1 U2052 ( .A(n72), .Z(n202) );
  BUF_X1 U2053 ( .A(n91), .Z(n211) );
  BUF_X1 U2054 ( .A(n90), .Z(n208) );
  BUF_X1 U2055 ( .A(n69), .Z(n205) );
  BUF_X1 U2056 ( .A(n76), .Z(n193) );
  BUF_X1 U2057 ( .A(n70), .Z(n190) );
  BUF_X1 U2058 ( .A(n74), .Z(n187) );
  BUF_X1 U2059 ( .A(n71), .Z(n184) );
  BUF_X1 U2060 ( .A(n77), .Z(n181) );
  BUF_X1 U2061 ( .A(n79), .Z(n178) );
  BUF_X1 U2062 ( .A(n78), .Z(n175) );
  BUF_X1 U2063 ( .A(n94), .Z(n172) );
  BUF_X1 U2064 ( .A(n100), .Z(n169) );
  BUF_X1 U2065 ( .A(n99), .Z(n166) );
  BUF_X1 U2066 ( .A(n79), .Z(n177) );
  BUF_X1 U2067 ( .A(n78), .Z(n174) );
  BUF_X1 U2068 ( .A(n89), .Z(n290) );
  BUF_X1 U2069 ( .A(n88), .Z(n287) );
  BUF_X1 U2070 ( .A(n87), .Z(n284) );
  BUF_X1 U2071 ( .A(n94), .Z(n171) );
  NOR2_X1 U2072 ( .A1(n210), .A2(n127), .ZN(\p[6][17] ) );
  NOR2_X1 U2073 ( .A1(n207), .A2(n127), .ZN(\p[6][18] ) );
  NOR2_X1 U2074 ( .A1(n204), .A2(n127), .ZN(\p[6][19] ) );
  NOR2_X1 U2075 ( .A1(n201), .A2(n127), .ZN(\p[6][20] ) );
  NOR2_X1 U2076 ( .A1(n198), .A2(n127), .ZN(\p[6][21] ) );
  NOR2_X1 U2077 ( .A1(n195), .A2(n127), .ZN(\p[6][22] ) );
  NOR2_X1 U2078 ( .A1(n192), .A2(n127), .ZN(\p[6][23] ) );
  NOR2_X1 U2079 ( .A1(n189), .A2(n127), .ZN(\p[6][24] ) );
  NOR2_X1 U2080 ( .A1(n186), .A2(n127), .ZN(\p[6][25] ) );
  NOR2_X1 U2081 ( .A1(n183), .A2(n127), .ZN(\p[6][26] ) );
  NOR2_X1 U2082 ( .A1(n222), .A2(n305), .ZN(\p[8][14] ) );
  NOR2_X1 U2083 ( .A1(n222), .A2(n297), .ZN(\p[11][17] ) );
  NOR2_X1 U2084 ( .A1(n222), .A2(n288), .ZN(\p[14][20] ) );
  NOR2_X1 U2085 ( .A1(n222), .A2(n279), .ZN(\p[17][23] ) );
  NOR2_X1 U2086 ( .A1(n222), .A2(n294), .ZN(\p[12][18] ) );
  NOR2_X1 U2087 ( .A1(n222), .A2(n285), .ZN(\p[15][21] ) );
  NOR2_X1 U2088 ( .A1(n222), .A2(n276), .ZN(\p[18][24] ) );
  NOR2_X1 U2089 ( .A1(n222), .A2(n300), .ZN(\p[10][16] ) );
  NOR2_X1 U2090 ( .A1(n222), .A2(n291), .ZN(\p[13][19] ) );
  NOR2_X1 U2091 ( .A1(n222), .A2(n282), .ZN(\p[16][22] ) );
  NOR2_X1 U2092 ( .A1(n222), .A2(n273), .ZN(\p[19][25] ) );
  NOR2_X1 U2093 ( .A1(n229), .A2(n305), .ZN(\p[8][11] ) );
  NOR2_X1 U2094 ( .A1(n229), .A2(n297), .ZN(\p[11][14] ) );
  NOR2_X1 U2095 ( .A1(n229), .A2(n288), .ZN(\p[14][17] ) );
  NOR2_X1 U2096 ( .A1(n229), .A2(n279), .ZN(\p[17][20] ) );
  NOR2_X1 U2097 ( .A1(n229), .A2(n270), .ZN(\p[20][23] ) );
  NOR2_X1 U2098 ( .A1(n229), .A2(n294), .ZN(\p[12][15] ) );
  NOR2_X1 U2099 ( .A1(n229), .A2(n285), .ZN(\p[15][18] ) );
  NOR2_X1 U2100 ( .A1(n229), .A2(n276), .ZN(\p[18][21] ) );
  NOR2_X1 U2101 ( .A1(n229), .A2(n267), .ZN(\p[21][24] ) );
  NOR2_X1 U2102 ( .A1(n194), .A2(n316), .ZN(\p[0][17] ) );
  NOR2_X1 U2103 ( .A1(n200), .A2(n317), .ZN(\p[0][15] ) );
  NOR2_X1 U2104 ( .A1(n197), .A2(n316), .ZN(\p[0][16] ) );
  NOR2_X1 U2105 ( .A1(n209), .A2(n317), .ZN(\p[0][12] ) );
  NOR2_X1 U2106 ( .A1(n212), .A2(n317), .ZN(\p[0][11] ) );
  NOR2_X1 U2107 ( .A1(n206), .A2(n317), .ZN(\p[0][13] ) );
  NOR2_X1 U2108 ( .A1(n203), .A2(n317), .ZN(\p[0][14] ) );
  NOR2_X1 U2109 ( .A1(n191), .A2(n316), .ZN(\p[0][18] ) );
  NOR2_X1 U2110 ( .A1(n188), .A2(n316), .ZN(\p[0][19] ) );
  NOR2_X1 U2111 ( .A1(n185), .A2(n316), .ZN(\p[0][20] ) );
  NOR2_X1 U2112 ( .A1(n182), .A2(n316), .ZN(\p[0][21] ) );
  NOR2_X1 U2113 ( .A1(n179), .A2(n316), .ZN(\p[0][22] ) );
  NOR2_X1 U2114 ( .A1(n176), .A2(n316), .ZN(\p[0][23] ) );
  NOR2_X1 U2115 ( .A1(n173), .A2(n316), .ZN(\p[0][24] ) );
  NOR2_X1 U2116 ( .A1(n170), .A2(n316), .ZN(\p[0][25] ) );
  NOR2_X1 U2117 ( .A1(n167), .A2(n316), .ZN(\p[0][26] ) );
  NOR2_X1 U2118 ( .A1(n230), .A2(n112), .ZN(\p[10][13] ) );
  NOR2_X1 U2119 ( .A1(n229), .A2(n291), .ZN(\p[13][16] ) );
  NOR2_X1 U2120 ( .A1(n229), .A2(n282), .ZN(\p[16][19] ) );
  NOR2_X1 U2121 ( .A1(n229), .A2(n273), .ZN(\p[19][22] ) );
  NOR2_X1 U2122 ( .A1(n229), .A2(n264), .ZN(\p[22][25] ) );
  NOR2_X1 U2123 ( .A1(n302), .A2(n228), .ZN(\p[9][12] ) );
  NOR2_X1 U2124 ( .A1(n302), .A2(n226), .ZN(\p[9][13] ) );
  NOR2_X1 U2125 ( .A1(n302), .A2(n222), .ZN(\p[9][15] ) );
  NOR2_X1 U2126 ( .A1(n204), .A2(n134), .ZN(\p[3][16] ) );
  NOR2_X1 U2127 ( .A1(n439), .A2(n136), .ZN(\p[3][10] ) );
  NOR2_X1 U2128 ( .A1(n189), .A2(n134), .ZN(\p[3][21] ) );
  NOR2_X1 U2129 ( .A1(n183), .A2(n134), .ZN(\p[3][23] ) );
  NOR2_X1 U2130 ( .A1(n213), .A2(n127), .ZN(\p[6][16] ) );
  NOR2_X1 U2131 ( .A1(n443), .A2(n294), .ZN(\p[12][12] ) );
  NOR2_X1 U2132 ( .A1(n442), .A2(n294), .ZN(\p[12][13] ) );
  NOR2_X1 U2133 ( .A1(n201), .A2(n134), .ZN(\p[3][17] ) );
  NOR2_X1 U2134 ( .A1(n207), .A2(n134), .ZN(\p[3][15] ) );
  NOR2_X1 U2135 ( .A1(n216), .A2(n134), .ZN(\p[3][12] ) );
  NOR2_X1 U2136 ( .A1(n117), .A2(n134), .ZN(\p[3][11] ) );
  NOR2_X1 U2137 ( .A1(n198), .A2(n134), .ZN(\p[3][18] ) );
  NOR2_X1 U2138 ( .A1(n186), .A2(n134), .ZN(\p[3][22] ) );
  NOR2_X1 U2139 ( .A1(n180), .A2(n134), .ZN(\p[3][24] ) );
  NOR2_X1 U2140 ( .A1(n171), .A2(n134), .ZN(\p[3][27] ) );
  NOR2_X1 U2141 ( .A1(n442), .A2(n297), .ZN(\p[11][12] ) );
  NOR2_X1 U2142 ( .A1(n221), .A2(n309), .ZN(\p[5][12] ) );
  NOR2_X1 U2143 ( .A1(n116), .A2(n309), .ZN(\p[5][13] ) );
  NOR2_X1 U2144 ( .A1(n226), .A2(n307), .ZN(\p[7][11] ) );
  NOR2_X1 U2145 ( .A1(n228), .A2(n119), .ZN(\p[7][10] ) );
  NOR2_X1 U2146 ( .A1(n217), .A2(n126), .ZN(\p[6][15] ) );
  NOR2_X1 U2147 ( .A1(n219), .A2(n126), .ZN(\p[6][14] ) );
  NOR2_X1 U2148 ( .A1(n232), .A2(n112), .ZN(\p[10][12] ) );
  NOR2_X1 U2149 ( .A1(n213), .A2(n135), .ZN(\p[3][13] ) );
  NOR2_X1 U2150 ( .A1(n210), .A2(n136), .ZN(\p[3][14] ) );
  NOR2_X1 U2151 ( .A1(n195), .A2(n135), .ZN(\p[3][19] ) );
  NOR2_X1 U2152 ( .A1(n192), .A2(n136), .ZN(\p[3][20] ) );
  NOR2_X1 U2153 ( .A1(n177), .A2(n135), .ZN(\p[3][25] ) );
  NOR2_X1 U2154 ( .A1(n174), .A2(n136), .ZN(\p[3][26] ) );
  NOR2_X1 U2155 ( .A1(n123), .A2(n316), .ZN(\p[0][1] ) );
  NOR2_X1 U2156 ( .A1(n237), .A2(n291), .ZN(\p[13][13] ) );
  NOR2_X1 U2157 ( .A1(n123), .A2(n291), .ZN(\p[13][14] ) );
  NOR2_X1 U2158 ( .A1(n442), .A2(n303), .ZN(\p[8][9] ) );
  NOR2_X1 U2159 ( .A1(n214), .A2(n110), .ZN(\p[1][11] ) );
  NOR2_X1 U2160 ( .A1(n216), .A2(n310), .ZN(\p[4][13] ) );
  NOR2_X1 U2161 ( .A1(n213), .A2(n311), .ZN(\p[4][14] ) );
  NOR2_X1 U2162 ( .A1(n215), .A2(n317), .ZN(\p[0][10] ) );
  NOR2_X1 U2163 ( .A1(n116), .A2(n314), .ZN(\p[2][10] ) );
  NOR2_X1 U2164 ( .A1(n237), .A2(n297), .ZN(\p[11][11] ) );
  NOR2_X1 U2165 ( .A1(n218), .A2(n110), .ZN(\p[1][10] ) );
  NOR2_X1 U2166 ( .A1(n443), .A2(n303), .ZN(\p[8][8] ) );
  AND2_X1 U2167 ( .A1(N189), .A2(n146), .ZN(N253) );
  AND2_X1 U2168 ( .A1(N190), .A2(n146), .ZN(N254) );
  AND2_X1 U2169 ( .A1(N179), .A2(n146), .ZN(N243) );
  AND2_X1 U2170 ( .A1(N180), .A2(n146), .ZN(N244) );
  AND2_X1 U2171 ( .A1(N181), .A2(n146), .ZN(N245) );
  AND2_X1 U2172 ( .A1(N182), .A2(n146), .ZN(N246) );
  AND2_X1 U2173 ( .A1(N183), .A2(n146), .ZN(N247) );
  AND2_X1 U2174 ( .A1(N184), .A2(n146), .ZN(N248) );
  AND2_X1 U2175 ( .A1(N185), .A2(n146), .ZN(N249) );
  AND2_X1 U2176 ( .A1(N186), .A2(n146), .ZN(N250) );
  AND2_X1 U2177 ( .A1(N187), .A2(n146), .ZN(N251) );
  AND2_X1 U2178 ( .A1(N188), .A2(n146), .ZN(N252) );
  AND2_X1 U2179 ( .A1(N193), .A2(n147), .ZN(N257) );
  AND2_X1 U2180 ( .A1(N192), .A2(n147), .ZN(N256) );
  AND2_X1 U2181 ( .A1(N191), .A2(n147), .ZN(N255) );
  BUF_X2 U2182 ( .A(\p[2][63] ), .Z(n414) );
  BUF_X2 U2183 ( .A(\p[5][63] ), .Z(n423) );
  BUF_X2 U2184 ( .A(\p[61][63] ), .Z(n399) );
  BUF_X2 U2185 ( .A(\p[9][63] ), .Z(n322) );
  BUF_X2 U2186 ( .A(\p[61][63] ), .Z(n400) );
  BUF_X2 U2187 ( .A(\p[7][63] ), .Z(n429) );
  BUF_X1 U2188 ( .A(\p[61][63] ), .Z(n401) );
  BUF_X1 U2189 ( .A(n97), .Z(n161) );
  BUF_X1 U2190 ( .A(n96), .Z(n158) );
  BUF_X1 U2191 ( .A(n95), .Z(n155) );
  BUF_X1 U2192 ( .A(n82), .Z(n266) );
  BUF_X1 U2193 ( .A(n81), .Z(n269) );
  BUF_X1 U2194 ( .A(n80), .Z(n263) );
  BUF_X1 U2195 ( .A(n89), .Z(n289) );
  BUF_X1 U2196 ( .A(n104), .Z(n260) );
  BUF_X1 U2197 ( .A(n103), .Z(n257) );
  BUF_X1 U2198 ( .A(n102), .Z(n254) );
  BUF_X1 U2199 ( .A(n88), .Z(n286) );
  BUF_X1 U2200 ( .A(n108), .Z(n248) );
  BUF_X1 U2201 ( .A(n87), .Z(n283) );
  BUF_X1 U2202 ( .A(n101), .Z(n251) );
  BUF_X1 U2203 ( .A(n107), .Z(n245) );
  BUF_X1 U2204 ( .A(n86), .Z(n280) );
  BUF_X1 U2205 ( .A(n105), .Z(n242) );
  BUF_X1 U2206 ( .A(n106), .Z(n239) );
  BUF_X1 U2207 ( .A(n85), .Z(n274) );
  BUF_X1 U2208 ( .A(n84), .Z(n277) );
  BUF_X1 U2209 ( .A(n83), .Z(n271) );
  BUF_X1 U2210 ( .A(n101), .Z(n252) );
  BUF_X1 U2211 ( .A(n107), .Z(n246) );
  BUF_X1 U2212 ( .A(n105), .Z(n243) );
  BUF_X1 U2213 ( .A(n106), .Z(n240) );
  BUF_X1 U2214 ( .A(n98), .Z(n163) );
  BUF_X1 U2215 ( .A(n97), .Z(n160) );
  BUF_X1 U2216 ( .A(n96), .Z(n157) );
  BUF_X1 U2217 ( .A(n95), .Z(n154) );
  BUF_X1 U2218 ( .A(n100), .Z(n168) );
  BUF_X1 U2219 ( .A(n99), .Z(n165) );
  BUF_X1 U2220 ( .A(n98), .Z(n162) );
  BUF_X1 U2221 ( .A(n97), .Z(n159) );
  BUF_X1 U2222 ( .A(n96), .Z(n156) );
  BUF_X1 U2223 ( .A(n95), .Z(n153) );
  NOR2_X1 U2224 ( .A1(n180), .A2(n127), .ZN(\p[6][27] ) );
  NOR2_X1 U2225 ( .A1(n177), .A2(n127), .ZN(\p[6][28] ) );
  NOR2_X1 U2226 ( .A1(n174), .A2(n127), .ZN(\p[6][29] ) );
  NOR2_X1 U2227 ( .A1(n171), .A2(n127), .ZN(\p[6][30] ) );
  NOR2_X1 U2228 ( .A1(n168), .A2(n127), .ZN(\p[6][31] ) );
  NOR2_X1 U2229 ( .A1(n165), .A2(n127), .ZN(\p[6][32] ) );
  NOR2_X1 U2230 ( .A1(n162), .A2(n127), .ZN(\p[6][33] ) );
  NOR2_X1 U2231 ( .A1(n159), .A2(n127), .ZN(\p[6][34] ) );
  NOR2_X1 U2232 ( .A1(n156), .A2(n127), .ZN(\p[6][35] ) );
  NOR2_X1 U2233 ( .A1(n222), .A2(n270), .ZN(\p[20][26] ) );
  NOR2_X1 U2234 ( .A1(n222), .A2(n261), .ZN(\p[23][29] ) );
  NOR2_X1 U2235 ( .A1(n222), .A2(n252), .ZN(\p[26][32] ) );
  NOR2_X1 U2236 ( .A1(n222), .A2(n243), .ZN(\p[29][35] ) );
  NOR2_X1 U2237 ( .A1(n222), .A2(n267), .ZN(\p[21][27] ) );
  NOR2_X1 U2238 ( .A1(n222), .A2(n258), .ZN(\p[24][30] ) );
  NOR2_X1 U2239 ( .A1(n222), .A2(n249), .ZN(\p[27][33] ) );
  NOR2_X1 U2240 ( .A1(n222), .A2(n240), .ZN(\p[30][36] ) );
  NOR2_X1 U2241 ( .A1(n230), .A2(n252), .ZN(\p[26][29] ) );
  NOR2_X1 U2242 ( .A1(n222), .A2(n264), .ZN(\p[22][28] ) );
  NOR2_X1 U2243 ( .A1(n222), .A2(n255), .ZN(\p[25][31] ) );
  NOR2_X1 U2244 ( .A1(n222), .A2(n246), .ZN(\p[28][34] ) );
  NOR2_X1 U2245 ( .A1(n229), .A2(n261), .ZN(\p[23][26] ) );
  NOR2_X1 U2246 ( .A1(n229), .A2(n243), .ZN(\p[29][32] ) );
  NOR2_X1 U2247 ( .A1(n229), .A2(n258), .ZN(\p[24][27] ) );
  NOR2_X1 U2248 ( .A1(n229), .A2(n249), .ZN(\p[27][30] ) );
  NOR2_X1 U2249 ( .A1(n229), .A2(n240), .ZN(\p[30][33] ) );
  NOR2_X1 U2250 ( .A1(n229), .A2(n255), .ZN(\p[25][28] ) );
  NOR2_X1 U2251 ( .A1(n229), .A2(n246), .ZN(\p[28][31] ) );
  NOR2_X1 U2252 ( .A1(n168), .A2(n134), .ZN(\p[3][28] ) );
  NOR2_X1 U2253 ( .A1(n153), .A2(n127), .ZN(\p[6][36] ) );
  NOR2_X1 U2254 ( .A1(n123), .A2(n243), .ZN(\p[29][30] ) );
  AND2_X1 U2255 ( .A1(n432), .A2(A_reg[0]), .ZN(\p[63][63] ) );
  AND2_X1 U2256 ( .A1(n114), .A2(n435), .ZN(\p[0][63] ) );
  AND2_X1 U2257 ( .A1(n432), .A2(A_reg[7]), .ZN(\p[56][63] ) );
  AND2_X1 U2258 ( .A1(n432), .A2(n109), .ZN(\p[60][63] ) );
  AND2_X1 U2259 ( .A1(n432), .A2(A_reg[4]), .ZN(\p[59][63] ) );
  AND2_X1 U2260 ( .A1(n432), .A2(A_reg[6]), .ZN(\p[57][63] ) );
  AND2_X1 U2261 ( .A1(B_reg[3]), .A2(n437), .ZN(\p[3][63] ) );
  AND2_X1 U2262 ( .A1(B_reg[6]), .A2(n437), .ZN(\p[6][63] ) );
  AND2_X1 U2263 ( .A1(n432), .A2(A_reg[1]), .ZN(\p[62][63] ) );
  AND2_X1 U2264 ( .A1(B_reg[1]), .A2(n435), .ZN(\p[1][63] ) );
  AND2_X1 U2265 ( .A1(N167), .A2(n145), .ZN(N231) );
  AND2_X1 U2266 ( .A1(N168), .A2(n145), .ZN(N232) );
  AND2_X1 U2267 ( .A1(N169), .A2(n145), .ZN(N233) );
  AND2_X1 U2268 ( .A1(N170), .A2(n145), .ZN(N234) );
  AND2_X1 U2269 ( .A1(N171), .A2(n145), .ZN(N235) );
  AND2_X1 U2270 ( .A1(N172), .A2(n145), .ZN(N236) );
  AND2_X1 U2271 ( .A1(N173), .A2(n145), .ZN(N237) );
  AND2_X1 U2272 ( .A1(N174), .A2(n145), .ZN(N238) );
  AND2_X1 U2273 ( .A1(N175), .A2(n145), .ZN(N239) );
  AND2_X1 U2274 ( .A1(N176), .A2(n145), .ZN(N240) );
  AND2_X1 U2275 ( .A1(N177), .A2(n145), .ZN(N241) );
  AND2_X1 U2276 ( .A1(N178), .A2(n145), .ZN(N242) );
  BUF_X1 U2277 ( .A(\p[50][63] ), .Z(n371) );
  BUF_X2 U2278 ( .A(\p[11][63] ), .Z(n326) );
  BUF_X2 U2279 ( .A(\p[2][63] ), .Z(n415) );
  BUF_X2 U2280 ( .A(\p[14][63] ), .Z(n332) );
  BUF_X2 U2281 ( .A(\p[5][63] ), .Z(n424) );
  BUF_X2 U2282 ( .A(\p[54][63] ), .Z(n378) );
  BUF_X2 U2283 ( .A(\p[51][63] ), .Z(n372) );
  BUF_X2 U2284 ( .A(\p[53][63] ), .Z(n376) );
  BUF_X2 U2285 ( .A(\p[52][63] ), .Z(n374) );
  BUF_X2 U2286 ( .A(\p[50][63] ), .Z(n370) );
  BUF_X2 U2287 ( .A(\p[49][63] ), .Z(n368) );
  BUF_X2 U2288 ( .A(\p[12][63] ), .Z(n328) );
  BUF_X2 U2289 ( .A(\p[10][63] ), .Z(n324) );
  BUF_X2 U2290 ( .A(\p[13][63] ), .Z(n330) );
  BUF_X2 U2291 ( .A(\p[7][63] ), .Z(n430) );
  BUF_X1 U2292 ( .A(\p[49][63] ), .Z(n369) );
  BUF_X1 U2293 ( .A(\p[51][63] ), .Z(n373) );
  BUF_X1 U2294 ( .A(n81), .Z(n268) );
  BUF_X1 U2295 ( .A(n82), .Z(n265) );
  BUF_X1 U2296 ( .A(n80), .Z(n262) );
  BUF_X1 U2297 ( .A(n104), .Z(n259) );
  BUF_X1 U2298 ( .A(n103), .Z(n256) );
  BUF_X1 U2299 ( .A(n102), .Z(n253) );
  BUF_X1 U2300 ( .A(n108), .Z(n247) );
  BUF_X1 U2301 ( .A(n101), .Z(n250) );
  BUF_X1 U2302 ( .A(n107), .Z(n244) );
  BUF_X1 U2303 ( .A(n105), .Z(n241) );
  BUF_X1 U2304 ( .A(n106), .Z(n238) );
  AND2_X1 U2305 ( .A1(N154), .A2(n143), .ZN(N218) );
  AND2_X1 U2306 ( .A1(N155), .A2(n144), .ZN(N219) );
  AND2_X1 U2307 ( .A1(N156), .A2(n144), .ZN(N220) );
  AND2_X1 U2308 ( .A1(N157), .A2(n144), .ZN(N221) );
  AND2_X1 U2309 ( .A1(N158), .A2(n144), .ZN(N222) );
  AND2_X1 U2310 ( .A1(N159), .A2(n144), .ZN(N223) );
  AND2_X1 U2311 ( .A1(N160), .A2(n144), .ZN(N224) );
  AND2_X1 U2312 ( .A1(N161), .A2(n144), .ZN(N225) );
  AND2_X1 U2313 ( .A1(N162), .A2(n144), .ZN(N226) );
  AND2_X1 U2314 ( .A1(N163), .A2(n144), .ZN(N227) );
  AND2_X1 U2315 ( .A1(N164), .A2(n144), .ZN(N228) );
  AND2_X1 U2316 ( .A1(N165), .A2(n144), .ZN(N229) );
  AND2_X1 U2317 ( .A1(N166), .A2(n144), .ZN(N230) );
  BUF_X1 U2318 ( .A(\p[13][63] ), .Z(n331) );
  BUF_X1 U2319 ( .A(\p[14][63] ), .Z(n333) );
  BUF_X1 U2320 ( .A(\p[2][63] ), .Z(n416) );
  BUF_X1 U2321 ( .A(\p[12][63] ), .Z(n329) );
  BUF_X1 U2322 ( .A(\p[5][63] ), .Z(n425) );
  NOR2_X1 U2323 ( .A1(n236), .A2(n317), .ZN(\p[0][0] ) );
  AND2_X1 U2324 ( .A1(n434), .A2(n437), .ZN(\p[32][63] ) );
  BUF_X1 U2325 ( .A(\p[7][63] ), .Z(n431) );
  AND2_X1 U2326 ( .A1(N133), .A2(n142), .ZN(N197) );
  AND2_X1 U2327 ( .A1(N134), .A2(n142), .ZN(N198) );
  AND2_X1 U2328 ( .A1(N135), .A2(n142), .ZN(N199) );
  AND2_X1 U2329 ( .A1(N142), .A2(n142), .ZN(N206) );
  AND2_X1 U2330 ( .A1(N143), .A2(n143), .ZN(N207) );
  AND2_X1 U2331 ( .A1(N144), .A2(n143), .ZN(N208) );
  AND2_X1 U2332 ( .A1(N145), .A2(n143), .ZN(N209) );
  AND2_X1 U2333 ( .A1(N146), .A2(n143), .ZN(N210) );
  AND2_X1 U2334 ( .A1(N147), .A2(n143), .ZN(N211) );
  AND2_X1 U2335 ( .A1(N148), .A2(n143), .ZN(N212) );
  AND2_X1 U2336 ( .A1(N149), .A2(n143), .ZN(N213) );
  AND2_X1 U2337 ( .A1(N150), .A2(n143), .ZN(N214) );
  AND2_X1 U2338 ( .A1(N151), .A2(n143), .ZN(N215) );
  AND2_X1 U2339 ( .A1(N152), .A2(n143), .ZN(N216) );
  AND2_X1 U2340 ( .A1(N153), .A2(n143), .ZN(N217) );
  AND2_X1 U2341 ( .A1(N136), .A2(n142), .ZN(N200) );
  AND2_X1 U2342 ( .A1(N137), .A2(n142), .ZN(N201) );
  AND2_X1 U2343 ( .A1(N138), .A2(n142), .ZN(N202) );
  AND2_X1 U2344 ( .A1(N139), .A2(n142), .ZN(N203) );
  AND2_X1 U2345 ( .A1(N140), .A2(n142), .ZN(N204) );
  AND2_X1 U2346 ( .A1(N141), .A2(n142), .ZN(N205) );
  BUF_X1 U2347 ( .A(n438), .Z(n150) );
  BUF_X1 U2348 ( .A(n438), .Z(n151) );
  BUF_X1 U2349 ( .A(n438), .Z(n149) );
  AND2_X1 U2350 ( .A1(n111), .A2(n114), .ZN(\p[0][5] ) );
  INV_X1 U2351 ( .A(A_reg[0]), .ZN(n443) );
  NOR2_X1 U2352 ( .A1(n139), .A2(n113), .ZN(\p[4][10] ) );
  NOR2_X1 U2353 ( .A1(n120), .A2(n125), .ZN(\p[6][6] ) );
  NOR2_X1 U2354 ( .A1(n223), .A2(n309), .ZN(\p[5][11] ) );
  NOR2_X1 U2355 ( .A1(n222), .A2(n307), .ZN(\p[7][13] ) );
  NOR2_X1 U2356 ( .A1(n117), .A2(n310), .ZN(\p[4][12] ) );
  NOR2_X1 U2357 ( .A1(n124), .A2(n112), .ZN(\p[10][11] ) );
  NOR2_X1 U2358 ( .A1(n124), .A2(n125), .ZN(\p[6][7] ) );
  NOR2_X1 U2359 ( .A1(n120), .A2(n112), .ZN(\p[10][10] ) );
  NOR2_X1 U2360 ( .A1(n302), .A2(n124), .ZN(\p[9][10] ) );
  AND2_X1 U2361 ( .A1(A_reg[6]), .A2(B_reg[6]), .ZN(\p[6][12] ) );
  AND2_X1 U2362 ( .A1(n109), .A2(B_reg[6]), .ZN(\p[6][9] ) );
  AND2_X1 U2363 ( .A1(A_reg[3]), .A2(B_reg[4]), .ZN(\p[4][7] ) );
  BUF_X1 U2364 ( .A(A_reg[31]), .Z(n435) );
  BUF_X1 U2365 ( .A(B_reg[31]), .Z(n432) );
  BUF_X1 U2366 ( .A(A_reg[31]), .Z(n437) );
  BUF_X1 U2367 ( .A(A_reg[31]), .Z(n436) );
  AND2_X1 U2368 ( .A1(B_reg[2]), .A2(n436), .ZN(\p[2][63] ) );
  AND2_X1 U2369 ( .A1(B_reg[5]), .A2(n437), .ZN(\p[5][63] ) );
  AND2_X1 U2370 ( .A1(B_reg[7]), .A2(n437), .ZN(\p[7][63] ) );
  AND2_X1 U2371 ( .A1(n437), .A2(B_reg[9]), .ZN(\p[9][63] ) );
  BUF_X1 U2372 ( .A(B_reg[31]), .Z(n433) );
  AND2_X1 U2373 ( .A1(n433), .A2(A_reg[12]), .ZN(\p[51][63] ) );
  AND2_X1 U2374 ( .A1(n432), .A2(A_reg[10]), .ZN(\p[53][63] ) );
  AND2_X1 U2375 ( .A1(n432), .A2(A_reg[11]), .ZN(\p[52][63] ) );
  AND2_X1 U2376 ( .A1(B_reg[10]), .A2(n435), .ZN(\p[10][63] ) );
  AND2_X1 U2377 ( .A1(B_reg[11]), .A2(n435), .ZN(\p[11][63] ) );
  AND2_X1 U2378 ( .A1(B_reg[12]), .A2(n435), .ZN(\p[12][63] ) );
  AND2_X1 U2379 ( .A1(B_reg[8]), .A2(n437), .ZN(\p[8][63] ) );
  AND2_X1 U2380 ( .A1(n433), .A2(A_reg[13]), .ZN(\p[50][63] ) );
  AND2_X1 U2381 ( .A1(n433), .A2(A_reg[14]), .ZN(\p[49][63] ) );
  AND2_X1 U2382 ( .A1(B_reg[13]), .A2(n435), .ZN(\p[13][63] ) );
  AND2_X1 U2383 ( .A1(B_reg[14]), .A2(n435), .ZN(\p[14][63] ) );
  AND2_X1 U2384 ( .A1(n433), .A2(A_reg[19]), .ZN(\p[44][63] ) );
  AND2_X1 U2385 ( .A1(n433), .A2(A_reg[18]), .ZN(\p[45][63] ) );
  AND2_X1 U2386 ( .A1(n433), .A2(A_reg[16]), .ZN(\p[47][63] ) );
  AND2_X1 U2387 ( .A1(n433), .A2(A_reg[17]), .ZN(\p[46][63] ) );
  AND2_X1 U2388 ( .A1(n433), .A2(A_reg[20]), .ZN(\p[43][63] ) );
  AND2_X1 U2389 ( .A1(n433), .A2(A_reg[15]), .ZN(\p[48][63] ) );
  AND2_X1 U2390 ( .A1(B_reg[18]), .A2(n435), .ZN(\p[18][63] ) );
  AND2_X1 U2391 ( .A1(B_reg[15]), .A2(n435), .ZN(\p[15][63] ) );
  AND2_X1 U2392 ( .A1(B_reg[16]), .A2(n435), .ZN(\p[16][63] ) );
  AND2_X1 U2393 ( .A1(B_reg[17]), .A2(n435), .ZN(\p[17][63] ) );
  AND2_X1 U2394 ( .A1(B_reg[19]), .A2(n435), .ZN(\p[19][63] ) );
  AND2_X1 U2395 ( .A1(n434), .A2(A_reg[25]), .ZN(\p[38][63] ) );
  AND2_X1 U2396 ( .A1(B_reg[25]), .A2(n436), .ZN(\p[25][63] ) );
  AND2_X1 U2397 ( .A1(B_reg[26]), .A2(n436), .ZN(\p[26][63] ) );
  AND2_X1 U2398 ( .A1(n434), .A2(A_reg[26]), .ZN(\p[37][63] ) );
  AND2_X1 U2399 ( .A1(B_reg[27]), .A2(n436), .ZN(\p[27][63] ) );
  AND2_X1 U2400 ( .A1(n434), .A2(A_reg[27]), .ZN(\p[36][63] ) );
  AND2_X1 U2401 ( .A1(n434), .A2(A_reg[28]), .ZN(\p[35][63] ) );
  AND2_X1 U2402 ( .A1(B_reg[28]), .A2(n436), .ZN(\p[28][63] ) );
  AND2_X1 U2403 ( .A1(B_reg[24]), .A2(n436), .ZN(\p[24][63] ) );
  AND2_X1 U2404 ( .A1(n434), .A2(A_reg[24]), .ZN(\p[39][63] ) );
  AND2_X1 U2405 ( .A1(B_reg[29]), .A2(n436), .ZN(\p[29][63] ) );
  AND2_X1 U2406 ( .A1(n434), .A2(A_reg[29]), .ZN(\p[34][63] ) );
  BUF_X1 U2407 ( .A(B_reg[31]), .Z(n434) );
  AND2_X1 U2408 ( .A1(B_reg[30]), .A2(n436), .ZN(\p[30][63] ) );
  AND2_X1 U2409 ( .A1(n434), .A2(A_reg[30]), .ZN(\p[33][63] ) );
  AND2_X1 U2410 ( .A1(B_reg[20]), .A2(n436), .ZN(\p[20][63] ) );
  AND2_X1 U2411 ( .A1(N131), .A2(n142), .ZN(N195) );
  INV_X1 U2412 ( .A(rst), .ZN(n438) );
  AND2_X1 U2413 ( .A1(A[8]), .A2(n148), .ZN(N43) );
  AND2_X1 U2414 ( .A1(A[9]), .A2(n148), .ZN(N44) );
  AND2_X1 U2415 ( .A1(A[10]), .A2(n148), .ZN(N45) );
  AND2_X1 U2416 ( .A1(A[11]), .A2(n148), .ZN(N46) );
  AND2_X1 U2417 ( .A1(A[12]), .A2(n148), .ZN(N47) );
  AND2_X1 U2418 ( .A1(A[13]), .A2(n148), .ZN(N48) );
  AND2_X1 U2419 ( .A1(A[14]), .A2(n148), .ZN(N49) );
  AND2_X1 U2420 ( .A1(A[15]), .A2(n148), .ZN(N50) );
  AND2_X1 U2421 ( .A1(A[16]), .A2(n148), .ZN(N51) );
  AND2_X1 U2422 ( .A1(A[17]), .A2(n148), .ZN(N52) );
  AND2_X1 U2423 ( .A1(A[18]), .A2(n148), .ZN(N53) );
  AND2_X1 U2424 ( .A1(A[19]), .A2(n148), .ZN(N54) );
  AND2_X1 U2425 ( .A1(A[0]), .A2(n147), .ZN(N35) );
  AND2_X1 U2426 ( .A1(A[1]), .A2(n147), .ZN(N36) );
  AND2_X1 U2427 ( .A1(A[2]), .A2(n147), .ZN(N37) );
  AND2_X1 U2428 ( .A1(A[3]), .A2(n147), .ZN(N38) );
  AND2_X1 U2429 ( .A1(A[4]), .A2(n147), .ZN(N39) );
  AND2_X1 U2430 ( .A1(A[5]), .A2(n147), .ZN(N40) );
  AND2_X1 U2431 ( .A1(A[6]), .A2(n147), .ZN(N41) );
  AND2_X1 U2432 ( .A1(A[7]), .A2(n147), .ZN(N42) );
  AND2_X1 U2433 ( .A1(B[24]), .A2(n152), .ZN(N91) );
  AND2_X1 U2434 ( .A1(B[25]), .A2(n152), .ZN(N92) );
  AND2_X1 U2435 ( .A1(B[26]), .A2(n152), .ZN(N93) );
  AND2_X1 U2436 ( .A1(B[27]), .A2(n152), .ZN(N94) );
  AND2_X1 U2437 ( .A1(B[28]), .A2(n152), .ZN(N95) );
  AND2_X1 U2438 ( .A1(B[29]), .A2(n152), .ZN(N96) );
  AND2_X1 U2439 ( .A1(B[30]), .A2(n152), .ZN(N97) );
  AND2_X1 U2440 ( .A1(B[31]), .A2(n152), .ZN(N98) );
  AND2_X1 U2441 ( .A1(B[0]), .A2(n150), .ZN(N67) );
  AND2_X1 U2442 ( .A1(B[1]), .A2(n150), .ZN(N68) );
  AND2_X1 U2443 ( .A1(B[2]), .A2(n150), .ZN(N69) );
  AND2_X1 U2444 ( .A1(B[3]), .A2(n150), .ZN(N70) );
  AND2_X1 U2445 ( .A1(B[4]), .A2(n150), .ZN(N71) );
  AND2_X1 U2446 ( .A1(B[5]), .A2(n150), .ZN(N72) );
  AND2_X1 U2447 ( .A1(B[6]), .A2(n150), .ZN(N73) );
  AND2_X1 U2448 ( .A1(B[7]), .A2(n150), .ZN(N74) );
  AND2_X1 U2449 ( .A1(B[8]), .A2(n150), .ZN(N75) );
  AND2_X1 U2450 ( .A1(B[9]), .A2(n150), .ZN(N76) );
  AND2_X1 U2451 ( .A1(B[10]), .A2(n150), .ZN(N77) );
  AND2_X1 U2452 ( .A1(B[11]), .A2(n150), .ZN(N78) );
  AND2_X1 U2453 ( .A1(B[12]), .A2(n151), .ZN(N79) );
  AND2_X1 U2454 ( .A1(B[13]), .A2(n151), .ZN(N80) );
  AND2_X1 U2455 ( .A1(B[14]), .A2(n151), .ZN(N81) );
  AND2_X1 U2456 ( .A1(B[15]), .A2(n151), .ZN(N82) );
  AND2_X1 U2457 ( .A1(B[16]), .A2(n151), .ZN(N83) );
  AND2_X1 U2458 ( .A1(B[17]), .A2(n151), .ZN(N84) );
  AND2_X1 U2459 ( .A1(B[18]), .A2(n151), .ZN(N85) );
  AND2_X1 U2460 ( .A1(B[19]), .A2(n151), .ZN(N86) );
  AND2_X1 U2461 ( .A1(B[20]), .A2(n151), .ZN(N87) );
  AND2_X1 U2462 ( .A1(B[21]), .A2(n151), .ZN(N88) );
  AND2_X1 U2463 ( .A1(B[22]), .A2(n151), .ZN(N89) );
  AND2_X1 U2464 ( .A1(B[23]), .A2(n151), .ZN(N90) );
  AND2_X1 U2465 ( .A1(A[20]), .A2(n149), .ZN(N55) );
  AND2_X1 U2466 ( .A1(A[21]), .A2(n149), .ZN(N56) );
  AND2_X1 U2467 ( .A1(A[22]), .A2(n149), .ZN(N57) );
  AND2_X1 U2468 ( .A1(A[23]), .A2(n149), .ZN(N58) );
  AND2_X1 U2469 ( .A1(A[24]), .A2(n149), .ZN(N59) );
  AND2_X1 U2470 ( .A1(A[25]), .A2(n149), .ZN(N60) );
  AND2_X1 U2471 ( .A1(A[26]), .A2(n149), .ZN(N61) );
  AND2_X1 U2472 ( .A1(A[27]), .A2(n149), .ZN(N62) );
  AND2_X1 U2473 ( .A1(A[28]), .A2(n149), .ZN(N63) );
  AND2_X1 U2474 ( .A1(A[29]), .A2(n149), .ZN(N64) );
  AND2_X1 U2475 ( .A1(A[30]), .A2(n149), .ZN(N65) );
  AND2_X1 U2476 ( .A1(A[31]), .A2(n149), .ZN(N66) );
  NOR2_X1 U2477 ( .A1(n439), .A2(n113), .ZN(\p[4][11] ) );
  INV_X1 U2478 ( .A(A_reg[7]), .ZN(n439) );
  CLKBUF_X1 U2479 ( .A(n117), .Z(n116) );
  CLKBUF_X1 U2480 ( .A(n125), .Z(n126) );
  INV_X1 U2481 ( .A(A_reg[4]), .ZN(n440) );
  NOR2_X1 U2482 ( .A1(n120), .A2(n115), .ZN(\p[9][9] ) );
  AND2_X1 U2483 ( .A1(n432), .A2(A_reg[9]), .ZN(\p[54][63] ) );
  NOR2_X1 U2484 ( .A1(n216), .A2(n284), .ZN(\p[15][24] ) );
  NOR2_X1 U2485 ( .A1(n217), .A2(n287), .ZN(\p[14][23] ) );
  NOR2_X1 U2486 ( .A1(n216), .A2(n290), .ZN(\p[13][22] ) );
  NOR2_X1 U2487 ( .A1(n216), .A2(n296), .ZN(\p[11][20] ) );
  NOR2_X1 U2488 ( .A1(n216), .A2(n293), .ZN(\p[12][21] ) );
  NOR2_X1 U2489 ( .A1(n217), .A2(n299), .ZN(\p[10][19] ) );
  CLKBUF_X1 U2490 ( .A(n118), .Z(n312) );
  CLKBUF_X1 U2491 ( .A(n119), .Z(n306) );
  AND2_X1 U2492 ( .A1(n111), .A2(B_reg[2]), .ZN(\p[2][7] ) );
  CLKBUF_X1 U2493 ( .A(n443), .Z(n237) );
  CLKBUF_X1 U2494 ( .A(n443), .Z(n235) );
  CLKBUF_X1 U2495 ( .A(n441), .Z(n231) );
  CLKBUF_X1 U2496 ( .A(n441), .Z(n233) );
  CLKBUF_X1 U2497 ( .A(n442), .Z(n123) );
  NOR2_X1 U2498 ( .A1(n439), .A2(n118), .ZN(\p[2][9] ) );
  NOR2_X1 U2499 ( .A1(n139), .A2(n118), .ZN(\p[2][8] ) );
  NOR2_X1 U2500 ( .A1(n440), .A2(n118), .ZN(\p[2][6] ) );
  NOR2_X1 U2501 ( .A1(n140), .A2(n118), .ZN(\p[2][5] ) );
  NOR2_X1 U2502 ( .A1(n442), .A2(n118), .ZN(\p[2][3] ) );
  NOR2_X1 U2503 ( .A1(n153), .A2(n312), .ZN(\p[2][32] ) );
  NOR2_X1 U2504 ( .A1(n156), .A2(n312), .ZN(\p[2][31] ) );
  NOR2_X1 U2505 ( .A1(n159), .A2(n312), .ZN(\p[2][30] ) );
  NOR2_X1 U2506 ( .A1(n235), .A2(n118), .ZN(\p[2][2] ) );
  NOR2_X1 U2507 ( .A1(n162), .A2(n312), .ZN(\p[2][29] ) );
  NOR2_X1 U2508 ( .A1(n137), .A2(n122), .ZN(\p[5][9] ) );
  NOR2_X1 U2509 ( .A1(n140), .A2(n122), .ZN(\p[5][8] ) );
  NOR2_X1 U2510 ( .A1(n124), .A2(n122), .ZN(\p[5][6] ) );
  NOR2_X1 U2511 ( .A1(n443), .A2(n122), .ZN(\p[5][5] ) );
  NOR2_X1 U2512 ( .A1(n153), .A2(n308), .ZN(\p[5][35] ) );
  NOR2_X1 U2513 ( .A1(n156), .A2(n308), .ZN(\p[5][34] ) );
  NOR2_X1 U2514 ( .A1(n159), .A2(n308), .ZN(\p[5][33] ) );
  NOR2_X1 U2515 ( .A1(n162), .A2(n308), .ZN(\p[5][32] ) );
  NOR2_X1 U2516 ( .A1(n165), .A2(n308), .ZN(\p[5][31] ) );
  NOR2_X1 U2517 ( .A1(n168), .A2(n308), .ZN(\p[5][30] ) );
  NOR2_X1 U2518 ( .A1(n171), .A2(n308), .ZN(\p[5][29] ) );
  NOR2_X1 U2519 ( .A1(n153), .A2(n307), .ZN(\p[7][37] ) );
  NOR2_X1 U2520 ( .A1(n156), .A2(n307), .ZN(\p[7][36] ) );
  NOR2_X1 U2521 ( .A1(n159), .A2(n306), .ZN(\p[7][35] ) );
  NOR2_X1 U2522 ( .A1(n162), .A2(n307), .ZN(\p[7][34] ) );
  NOR2_X1 U2523 ( .A1(n165), .A2(n306), .ZN(\p[7][33] ) );
  NOR2_X1 U2524 ( .A1(n168), .A2(n307), .ZN(\p[7][32] ) );
  NOR2_X1 U2525 ( .A1(n171), .A2(n307), .ZN(\p[7][31] ) );
  NOR2_X1 U2526 ( .A1(n174), .A2(n307), .ZN(\p[7][30] ) );
  NOR2_X1 U2527 ( .A1(n177), .A2(n307), .ZN(\p[7][29] ) );
  NOR2_X1 U2528 ( .A1(n124), .A2(n119), .ZN(\p[7][8] ) );
  NOR2_X1 U2529 ( .A1(n120), .A2(n119), .ZN(\p[7][7] ) );
  NOR2_X1 U2530 ( .A1(n441), .A2(n252), .ZN(\p[26][28] ) );
  NOR2_X1 U2531 ( .A1(n441), .A2(n255), .ZN(\p[25][27] ) );
  NOR2_X1 U2532 ( .A1(n232), .A2(n258), .ZN(\p[24][26] ) );
  NOR2_X1 U2533 ( .A1(n231), .A2(n264), .ZN(\p[22][24] ) );
  NOR2_X1 U2534 ( .A1(n232), .A2(n270), .ZN(\p[20][22] ) );
  NOR2_X1 U2535 ( .A1(n232), .A2(n273), .ZN(\p[19][21] ) );
  NOR2_X1 U2536 ( .A1(n231), .A2(n279), .ZN(\p[17][19] ) );
  NOR2_X1 U2537 ( .A1(n232), .A2(n282), .ZN(\p[16][18] ) );
  NOR2_X1 U2538 ( .A1(n231), .A2(n285), .ZN(\p[15][17] ) );
  NOR2_X1 U2539 ( .A1(n232), .A2(n288), .ZN(\p[14][16] ) );
  NOR2_X1 U2540 ( .A1(n232), .A2(n291), .ZN(\p[13][15] ) );
  NOR2_X1 U2541 ( .A1(n232), .A2(n297), .ZN(\p[11][13] ) );
  AND2_X1 U2542 ( .A1(A_reg[8]), .A2(B_reg[0]), .ZN(\p[0][8] ) );
  INV_X1 U2543 ( .A(n224), .ZN(n129) );
  CLKBUF_X1 U2544 ( .A(n128), .Z(n224) );
  NOR2_X1 U2545 ( .A1(n441), .A2(n243), .ZN(\p[29][31] ) );
  NOR2_X1 U2546 ( .A1(n441), .A2(n240), .ZN(\p[30][32] ) );
  AND2_X1 U2547 ( .A1(n432), .A2(A_reg[2]), .ZN(\p[61][63] ) );
  NOR2_X1 U2548 ( .A1(n441), .A2(n246), .ZN(\p[28][30] ) );
  NOR2_X1 U2549 ( .A1(n231), .A2(n249), .ZN(\p[27][29] ) );
  NOR2_X1 U2550 ( .A1(n232), .A2(n305), .ZN(\p[8][10] ) );
  NOR2_X1 U2551 ( .A1(n233), .A2(n118), .ZN(\p[2][4] ) );
  NOR2_X1 U2552 ( .A1(n441), .A2(n119), .ZN(\p[7][9] ) );
  NOR2_X1 U2553 ( .A1(n302), .A2(n233), .ZN(\p[9][11] ) );
  NOR2_X1 U2554 ( .A1(n121), .A2(n122), .ZN(\p[5][7] ) );
  NOR2_X1 U2555 ( .A1(n121), .A2(n125), .ZN(\p[6][8] ) );
  AND2_X1 U2556 ( .A1(n432), .A2(n129), .ZN(\p[58][63] ) );
  NOR2_X1 U2557 ( .A1(n225), .A2(n252), .ZN(\p[26][31] ) );
  NOR2_X1 U2558 ( .A1(n225), .A2(n255), .ZN(\p[25][30] ) );
  NOR2_X1 U2559 ( .A1(n225), .A2(n258), .ZN(\p[24][29] ) );
  NOR2_X1 U2560 ( .A1(n225), .A2(n261), .ZN(\p[23][28] ) );
  NOR2_X1 U2561 ( .A1(n225), .A2(n264), .ZN(\p[22][27] ) );
  NOR2_X1 U2562 ( .A1(n225), .A2(n270), .ZN(\p[20][25] ) );
  NOR2_X1 U2563 ( .A1(n225), .A2(n267), .ZN(\p[21][26] ) );
  NOR2_X1 U2564 ( .A1(n225), .A2(n273), .ZN(\p[19][24] ) );
  NOR2_X1 U2565 ( .A1(n225), .A2(n279), .ZN(\p[17][22] ) );
  NOR2_X1 U2566 ( .A1(n225), .A2(n276), .ZN(\p[18][23] ) );
  NOR2_X1 U2567 ( .A1(n225), .A2(n282), .ZN(\p[16][21] ) );
  CLKBUF_X1 U2568 ( .A(n444), .Z(n310) );
  BUF_X2 U2569 ( .A(n133), .Z(n134) );
  BUF_X1 U2570 ( .A(n133), .Z(n135) );
  INV_X1 U2571 ( .A(B_reg[1]), .ZN(n445) );
  NOR2_X1 U2572 ( .A1(n225), .A2(n243), .ZN(\p[29][34] ) );
  NOR2_X1 U2573 ( .A1(n225), .A2(n240), .ZN(\p[30][35] ) );
  NOR2_X1 U2574 ( .A1(n225), .A2(n246), .ZN(\p[28][33] ) );
  NOR2_X1 U2575 ( .A1(n225), .A2(n249), .ZN(\p[27][32] ) );
  NOR2_X1 U2576 ( .A1(n225), .A2(n305), .ZN(\p[8][13] ) );
  NOR2_X1 U2577 ( .A1(n302), .A2(n224), .ZN(\p[9][14] ) );
  NOR2_X1 U2578 ( .A1(n224), .A2(n306), .ZN(\p[7][12] ) );
  NOR2_X1 U2579 ( .A1(n128), .A2(n309), .ZN(\p[5][10] ) );
  NOR2_X1 U2580 ( .A1(n128), .A2(n126), .ZN(\p[6][11] ) );
  AND2_X1 U2581 ( .A1(B_reg[4]), .A2(n437), .ZN(\p[4][63] ) );
  INV_X1 U2582 ( .A(B_reg[4]), .ZN(n444) );
  AND2_X1 U2583 ( .A1(A_reg[6]), .A2(B_reg[1]), .ZN(\p[1][7] ) );
  AND2_X1 U2584 ( .A1(B_reg[3]), .A2(A_reg[4]), .ZN(\p[3][7] ) );
  AND2_X1 U2585 ( .A1(n432), .A2(A_reg[8]), .ZN(\p[55][63] ) );
  NOR2_X1 U2586 ( .A1(n219), .A2(n284), .ZN(\p[15][23] ) );
  NOR2_X1 U2587 ( .A1(n219), .A2(n287), .ZN(\p[14][22] ) );
  NOR2_X1 U2588 ( .A1(n219), .A2(n290), .ZN(\p[13][21] ) );
  NOR2_X1 U2589 ( .A1(n219), .A2(n296), .ZN(\p[11][19] ) );
  NOR2_X1 U2590 ( .A1(n219), .A2(n293), .ZN(\p[12][20] ) );
  NOR2_X1 U2591 ( .A1(n219), .A2(n299), .ZN(\p[10][18] ) );
  CLKBUF_X1 U2592 ( .A(n440), .Z(n137) );
  CLKBUF_X1 U2593 ( .A(n139), .Z(n223) );
  CLKBUF_X1 U2594 ( .A(n140), .Z(n230) );
  CLKBUF_X1 U2595 ( .A(n140), .Z(n228) );
  CLKBUF_X1 U2596 ( .A(n439), .Z(n221) );
  NOR2_X1 U2597 ( .A1(n218), .A2(n132), .ZN(\p[0][9] ) );
  NOR2_X1 U2598 ( .A1(n440), .A2(n132), .ZN(\p[0][4] ) );
  NOR2_X1 U2599 ( .A1(n140), .A2(n132), .ZN(\p[0][3] ) );
  NOR2_X1 U2600 ( .A1(n155), .A2(n316), .ZN(\p[0][30] ) );
  NOR2_X1 U2601 ( .A1(n231), .A2(n316), .ZN(\p[0][2] ) );
  NOR2_X1 U2602 ( .A1(n158), .A2(n316), .ZN(\p[0][29] ) );
  NOR2_X1 U2603 ( .A1(n161), .A2(n316), .ZN(\p[0][28] ) );
  NOR2_X1 U2604 ( .A1(n164), .A2(n316), .ZN(\p[0][27] ) );
  NOR2_X1 U2605 ( .A1(n154), .A2(n315), .ZN(\p[1][31] ) );
  NOR2_X1 U2606 ( .A1(n157), .A2(n315), .ZN(\p[1][30] ) );
  NOR2_X1 U2607 ( .A1(n160), .A2(n315), .ZN(\p[1][29] ) );
  NOR2_X1 U2608 ( .A1(n163), .A2(n315), .ZN(\p[1][28] ) );
  NOR2_X1 U2609 ( .A1(n442), .A2(n315), .ZN(\p[1][2] ) );
  NOR2_X1 U2610 ( .A1(n441), .A2(n110), .ZN(\p[1][3] ) );
  NOR2_X1 U2611 ( .A1(n138), .A2(n445), .ZN(\p[1][5] ) );
  NOR2_X1 U2612 ( .A1(n117), .A2(n131), .ZN(\p[1][9] ) );
  NOR2_X1 U2613 ( .A1(n140), .A2(n131), .ZN(\p[1][4] ) );
  NOR2_X1 U2614 ( .A1(n131), .A2(n141), .ZN(\p[1][8] ) );
  NOR2_X1 U2615 ( .A1(n128), .A2(n131), .ZN(\p[1][6] ) );
  NOR2_X1 U2616 ( .A1(n153), .A2(n134), .ZN(\p[3][33] ) );
  NOR2_X1 U2617 ( .A1(n156), .A2(n134), .ZN(\p[3][32] ) );
  NOR2_X1 U2618 ( .A1(n159), .A2(n136), .ZN(\p[3][31] ) );
  NOR2_X1 U2619 ( .A1(n162), .A2(n135), .ZN(\p[3][30] ) );
  NOR2_X1 U2620 ( .A1(n165), .A2(n134), .ZN(\p[3][29] ) );
  NOR2_X1 U2621 ( .A1(n120), .A2(n134), .ZN(\p[3][3] ) );
  NOR2_X1 U2622 ( .A1(n121), .A2(n133), .ZN(\p[3][5] ) );
  NOR2_X1 U2623 ( .A1(n139), .A2(n135), .ZN(\p[3][9] ) );
  NOR2_X1 U2624 ( .A1(n124), .A2(n136), .ZN(\p[3][4] ) );
  NOR2_X1 U2625 ( .A1(n153), .A2(n311), .ZN(\p[4][34] ) );
  NOR2_X1 U2626 ( .A1(n156), .A2(n311), .ZN(\p[4][33] ) );
  NOR2_X1 U2627 ( .A1(n159), .A2(n311), .ZN(\p[4][32] ) );
  NOR2_X1 U2628 ( .A1(n162), .A2(n311), .ZN(\p[4][31] ) );
  NOR2_X1 U2629 ( .A1(n165), .A2(n311), .ZN(\p[4][30] ) );
  NOR2_X1 U2630 ( .A1(n168), .A2(n311), .ZN(\p[4][29] ) );
  NOR2_X1 U2631 ( .A1(n124), .A2(n444), .ZN(\p[4][5] ) );
  NOR2_X1 U2632 ( .A1(n128), .A2(n113), .ZN(\p[4][9] ) );
  NOR2_X1 U2633 ( .A1(n120), .A2(n113), .ZN(\p[4][4] ) );
  NOR2_X1 U2634 ( .A1(n138), .A2(n130), .ZN(\p[4][8] ) );
  NOR2_X1 U2635 ( .A1(n121), .A2(n130), .ZN(\p[4][6] ) );
  AND2_X1 U2636 ( .A1(N194), .A2(n147), .ZN(N258) );
  BUF_X4 U2637 ( .A(n117), .Z(n219) );
  BUF_X4 U2638 ( .A(n439), .Z(n220) );
  BUF_X1 U2639 ( .A(n438), .Z(n142) );
  BUF_X1 U2640 ( .A(n438), .Z(n143) );
  BUF_X1 U2641 ( .A(n438), .Z(n144) );
  BUF_X1 U2642 ( .A(n438), .Z(n145) );
  BUF_X1 U2643 ( .A(n438), .Z(n146) );
  BUF_X1 U2644 ( .A(n438), .Z(n147) );
  BUF_X1 U2645 ( .A(n438), .Z(n148) );
  BUF_X1 U2646 ( .A(n438), .Z(n152) );
  BUF_X1 U2647 ( .A(\p[8][63] ), .Z(n318) );
  BUF_X1 U2648 ( .A(\p[8][63] ), .Z(n319) );
  BUF_X1 U2649 ( .A(\p[8][63] ), .Z(n320) );
  BUF_X1 U2650 ( .A(\p[8][63] ), .Z(n321) );
  BUF_X1 U2651 ( .A(\p[15][63] ), .Z(n334) );
  BUF_X1 U2652 ( .A(\p[15][63] ), .Z(n335) );
  BUF_X1 U2653 ( .A(\p[15][63] ), .Z(n336) );
  BUF_X1 U2654 ( .A(\p[16][63] ), .Z(n337) );
  BUF_X1 U2655 ( .A(\p[16][63] ), .Z(n338) );
  BUF_X1 U2656 ( .A(\p[16][63] ), .Z(n339) );
  BUF_X1 U2657 ( .A(\p[17][63] ), .Z(n340) );
  BUF_X1 U2658 ( .A(\p[17][63] ), .Z(n341) );
  BUF_X1 U2659 ( .A(\p[17][63] ), .Z(n342) );
  BUF_X1 U2660 ( .A(\p[18][63] ), .Z(n343) );
  BUF_X1 U2661 ( .A(\p[18][63] ), .Z(n344) );
  BUF_X1 U2662 ( .A(\p[18][63] ), .Z(n345) );
  BUF_X1 U2663 ( .A(\p[19][63] ), .Z(n346) );
  BUF_X1 U2664 ( .A(\p[19][63] ), .Z(n347) );
  BUF_X1 U2665 ( .A(\p[19][63] ), .Z(n348) );
  BUF_X1 U2666 ( .A(\p[20][63] ), .Z(n349) );
  BUF_X1 U2667 ( .A(\p[20][63] ), .Z(n350) );
  BUF_X1 U2668 ( .A(\p[43][63] ), .Z(n351) );
  BUF_X1 U2669 ( .A(\p[43][63] ), .Z(n352) );
  BUF_X1 U2670 ( .A(\p[44][63] ), .Z(n353) );
  BUF_X1 U2671 ( .A(\p[44][63] ), .Z(n354) );
  BUF_X1 U2672 ( .A(\p[44][63] ), .Z(n355) );
  BUF_X1 U2673 ( .A(\p[45][63] ), .Z(n356) );
  BUF_X1 U2674 ( .A(\p[45][63] ), .Z(n357) );
  BUF_X1 U2675 ( .A(\p[45][63] ), .Z(n358) );
  BUF_X1 U2676 ( .A(\p[46][63] ), .Z(n359) );
  BUF_X1 U2677 ( .A(\p[46][63] ), .Z(n360) );
  BUF_X1 U2678 ( .A(\p[46][63] ), .Z(n361) );
  BUF_X1 U2679 ( .A(\p[47][63] ), .Z(n362) );
  BUF_X1 U2680 ( .A(\p[47][63] ), .Z(n363) );
  BUF_X1 U2681 ( .A(\p[47][63] ), .Z(n364) );
  BUF_X1 U2682 ( .A(\p[48][63] ), .Z(n365) );
  BUF_X1 U2683 ( .A(\p[48][63] ), .Z(n366) );
  BUF_X1 U2684 ( .A(\p[48][63] ), .Z(n367) );
  BUF_X1 U2685 ( .A(\p[55][63] ), .Z(n380) );
  BUF_X1 U2686 ( .A(\p[55][63] ), .Z(n381) );
  BUF_X1 U2687 ( .A(\p[55][63] ), .Z(n382) );
  BUF_X1 U2688 ( .A(\p[55][63] ), .Z(n383) );
endmodule

