
module SeqMult_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [0:0] B;
  output [32:0] PRODUCT;
  input TC;
  wire   n1, n2, n3, n4, n5;

  AND2X1 U2 ( .IN1(A[12]), .IN2(n5), .Q(PRODUCT[12]) );
  AND2X1 U3 ( .IN1(A[28]), .IN2(n2), .Q(PRODUCT[28]) );
  AND2X1 U4 ( .IN1(n3), .IN2(A[11]), .Q(PRODUCT[11]) );
  AND2X1 U5 ( .IN1(n5), .IN2(A[7]), .Q(PRODUCT[7]) );
  AND2X1 U6 ( .IN1(A[8]), .IN2(n5), .Q(PRODUCT[8]) );
  AND2X1 U7 ( .IN1(n3), .IN2(A[16]), .Q(PRODUCT[16]) );
  AND2X1 U8 ( .IN1(A[18]), .IN2(n3), .Q(PRODUCT[18]) );
  AND2X1 U9 ( .IN1(A[29]), .IN2(n2), .Q(PRODUCT[29]) );
  AND2X1 U10 ( .IN1(A[30]), .IN2(n3), .Q(PRODUCT[30]) );
  AND2X1 U11 ( .IN1(A[31]), .IN2(n2), .Q(PRODUCT[31]) );
  AND2X1 U12 ( .IN1(A[22]), .IN2(n3), .Q(PRODUCT[22]) );
  AND2X1 U13 ( .IN1(A[20]), .IN2(n2), .Q(PRODUCT[20]) );
  AND2X1 U14 ( .IN1(A[15]), .IN2(n3), .Q(PRODUCT[15]) );
  AND2X1 U15 ( .IN1(A[23]), .IN2(n2), .Q(PRODUCT[23]) );
  AND2X1 U16 ( .IN1(A[27]), .IN2(n5), .Q(PRODUCT[27]) );
  AND2X1 U17 ( .IN1(A[19]), .IN2(n5), .Q(PRODUCT[19]) );
  AND2X1 U18 ( .IN1(n3), .IN2(A[5]), .Q(PRODUCT[5]) );
  AND2X1 U19 ( .IN1(n5), .IN2(A[13]), .Q(PRODUCT[13]) );
  AND2X1 U20 ( .IN1(n3), .IN2(A[9]), .Q(PRODUCT[9]) );
  AND2X1 U21 ( .IN1(n4), .IN2(A[4]), .Q(PRODUCT[4]) );
  AND2X1 U22 ( .IN1(A[24]), .IN2(n2), .Q(PRODUCT[24]) );
  AND2X1 U23 ( .IN1(A[25]), .IN2(n2), .Q(PRODUCT[25]) );
  INVX0 U24 ( .INP(n5), .ZN(n1) );
  INVX0 U25 ( .INP(n1), .ZN(n2) );
  NBUFFX2 U26 ( .INP(B[0]), .Z(n4) );
  AND2X1 U27 ( .IN1(A[14]), .IN2(n3), .Q(PRODUCT[14]) );
  AND2X1 U28 ( .IN1(n4), .IN2(A[6]), .Q(PRODUCT[6]) );
  AND2X1 U29 ( .IN1(n4), .IN2(A[1]), .Q(PRODUCT[1]) );
  AND2X1 U30 ( .IN1(A[3]), .IN2(n4), .Q(PRODUCT[3]) );
  AND2X1 U31 ( .IN1(A[17]), .IN2(n3), .Q(PRODUCT[17]) );
  AND2X1 U32 ( .IN1(A[0]), .IN2(n5), .Q(PRODUCT[0]) );
  NBUFFX2 U33 ( .INP(B[0]), .Z(n3) );
  NBUFFX2 U34 ( .INP(B[0]), .Z(n5) );
  AND2X1 U35 ( .IN1(n4), .IN2(A[2]), .Q(PRODUCT[2]) );
  AND2X1 U36 ( .IN1(A[10]), .IN2(n5), .Q(PRODUCT[10]) );
  AND2X1 U37 ( .IN1(A[21]), .IN2(n2), .Q(PRODUCT[21]) );
  AND2X1 U38 ( .IN1(A[26]), .IN2(n2), .Q(PRODUCT[26]) );
endmodule


module SeqMult_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  INVX0 U3 ( .INP(B[28]), .ZN(n49) );
  XNOR2X1 U4 ( .IN1(n45), .IN2(\B[0] ), .Q(DIFF[1]) );
  AND2X1 U5 ( .IN1(n43), .IN2(n45), .Q(n30) );
  NAND3X0 U6 ( .IN1(n43), .IN2(n44), .IN3(n45), .QN(n42) );
  XOR2X1 U7 ( .IN1(n40), .IN2(n26), .Q(DIFF[5]) );
  XNOR2X1 U8 ( .IN1(n13), .IN2(B[28]), .Q(DIFF[28]) );
  XNOR2X1 U9 ( .IN1(n31), .IN2(B[29]), .Q(DIFF[29]) );
  AND2X1 U10 ( .IN1(n41), .IN2(n8), .Q(n26) );
  AND2X1 U11 ( .IN1(n26), .IN2(n40), .Q(n27) );
  AND2X1 U12 ( .IN1(n12), .IN2(n8), .Q(n9) );
  AND2X1 U13 ( .IN1(n37), .IN2(n9), .Q(n21) );
  AND2X1 U14 ( .IN1(n11), .IN2(n9), .Q(n10) );
  AND4X1 U15 ( .IN1(n20), .IN2(n51), .IN3(n50), .IN4(n3), .Q(n32) );
  INVX0 U16 ( .INP(B[29]), .ZN(n48) );
  XOR2X1 U17 ( .IN1(n6), .IN2(n35), .Q(DIFF[17]) );
  XOR2X1 U18 ( .IN1(n59), .IN2(n60), .Q(DIFF[18]) );
  XOR2X1 U19 ( .IN1(n15), .IN2(n54), .Q(DIFF[23]) );
  XOR2X1 U20 ( .IN1(n17), .IN2(n53), .Q(DIFF[24]) );
  XOR2X1 U21 ( .IN1(n18), .IN2(n52), .Q(DIFF[25]) );
  XOR2X1 U22 ( .IN1(n20), .IN2(n51), .Q(DIFF[26]) );
  AND2X1 U23 ( .IN1(n59), .IN2(n60), .Q(n1) );
  NAND4X0 U24 ( .IN1(n62), .IN2(n8), .IN3(n11), .IN4(n12), .QN(n2) );
  AND2X1 U25 ( .IN1(n48), .IN2(n49), .Q(n3) );
  AND3X1 U26 ( .IN1(n14), .IN2(n61), .IN3(n35), .Q(n59) );
  NOR4X1 U27 ( .IN1(B[11]), .IN2(B[10]), .IN3(B[9]), .IN4(B[8]), .QN(n11) );
  AND2X1 U28 ( .IN1(n4), .IN2(n5), .Q(n62) );
  NOR2X0 U29 ( .IN1(B[14]), .IN2(B[15]), .QN(n4) );
  NOR2X0 U30 ( .IN1(B[12]), .IN2(B[13]), .QN(n5) );
  NOR4X1 U31 ( .IN1(B[4]), .IN2(B[6]), .IN3(B[5]), .IN4(B[7]), .QN(n12) );
  AND2X1 U32 ( .IN1(n14), .IN2(n61), .Q(n6) );
  AND2X1 U33 ( .IN1(n59), .IN2(n7), .Q(n15) );
  NOR2X0 U34 ( .IN1(n16), .IN2(B[18]), .QN(n7) );
  XOR2X1 U35 ( .IN1(n19), .IN2(n50), .Q(DIFF[27]) );
  NOR4X1 U36 ( .IN1(B[1]), .IN2(\B[0] ), .IN3(B[2]), .IN4(B[3]), .QN(n8) );
  XNOR2X1 U37 ( .IN1(n32), .IN2(B[30]), .Q(DIFF[30]) );
  XOR2X1 U38 ( .IN1(n46), .IN2(B[31]), .Q(DIFF[31]) );
  XOR2X1 U39 ( .IN1(n28), .IN2(n65), .Q(DIFF[14]) );
  AND2X1 U40 ( .IN1(n19), .IN2(n50), .Q(n13) );
  AND4X1 U41 ( .IN1(n62), .IN2(n8), .IN3(n11), .IN4(n12), .Q(n14) );
  NAND2X1 U42 ( .IN1(n58), .IN2(n33), .QN(n16) );
  AND2X1 U43 ( .IN1(n15), .IN2(n54), .Q(n17) );
  AND2X1 U44 ( .IN1(n17), .IN2(n53), .Q(n18) );
  AND2X1 U45 ( .IN1(n20), .IN2(n51), .Q(n19) );
  AND2X1 U46 ( .IN1(n18), .IN2(n52), .Q(n20) );
  AND2X1 U47 ( .IN1(n23), .IN2(n57), .Q(n22) );
  AND2X1 U48 ( .IN1(n1), .IN2(n58), .Q(n23) );
  AND2X1 U49 ( .IN1(n10), .IN2(n63), .Q(n24) );
  AND2X1 U50 ( .IN1(n57), .IN2(n34), .Q(n33) );
  AND2X1 U51 ( .IN1(n56), .IN2(n55), .Q(n34) );
  AND2X1 U52 ( .IN1(n36), .IN2(n21), .Q(n25) );
  AND2X1 U53 ( .IN1(n24), .IN2(n64), .Q(n28) );
  AND2X1 U54 ( .IN1(n22), .IN2(n56), .Q(n29) );
  INVX0 U55 ( .INP(B[30]), .ZN(n47) );
  INVX0 U56 ( .INP(B[13]), .ZN(n64) );
  INVX0 U57 ( .INP(B[1]), .ZN(n45) );
  INVX0 U58 ( .INP(B[9]), .ZN(n36) );
  INVX0 U59 ( .INP(B[4]), .ZN(n41) );
  INVX0 U60 ( .INP(B[8]), .ZN(n37) );
  INVX0 U61 ( .INP(B[5]), .ZN(n40) );
  INVX0 U62 ( .INP(B[6]), .ZN(n39) );
  INVX0 U63 ( .INP(B[10]), .ZN(n67) );
  INVX0 U64 ( .INP(B[12]), .ZN(n63) );
  INVX0 U65 ( .INP(B[14]), .ZN(n65) );
  AND2X1 U66 ( .IN1(n49), .IN2(n13), .Q(n31) );
  INVX0 U67 ( .INP(B[2]), .ZN(n44) );
  XOR2X1 U68 ( .IN1(n29), .IN2(n55), .Q(DIFF[22]) );
  XOR2X1 U69 ( .IN1(n1), .IN2(n58), .Q(DIFF[19]) );
  XOR2X1 U70 ( .IN1(n22), .IN2(n56), .Q(DIFF[21]) );
  XOR2X1 U71 ( .IN1(n24), .IN2(n64), .Q(DIFF[13]) );
  XNOR2X1 U72 ( .IN1(n2), .IN2(n61), .Q(DIFF[16]) );
  XOR2X1 U73 ( .IN1(n21), .IN2(n36), .Q(DIFF[9]) );
  XOR2X1 U74 ( .IN1(n25), .IN2(n67), .Q(DIFF[10]) );
  XOR2X1 U75 ( .IN1(n27), .IN2(n39), .Q(DIFF[6]) );
  XOR2X1 U76 ( .IN1(n68), .IN2(B[11]), .Q(DIFF[11]) );
  XOR2X1 U77 ( .IN1(n38), .IN2(B[7]), .Q(DIFF[7]) );
  XOR2X1 U78 ( .IN1(n10), .IN2(n63), .Q(DIFF[12]) );
  XOR2X1 U79 ( .IN1(n9), .IN2(n37), .Q(DIFF[8]) );
  XNOR2X1 U80 ( .IN1(n30), .IN2(B[2]), .Q(DIFF[2]) );
  XOR2X1 U81 ( .IN1(n42), .IN2(B[3]), .Q(DIFF[3]) );
  XOR2X1 U82 ( .IN1(n8), .IN2(n41), .Q(DIFF[4]) );
  INVX0 U83 ( .INP(B[21]), .ZN(n56) );
  INVX0 U84 ( .INP(B[19]), .ZN(n58) );
  INVX0 U85 ( .INP(B[20]), .ZN(n57) );
  INVX0 U86 ( .INP(B[17]), .ZN(n35) );
  XOR2X1 U87 ( .IN1(n66), .IN2(B[15]), .Q(DIFF[15]) );
  INVX0 U88 ( .INP(B[22]), .ZN(n55) );
  INVX0 U89 ( .INP(B[16]), .ZN(n61) );
  INVX0 U90 ( .INP(B[18]), .ZN(n60) );
  INVX0 U91 ( .INP(B[24]), .ZN(n53) );
  INVX0 U92 ( .INP(B[23]), .ZN(n54) );
  INVX0 U93 ( .INP(B[25]), .ZN(n52) );
  INVX0 U94 ( .INP(B[26]), .ZN(n51) );
  INVX0 U95 ( .INP(B[27]), .ZN(n50) );
  XOR2X1 U96 ( .IN1(n23), .IN2(n57), .Q(DIFF[20]) );
  NAND2X0 U97 ( .IN1(n25), .IN2(n67), .QN(n68) );
  NAND2X0 U98 ( .IN1(n27), .IN2(n39), .QN(n38) );
  INVX0 U99 ( .INP(\B[0] ), .ZN(n43) );
  NAND2X0 U100 ( .IN1(n28), .IN2(n65), .QN(n66) );
  NAND2X0 U101 ( .IN1(n47), .IN2(n32), .QN(n46) );
endmodule


module SeqMult_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;

  NAND3X0 U2 ( .IN1(A[28]), .IN2(A[29]), .IN3(n17), .QN(n15) );
  XNOR2X1 U3 ( .IN1(A[29]), .IN2(n1), .Q(SUM[29]) );
  XOR2X1 U4 ( .IN1(A[28]), .IN2(n17), .Q(SUM[28]) );
  XOR2X1 U5 ( .IN1(A[20]), .IN2(n32), .Q(SUM[20]) );
  XOR2X1 U6 ( .IN1(A[16]), .IN2(n41), .Q(SUM[16]) );
  XOR2X1 U7 ( .IN1(A[11]), .IN2(n56), .Q(SUM[11]) );
  NAND2X0 U8 ( .IN1(A[3]), .IN2(A[2]), .QN(n61) );
  NAND2X0 U9 ( .IN1(A[28]), .IN2(n17), .QN(n1) );
  NOR2X0 U10 ( .IN1(n6), .IN2(n59), .QN(n4) );
  NOR2X0 U11 ( .IN1(n54), .IN2(n55), .QN(n50) );
  NOR2X0 U12 ( .IN1(n12), .IN2(n61), .QN(n10) );
  NOR2X0 U13 ( .IN1(n36), .IN2(n37), .QN(n32) );
  NAND2X1 U14 ( .IN1(A[19]), .IN2(A[18]), .QN(n37) );
  NOR2X0 U15 ( .IN1(n45), .IN2(n46), .QN(n41) );
  NOR2X0 U16 ( .IN1(n27), .IN2(n28), .QN(n23) );
  NAND2X1 U17 ( .IN1(A[23]), .IN2(A[22]), .QN(n28) );
  NAND2X1 U18 ( .IN1(n58), .IN2(n4), .QN(n54) );
  NOR2X0 U19 ( .IN1(n2), .IN2(n63), .QN(n58) );
  INVX0 U20 ( .INP(A[8]), .ZN(n63) );
  NAND2X1 U21 ( .IN1(n49), .IN2(n50), .QN(n45) );
  NOR2X0 U22 ( .IN1(n51), .IN2(n52), .QN(n49) );
  INVX0 U23 ( .INP(A[12]), .ZN(n52) );
  NOR2X0 U24 ( .IN1(n18), .IN2(n19), .QN(n17) );
  NAND2X1 U25 ( .IN1(A[27]), .IN2(A[26]), .QN(n19) );
  NAND2X1 U26 ( .IN1(n40), .IN2(n41), .QN(n36) );
  NOR2X0 U27 ( .IN1(n42), .IN2(n43), .QN(n40) );
  INVX0 U28 ( .INP(A[16]), .ZN(n43) );
  NAND2X1 U29 ( .IN1(A[1]), .IN2(A[0]), .QN(n12) );
  NAND2X1 U30 ( .IN1(n31), .IN2(n32), .QN(n27) );
  NOR2X0 U31 ( .IN1(n33), .IN2(n34), .QN(n31) );
  INVX0 U32 ( .INP(A[20]), .ZN(n34) );
  NAND2X1 U33 ( .IN1(n60), .IN2(n10), .QN(n6) );
  NOR2X0 U34 ( .IN1(n8), .IN2(n62), .QN(n60) );
  INVX0 U35 ( .INP(A[4]), .ZN(n62) );
  NAND2X1 U36 ( .IN1(n22), .IN2(n23), .QN(n18) );
  NOR2X0 U37 ( .IN1(n24), .IN2(n25), .QN(n22) );
  INVX0 U38 ( .INP(A[13]), .ZN(n51) );
  INVX0 U39 ( .INP(A[5]), .ZN(n8) );
  INVX0 U40 ( .INP(A[9]), .ZN(n2) );
  XOR2X1 U41 ( .IN1(A[24]), .IN2(n23), .Q(SUM[24]) );
  NOR2X0 U42 ( .IN1(n15), .IN2(n16), .QN(n14) );
  NOR2X0 U43 ( .IN1(n18), .IN2(n21), .QN(n20) );
  NOR2X0 U44 ( .IN1(n27), .IN2(n30), .QN(n29) );
  NAND2X0 U45 ( .IN1(A[20]), .IN2(n32), .QN(n35) );
  INVX0 U46 ( .INP(A[21]), .ZN(n33) );
  INVX0 U47 ( .INP(A[17]), .ZN(n42) );
  XOR2X1 U48 ( .IN1(A[15]), .IN2(n47), .Q(SUM[15]) );
  NOR2X0 U49 ( .IN1(n45), .IN2(n48), .QN(n47) );
  XOR2X1 U50 ( .IN1(A[7]), .IN2(n5), .Q(SUM[7]) );
  NOR2X0 U51 ( .IN1(n6), .IN2(n7), .QN(n5) );
  NOR2X0 U52 ( .IN1(n12), .IN2(n13), .QN(n11) );
  INVX0 U53 ( .INP(A[0]), .ZN(SUM[0]) );
  NOR2X0 U54 ( .IN1(n36), .IN2(n39), .QN(n38) );
  NAND2X0 U55 ( .IN1(A[12]), .IN2(n50), .QN(n53) );
  NOR2X0 U56 ( .IN1(n54), .IN2(n57), .QN(n56) );
  NAND2X0 U57 ( .IN1(A[8]), .IN2(n4), .QN(n3) );
  NAND2X0 U58 ( .IN1(A[4]), .IN2(n10), .QN(n9) );
  INVX0 U59 ( .INP(A[6]), .ZN(n7) );
  INVX0 U60 ( .INP(A[26]), .ZN(n21) );
  INVX0 U61 ( .INP(A[22]), .ZN(n30) );
  INVX0 U62 ( .INP(A[18]), .ZN(n39) );
  INVX0 U63 ( .INP(A[2]), .ZN(n13) );
  INVX0 U64 ( .INP(A[14]), .ZN(n48) );
  INVX0 U65 ( .INP(A[10]), .ZN(n57) );
  INVX0 U66 ( .INP(A[25]), .ZN(n24) );
  INVX0 U67 ( .INP(A[30]), .ZN(n16) );
  NAND2X0 U68 ( .IN1(A[7]), .IN2(A[6]), .QN(n59) );
  INVX0 U69 ( .INP(A[24]), .ZN(n25) );
  NAND2X0 U70 ( .IN1(A[11]), .IN2(A[10]), .QN(n55) );
  NAND2X0 U71 ( .IN1(A[15]), .IN2(A[14]), .QN(n46) );
  NAND2X0 U72 ( .IN1(A[16]), .IN2(n41), .QN(n44) );
  NAND2X0 U73 ( .IN1(A[24]), .IN2(n23), .QN(n26) );
  XOR2X1 U74 ( .IN1(n2), .IN2(n3), .Q(SUM[9]) );
  XOR2X1 U75 ( .IN1(A[8]), .IN2(n4), .Q(SUM[8]) );
  XOR2X1 U76 ( .IN1(n7), .IN2(n6), .Q(SUM[6]) );
  XOR2X1 U77 ( .IN1(n8), .IN2(n9), .Q(SUM[5]) );
  XOR2X1 U78 ( .IN1(A[4]), .IN2(n10), .Q(SUM[4]) );
  XOR2X1 U79 ( .IN1(A[3]), .IN2(n11), .Q(SUM[3]) );
  XOR2X1 U80 ( .IN1(A[31]), .IN2(n14), .Q(SUM[31]) );
  XOR2X1 U81 ( .IN1(n16), .IN2(n15), .Q(SUM[30]) );
  XOR2X1 U82 ( .IN1(n13), .IN2(n12), .Q(SUM[2]) );
  XOR2X1 U83 ( .IN1(A[27]), .IN2(n20), .Q(SUM[27]) );
  XOR2X1 U84 ( .IN1(n21), .IN2(n18), .Q(SUM[26]) );
  XOR2X1 U85 ( .IN1(n24), .IN2(n26), .Q(SUM[25]) );
  XOR2X1 U86 ( .IN1(A[23]), .IN2(n29), .Q(SUM[23]) );
  XOR2X1 U87 ( .IN1(n30), .IN2(n27), .Q(SUM[22]) );
  XOR2X1 U88 ( .IN1(n33), .IN2(n35), .Q(SUM[21]) );
  XOR2X1 U89 ( .IN1(A[1]), .IN2(A[0]), .Q(SUM[1]) );
  XOR2X1 U90 ( .IN1(A[19]), .IN2(n38), .Q(SUM[19]) );
  XOR2X1 U91 ( .IN1(n39), .IN2(n36), .Q(SUM[18]) );
  XOR2X1 U92 ( .IN1(n42), .IN2(n44), .Q(SUM[17]) );
  XOR2X1 U93 ( .IN1(n48), .IN2(n45), .Q(SUM[14]) );
  XOR2X1 U94 ( .IN1(n51), .IN2(n53), .Q(SUM[13]) );
  XOR2X1 U95 ( .IN1(A[12]), .IN2(n50), .Q(SUM[12]) );
  XOR2X1 U96 ( .IN1(n57), .IN2(n54), .Q(SUM[10]) );
endmodule


module SeqMult_DW01_sub_8 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  NOR4X1 U3 ( .IN1(B[46]), .IN2(B[45]), .IN3(B[47]), .IN4(B[44]), .QN(n146) );
  NOR4X0 U4 ( .IN1(B[7]), .IN2(B[6]), .IN3(B[5]), .IN4(B[4]), .QN(n94) );
  NOR4X0 U5 ( .IN1(B[11]), .IN2(B[10]), .IN3(B[9]), .IN4(B[8]), .QN(n93) );
  NBUFFX2 U6 ( .INP(B[57]), .Z(n6) );
  AND2X1 U7 ( .IN1(n20), .IN2(n139), .Q(n22) );
  AND2X1 U8 ( .IN1(n11), .IN2(n8), .Q(n118) );
  AND2X1 U9 ( .IN1(n10), .IN2(n163), .Q(n81) );
  AND2X1 U10 ( .IN1(n92), .IN2(n37), .Q(n85) );
  NBUFFX4 U11 ( .INP(B[58]), .Z(n46) );
  AND2X1 U12 ( .IN1(n22), .IN2(n45), .Q(n51) );
  AND2X1 U13 ( .IN1(n22), .IN2(n138), .Q(n63) );
  AND2X1 U14 ( .IN1(n77), .IN2(n84), .Q(n56) );
  AND2X1 U15 ( .IN1(n73), .IN2(n10), .Q(n79) );
  AND2X1 U16 ( .IN1(n37), .IN2(n187), .Q(n95) );
  AND2X1 U17 ( .IN1(n82), .IN2(n194), .Q(n106) );
  AND2X1 U18 ( .IN1(n120), .IN2(n103), .Q(n104) );
  AND2X1 U19 ( .IN1(n127), .IN2(n2), .Q(n36) );
  AND2X1 U20 ( .IN1(n22), .IN2(n53), .Q(n71) );
  AND2X1 U21 ( .IN1(n12), .IN2(n10), .Q(n80) );
  AND2X1 U22 ( .IN1(n75), .IN2(n165), .Q(n76) );
  AND2X1 U23 ( .IN1(n99), .IN2(n176), .Q(n90) );
  XNOR2X1 U24 ( .IN1(n91), .IN2(B[28]), .Q(DIFF[28]) );
  AND2X1 U25 ( .IN1(n98), .IN2(n183), .Q(n102) );
  XNOR2X1 U26 ( .IN1(n202), .IN2(n208), .Q(DIFF[12]) );
  XNOR2X1 U27 ( .IN1(n122), .IN2(n121), .Q(DIFF[8]) );
  XNOR2X1 U28 ( .IN1(n125), .IN2(n131), .Q(DIFF[5]) );
  XNOR2X1 U29 ( .IN1(n132), .IN2(n143), .Q(DIFF[4]) );
  XNOR2X1 U30 ( .IN1(n179), .IN2(\B[0] ), .Q(DIFF[1]) );
  NBUFFX4 U31 ( .INP(B[61]), .Z(n1) );
  AND3X1 U32 ( .IN1(n26), .IN2(n21), .IN3(n130), .Q(n2) );
  INVX0 U33 ( .INP(n135), .ZN(n3) );
  OR2X1 U34 ( .IN1(B[39]), .IN2(B[37]), .Q(n4) );
  NAND2X1 U35 ( .IN1(n195), .IN2(n89), .QN(n5) );
  NOR4X1 U36 ( .IN1(B[43]), .IN2(B[42]), .IN3(B[41]), .IN4(B[40]), .QN(n11) );
  AND2X1 U37 ( .IN1(n32), .IN2(n53), .Q(n72) );
  AND2X1 U38 ( .IN1(n51), .IN2(n53), .Q(n69) );
  AND2X1 U39 ( .IN1(n63), .IN2(n53), .Q(n70) );
  AND2X1 U40 ( .IN1(n53), .IN2(n140), .Q(n74) );
  NOR2X0 U41 ( .IN1(n17), .IN2(n18), .QN(n53) );
  DELLN1X2 U42 ( .INP(B[53]), .Z(n7) );
  NOR3X0 U43 ( .IN1(B[38]), .IN2(B[36]), .IN3(n4), .QN(n8) );
  INVX0 U44 ( .INP(n140), .ZN(n9) );
  NOR3X0 U45 ( .IN1(n23), .IN2(B[28]), .IN3(n24), .QN(n10) );
  AND2X1 U46 ( .IN1(n52), .IN2(n35), .Q(n27) );
  AND4X1 U47 ( .IN1(n51), .IN2(n12), .IN3(n13), .IN4(n137), .Q(n55) );
  INVX0 U48 ( .INP(n17), .ZN(n12) );
  INVX0 U49 ( .INP(n18), .ZN(n13) );
  NOR3X0 U50 ( .IN1(B[57]), .IN2(B[56]), .IN3(B[55]), .QN(n19) );
  AND3X1 U51 ( .IN1(n183), .IN2(n174), .IN3(n175), .Q(n173) );
  NOR4X1 U52 ( .IN1(n5), .IN2(B[19]), .IN3(n199), .IN4(n83), .QN(n37) );
  NAND4X0 U53 ( .IN1(n128), .IN2(n130), .IN3(n54), .IN4(n40), .QN(n129) );
  NOR2X0 U54 ( .IN1(B[56]), .IN2(B[55]), .QN(n14) );
  NOR4X1 U55 ( .IN1(B[2]), .IN2(\B[0] ), .IN3(B[1]), .IN4(B[3]), .QN(n15) );
  NOR2X0 U56 ( .IN1(n16), .IN2(B[58]), .QN(n40) );
  NAND2X0 U57 ( .IN1(n134), .IN2(n14), .QN(n16) );
  NAND4X0 U58 ( .IN1(n146), .IN2(n8), .IN3(n11), .IN4(n73), .QN(n17) );
  NAND2X0 U59 ( .IN1(n10), .IN2(n145), .QN(n18) );
  NOR2X0 U60 ( .IN1(B[49]), .IN2(B[50]), .QN(n20) );
  AND2X1 U61 ( .IN1(n133), .IN2(n19), .Q(n21) );
  XNOR2X1 U62 ( .IN1(n25), .IN2(B[60]), .Q(DIFF[60]) );
  NOR4X0 U63 ( .IN1(B[43]), .IN2(B[42]), .IN3(B[41]), .IN4(B[40]), .QN(n31) );
  NOR3X0 U64 ( .IN1(n23), .IN2(B[28]), .IN3(n24), .QN(n88) );
  NAND4X0 U65 ( .IN1(n37), .IN2(n92), .IN3(n172), .IN4(n173), .QN(n23) );
  NAND2X0 U66 ( .IN1(n41), .IN2(n176), .QN(n24) );
  AND3X1 U67 ( .IN1(n26), .IN2(n130), .IN3(n40), .Q(n25) );
  AND3X1 U68 ( .IN1(n34), .IN2(n78), .IN3(n137), .Q(n26) );
  NAND2X0 U69 ( .IN1(n58), .IN2(n35), .QN(n28) );
  INVX0 U70 ( .INP(B[56]), .ZN(n29) );
  INVX0 U71 ( .INP(n29), .ZN(n30) );
  NOR2X0 U72 ( .IN1(n142), .IN2(n9), .QN(n32) );
  XOR2X1 U73 ( .IN1(B[62]), .IN2(n33), .Q(DIFF[62]) );
  NAND2X0 U74 ( .IN1(n42), .IN2(n127), .QN(n33) );
  AND2X1 U75 ( .IN1(n60), .IN2(n45), .Q(n34) );
  INVX0 U76 ( .INP(B[45]), .ZN(n35) );
  NOR2X0 U77 ( .IN1(n3), .IN2(n30), .QN(n38) );
  XOR2X1 U78 ( .IN1(n6), .IN2(n48), .Q(DIFF[57]) );
  NOR3X0 U79 ( .IN1(B[38]), .IN2(B[36]), .IN3(n4), .QN(n84) );
  INVX0 U80 ( .INP(B[53]), .ZN(n39) );
  NOR2X0 U81 ( .IN1(B[26]), .IN2(n182), .QN(n181) );
  NOR2X0 U82 ( .IN1(B[29]), .IN2(B[31]), .QN(n41) );
  AND3X1 U83 ( .IN1(n26), .IN2(n21), .IN3(n130), .Q(n42) );
  NOR2X0 U84 ( .IN1(n43), .IN2(n44), .QN(n78) );
  NAND4X0 U85 ( .IN1(n146), .IN2(n84), .IN3(n31), .IN4(n73), .QN(n43) );
  NAND2X0 U86 ( .IN1(n145), .IN2(n10), .QN(n44) );
  AND2X1 U87 ( .IN1(n56), .IN2(n152), .Q(n57) );
  AND2X1 U88 ( .IN1(n39), .IN2(n138), .Q(n45) );
  NOR2X0 U89 ( .IN1(B[49]), .IN2(B[50]), .QN(n62) );
  XOR2X1 U90 ( .IN1(n30), .IN2(n47), .Q(DIFF[56]) );
  NAND2X0 U91 ( .IN1(n55), .IN2(n135), .QN(n47) );
  NAND2X0 U92 ( .IN1(n126), .IN2(n36), .QN(DIFF[63]) );
  NAND2X0 U93 ( .IN1(n38), .IN2(n55), .QN(n48) );
  XOR2X1 U94 ( .IN1(n49), .IN2(n46), .Q(DIFF[58]) );
  NAND2X0 U95 ( .IN1(n55), .IN2(n19), .QN(n49) );
  XOR2X1 U96 ( .IN1(B[59]), .IN2(n50), .Q(DIFF[59]) );
  NAND2X0 U97 ( .IN1(n55), .IN2(n21), .QN(n50) );
  XOR2X1 U98 ( .IN1(n1), .IN2(n129), .Q(DIFF[61]) );
  INVX0 U99 ( .INP(B[46]), .ZN(n52) );
  AND3X1 U100 ( .IN1(n34), .IN2(n137), .IN3(n78), .Q(n54) );
  NAND2X0 U101 ( .IN1(n202), .IN2(n203), .QN(n201) );
  NAND2X0 U102 ( .IN1(n174), .IN2(n175), .QN(n182) );
  NAND2X0 U103 ( .IN1(n204), .IN2(n205), .QN(n200) );
  INVX0 U104 ( .INP(n64), .ZN(n153) );
  INVX0 U105 ( .INP(n61), .ZN(n161) );
  INVX0 U106 ( .INP(n57), .ZN(n154) );
  INVX0 U107 ( .INP(n75), .ZN(n167) );
  INVX0 U108 ( .INP(n66), .ZN(n159) );
  AND2X1 U109 ( .IN1(n67), .IN2(n147), .Q(n58) );
  AND2X1 U110 ( .IN1(n64), .IN2(n150), .Q(n59) );
  AND2X1 U111 ( .IN1(n139), .IN2(n62), .Q(n60) );
  AND2X1 U112 ( .IN1(n77), .IN2(n157), .Q(n61) );
  AND2X1 U113 ( .IN1(n57), .IN2(n151), .Q(n64) );
  AND2X1 U114 ( .IN1(n66), .IN2(n156), .Q(n65) );
  AND2X1 U115 ( .IN1(n61), .IN2(n160), .Q(n66) );
  AND2X1 U116 ( .IN1(n118), .IN2(n79), .Q(n67) );
  AND2X1 U117 ( .IN1(n27), .IN2(n58), .Q(n68) );
  AND4X1 U118 ( .IN1(n163), .IN2(n164), .IN3(n165), .IN4(n166), .Q(n73) );
  AND2X1 U119 ( .IN1(n81), .IN2(n164), .Q(n75) );
  INVX0 U120 ( .INP(n53), .ZN(n144) );
  INVX0 U121 ( .INP(n81), .ZN(n168) );
  INVX0 U122 ( .INP(n79), .ZN(n162) );
  INVX0 U123 ( .INP(B[33]), .ZN(n164) );
  INVX0 U124 ( .INP(n15), .ZN(n143) );
  INVX0 U125 ( .INP(n37), .ZN(n192) );
  INVX0 U126 ( .INP(n82), .ZN(n198) );
  INVX0 U127 ( .INP(n86), .ZN(n121) );
  INVX0 U128 ( .INP(n85), .ZN(n185) );
  INVX0 U129 ( .INP(n87), .ZN(n208) );
  INVX0 U130 ( .INP(n141), .ZN(n142) );
  AND2X1 U131 ( .IN1(n73), .IN2(n88), .Q(n77) );
  INVX0 U132 ( .INP(B[57]), .ZN(n134) );
  INVX0 U133 ( .INP(B[49]), .ZN(n140) );
  INVX0 U134 ( .INP(B[50]), .ZN(n141) );
  INVX0 U135 ( .INP(B[34]), .ZN(n165) );
  INVX0 U136 ( .INP(B[38]), .ZN(n156) );
  NOR2X0 U137 ( .IN1(n199), .IN2(n83), .QN(n82) );
  OR2X1 U138 ( .IN1(n200), .IN2(n201), .Q(n83) );
  INVX0 U139 ( .INP(B[52]), .ZN(n138) );
  INVX0 U140 ( .INP(B[58]), .ZN(n133) );
  INVX0 U141 ( .INP(B[40]), .ZN(n152) );
  INVX0 U142 ( .INP(B[36]), .ZN(n157) );
  INVX0 U143 ( .INP(B[41]), .ZN(n151) );
  INVX0 U144 ( .INP(B[42]), .ZN(n150) );
  INVX0 U145 ( .INP(B[44]), .ZN(n147) );
  INVX0 U146 ( .INP(B[55]), .ZN(n135) );
  INVX0 U147 ( .INP(B[48]), .ZN(n145) );
  INVX0 U148 ( .INP(B[54]), .ZN(n137) );
  INVX0 U149 ( .INP(B[35]), .ZN(n166) );
  INVX0 U150 ( .INP(B[51]), .ZN(n139) );
  INVX0 U151 ( .INP(n100), .ZN(n180) );
  AND2X1 U152 ( .IN1(n94), .IN2(n15), .Q(n86) );
  INVX0 U153 ( .INP(B[37]), .ZN(n160) );
  INVX0 U154 ( .INP(B[32]), .ZN(n163) );
  AND2X1 U155 ( .IN1(n93), .IN2(n86), .Q(n87) );
  INVX0 U156 ( .INP(n97), .ZN(n184) );
  INVX0 U157 ( .INP(n106), .ZN(n197) );
  INVX0 U158 ( .INP(n111), .ZN(n206) );
  INVX0 U159 ( .INP(n108), .ZN(n207) );
  INVX0 U160 ( .INP(n109), .ZN(n196) );
  INVX0 U161 ( .INP(n103), .ZN(n119) );
  INVX0 U162 ( .INP(n95), .ZN(n191) );
  INVX0 U163 ( .INP(n110), .ZN(n124) );
  INVX0 U164 ( .INP(n107), .ZN(n177) );
  INVX0 U165 ( .INP(n96), .ZN(n190) );
  INVX0 U166 ( .INP(n104), .ZN(n210) );
  INVX0 U167 ( .INP(n105), .ZN(n131) );
  AND2X1 U168 ( .IN1(n193), .IN2(n194), .Q(n89) );
  AND3X1 U169 ( .IN1(n85), .IN2(n172), .IN3(n181), .Q(n91) );
  AND4X1 U170 ( .IN1(n186), .IN2(n187), .IN3(n188), .IN4(n189), .Q(n92) );
  INVX0 U171 ( .INP(B[59]), .ZN(n130) );
  AND2X1 U172 ( .IN1(n95), .IN2(n186), .Q(n96) );
  INVX0 U173 ( .INP(B[60]), .ZN(n128) );
  AND2X1 U174 ( .IN1(n85), .IN2(n175), .Q(n97) );
  AND2X1 U175 ( .IN1(n97), .IN2(n174), .Q(n98) );
  AND2X1 U176 ( .IN1(n100), .IN2(n171), .Q(n99) );
  AND2X1 U177 ( .IN1(n91), .IN2(n170), .Q(n100) );
  AND2X1 U178 ( .IN1(n96), .IN2(n188), .Q(n101) );
  AND2X1 U179 ( .IN1(n122), .IN2(n86), .Q(n103) );
  AND2X1 U180 ( .IN1(n132), .IN2(n15), .Q(n105) );
  AND2X1 U181 ( .IN1(n178), .IN2(n179), .Q(n107) );
  AND2X1 U182 ( .IN1(n87), .IN2(n202), .Q(n108) );
  AND2X1 U183 ( .IN1(n106), .IN2(n195), .Q(n109) );
  AND2X1 U184 ( .IN1(n105), .IN2(n125), .Q(n110) );
  AND2X1 U185 ( .IN1(n108), .IN2(n204), .Q(n111) );
  AND2X1 U186 ( .IN1(n109), .IN2(n193), .Q(n112) );
  AND2X1 U187 ( .IN1(n104), .IN2(n209), .Q(n113) );
  AND2X1 U188 ( .IN1(n111), .IN2(n203), .Q(n114) );
  AND2X1 U189 ( .IN1(n107), .IN2(n158), .Q(n115) );
  AND2X1 U190 ( .IN1(n110), .IN2(n123), .Q(n116) );
  INVX0 U191 ( .INP(B[29]), .ZN(n171) );
  INVX0 U192 ( .INP(B[30]), .ZN(n176) );
  INVX0 U193 ( .INP(B[24]), .ZN(n175) );
  INVX0 U194 ( .INP(B[25]), .ZN(n174) );
  INVX0 U195 ( .INP(B[16]), .ZN(n194) );
  INVX0 U196 ( .INP(B[14]), .ZN(n203) );
  INVX0 U197 ( .INP(B[18]), .ZN(n193) );
  INVX0 U198 ( .INP(B[13]), .ZN(n204) );
  INVX0 U199 ( .INP(B[12]), .ZN(n202) );
  INVX0 U200 ( .INP(B[17]), .ZN(n195) );
  INVX0 U201 ( .INP(B[28]), .ZN(n170) );
  INVX0 U202 ( .INP(B[5]), .ZN(n125) );
  INVX0 U203 ( .INP(B[20]), .ZN(n187) );
  INVX0 U204 ( .INP(B[10]), .ZN(n209) );
  INVX0 U205 ( .INP(B[6]), .ZN(n123) );
  INVX0 U206 ( .INP(B[1]), .ZN(n179) );
  INVX0 U207 ( .INP(B[9]), .ZN(n120) );
  INVX0 U208 ( .INP(B[8]), .ZN(n122) );
  INVX0 U209 ( .INP(B[4]), .ZN(n132) );
  INVX0 U210 ( .INP(B[21]), .ZN(n186) );
  INVX0 U211 ( .INP(B[2]), .ZN(n158) );
  INVX0 U212 ( .INP(B[26]), .ZN(n183) );
  INVX0 U213 ( .INP(B[15]), .ZN(n205) );
  INVX0 U214 ( .INP(\B[0] ), .ZN(n178) );
  INVX0 U215 ( .INP(B[27]), .ZN(n172) );
  INVX0 U216 ( .INP(B[23]), .ZN(n189) );
  INVX0 U217 ( .INP(B[22]), .ZN(n188) );
  XNOR2X1 U218 ( .IN1(n59), .IN2(B[43]), .Q(DIFF[43]) );
  XNOR2X1 U219 ( .IN1(n68), .IN2(B[47]), .Q(DIFF[47]) );
  XNOR2X1 U220 ( .IN1(n65), .IN2(B[39]), .Q(DIFF[39]) );
  XNOR2X1 U221 ( .IN1(n153), .IN2(n150), .Q(DIFF[42]) );
  XNOR2X1 U222 ( .IN1(n28), .IN2(n52), .Q(DIFF[46]) );
  XNOR2X1 U223 ( .IN1(n159), .IN2(n156), .Q(DIFF[38]) );
  XNOR2X1 U224 ( .IN1(n76), .IN2(B[35]), .Q(DIFF[35]) );
  XNOR2X1 U225 ( .IN1(n154), .IN2(n151), .Q(DIFF[41]) );
  XNOR2X1 U226 ( .IN1(n148), .IN2(n35), .Q(DIFF[45]) );
  XNOR2X1 U227 ( .IN1(n167), .IN2(n165), .Q(DIFF[34]) );
  XNOR2X1 U228 ( .IN1(n161), .IN2(n160), .Q(DIFF[37]) );
  XNOR2X1 U229 ( .IN1(n90), .IN2(B[31]), .Q(DIFF[31]) );
  XNOR2X1 U230 ( .IN1(n149), .IN2(n147), .Q(DIFF[44]) );
  XNOR2X1 U231 ( .IN1(n155), .IN2(n152), .Q(DIFF[40]) );
  XNOR2X1 U232 ( .IN1(n74), .IN2(n142), .Q(DIFF[50]) );
  XNOR2X1 U233 ( .IN1(n69), .IN2(B[54]), .Q(DIFF[54]) );
  XNOR2X1 U234 ( .IN1(n70), .IN2(n7), .Q(DIFF[53]) );
  XNOR2X1 U235 ( .IN1(n71), .IN2(B[52]), .Q(DIFF[52]) );
  XNOR2X1 U236 ( .IN1(n72), .IN2(B[51]), .Q(DIFF[51]) );
  XNOR2X1 U237 ( .IN1(n102), .IN2(B[27]), .Q(DIFF[27]) );
  XNOR2X1 U238 ( .IN1(n168), .IN2(n164), .Q(DIFF[33]) );
  XNOR2X1 U239 ( .IN1(n162), .IN2(n157), .Q(DIFF[36]) );
  XNOR2X1 U240 ( .IN1(n99), .IN2(B[30]), .Q(DIFF[30]) );
  XNOR2X1 U241 ( .IN1(n80), .IN2(B[48]), .Q(DIFF[48]) );
  XNOR2X1 U242 ( .IN1(n180), .IN2(n171), .Q(DIFF[29]) );
  XNOR2X1 U243 ( .IN1(n98), .IN2(B[26]), .Q(DIFF[26]) );
  XNOR2X1 U244 ( .IN1(n169), .IN2(n163), .Q(DIFF[32]) );
  XNOR2X1 U245 ( .IN1(n101), .IN2(B[23]), .Q(DIFF[23]) );
  XNOR2X1 U246 ( .IN1(n136), .IN2(n135), .Q(DIFF[55]) );
  XNOR2X1 U247 ( .IN1(n144), .IN2(n140), .Q(DIFF[49]) );
  XNOR2X1 U248 ( .IN1(n114), .IN2(B[15]), .Q(DIFF[15]) );
  XNOR2X1 U249 ( .IN1(n190), .IN2(n188), .Q(DIFF[22]) );
  XNOR2X1 U250 ( .IN1(n206), .IN2(n203), .Q(DIFF[14]) );
  XNOR2X1 U251 ( .IN1(n112), .IN2(B[19]), .Q(DIFF[19]) );
  XNOR2X1 U252 ( .IN1(n113), .IN2(B[11]), .Q(DIFF[11]) );
  XNOR2X1 U253 ( .IN1(n191), .IN2(n186), .Q(DIFF[21]) );
  XNOR2X1 U254 ( .IN1(n196), .IN2(n193), .Q(DIFF[18]) );
  XNOR2X1 U255 ( .IN1(n210), .IN2(n209), .Q(DIFF[10]) );
  XNOR2X1 U256 ( .IN1(n207), .IN2(n204), .Q(DIFF[13]) );
  XNOR2X1 U257 ( .IN1(n116), .IN2(B[7]), .Q(DIFF[7]) );
  XNOR2X1 U258 ( .IN1(n192), .IN2(n187), .Q(DIFF[20]) );
  XNOR2X1 U259 ( .IN1(n197), .IN2(n195), .Q(DIFF[17]) );
  XNOR2X1 U260 ( .IN1(n119), .IN2(n120), .Q(DIFF[9]) );
  XNOR2X1 U261 ( .IN1(n124), .IN2(n123), .Q(DIFF[6]) );
  XNOR2X1 U262 ( .IN1(n198), .IN2(n194), .Q(DIFF[16]) );
  XNOR2X1 U263 ( .IN1(n115), .IN2(B[3]), .Q(DIFF[3]) );
  XNOR2X1 U264 ( .IN1(n177), .IN2(n158), .Q(DIFF[2]) );
  XNOR2X1 U265 ( .IN1(n184), .IN2(n174), .Q(DIFF[25]) );
  XNOR2X1 U266 ( .IN1(n185), .IN2(n175), .Q(DIFF[24]) );
  INVX0 U267 ( .INP(n67), .ZN(n149) );
  INVX0 U268 ( .INP(n10), .ZN(n169) );
  INVX0 U269 ( .INP(n58), .ZN(n148) );
  INVX0 U270 ( .INP(n55), .ZN(n136) );
  NOR2X0 U271 ( .IN1(B[60]), .IN2(B[61]), .QN(n127) );
  INVX0 U272 ( .INP(n56), .ZN(n155) );
  INVX0 U273 ( .INP(B[62]), .ZN(n126) );
  NAND3X0 U274 ( .IN1(n15), .IN2(n94), .IN3(n93), .QN(n199) );
endmodule


module SeqMult_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379;

  OR2X2 U2 ( .IN1(B[5]), .IN2(A[5]), .Q(n119) );
  NAND2X1 U3 ( .IN1(A[5]), .IN2(B[5]), .QN(n191) );
  INVX0 U4 ( .INP(n294), .ZN(n1) );
  NAND2X1 U5 ( .IN1(n2), .IN2(n25), .QN(n276) );
  NOR2X0 U6 ( .IN1(n165), .IN2(n1), .QN(n2) );
  XOR2X2 U7 ( .IN1(n271), .IN2(n272), .Q(SUM[21]) );
  OR2X1 U8 ( .IN1(B[15]), .IN2(A[15]), .Q(n71) );
  OR2X1 U9 ( .IN1(B[7]), .IN2(A[7]), .Q(n187) );
  OR2X1 U10 ( .IN1(B[15]), .IN2(A[15]), .Q(n317) );
  NAND3X0 U11 ( .IN1(n315), .IN2(n316), .IN3(n71), .QN(n306) );
  OR2X1 U12 ( .IN1(n332), .IN2(n333), .Q(n166) );
  NBUFFX2 U13 ( .INP(n191), .Z(n28) );
  AND2X1 U14 ( .IN1(n240), .IN2(n242), .Q(n170) );
  XOR2X1 U15 ( .IN1(n98), .IN2(n211), .Q(SUM[4]) );
  XOR3X1 U16 ( .IN1(B[28]), .IN2(A[28]), .IN3(n60), .Q(SUM[28]) );
  XNOR2X1 U17 ( .IN1(n130), .IN2(B[31]), .Q(SUM[31]) );
  AND2X1 U18 ( .IN1(B[16]), .IN2(A[16]), .Q(n150) );
  AND2X1 U19 ( .IN1(n65), .IN2(n6), .Q(n70) );
  INVX0 U20 ( .INP(n243), .ZN(n94) );
  AND2X1 U21 ( .IN1(n244), .IN2(n136), .Q(n110) );
  XNOR2X1 U22 ( .IN1(n184), .IN2(n185), .Q(SUM[7]) );
  AND2X1 U23 ( .IN1(B[8]), .IN2(A[8]), .Q(n173) );
  XOR2X1 U24 ( .IN1(n357), .IN2(n358), .Q(SUM[11]) );
  NBUFFX2 U25 ( .INP(B[13]), .Z(n26) );
  AND2X1 U26 ( .IN1(n146), .IN2(n152), .Q(n103) );
  XNOR2X1 U27 ( .IN1(n160), .IN2(n347), .Q(SUM[12]) );
  AND2X1 U28 ( .IN1(n299), .IN2(n298), .Q(n72) );
  XOR2X1 U29 ( .IN1(n77), .IN2(n76), .Q(SUM[18]) );
  AND2X1 U30 ( .IN1(n294), .IN2(n292), .Q(n76) );
  AND2X1 U31 ( .IN1(n142), .IN2(n111), .Q(n141) );
  XOR2X1 U32 ( .IN1(n256), .IN2(n257), .Q(SUM[24]) );
  AND2X1 U33 ( .IN1(n315), .IN2(n317), .Q(n310) );
  AND2X2 U34 ( .IN1(B[25]), .IN2(A[25]), .Q(n3) );
  NAND2X0 U35 ( .IN1(n179), .IN2(n354), .QN(n4) );
  NOR2X0 U36 ( .IN1(n374), .IN2(n375), .QN(n5) );
  OR2X1 U37 ( .IN1(B[8]), .IN2(A[8]), .Q(n6) );
  AND2X1 U38 ( .IN1(n179), .IN2(n349), .Q(n7) );
  AND2X1 U39 ( .IN1(n30), .IN2(n313), .Q(n8) );
  OR2X1 U40 ( .IN1(B[19]), .IN2(A[19]), .Q(n285) );
  OR2X1 U41 ( .IN1(B[3]), .IN2(A[3]), .Q(n368) );
  AND2X1 U42 ( .IN1(n278), .IN2(n279), .Q(n9) );
  AND2X1 U43 ( .IN1(n250), .IN2(n251), .Q(n10) );
  AND2X1 U44 ( .IN1(B[30]), .IN2(A[30]), .Q(n11) );
  NOR2X0 U45 ( .IN1(B[29]), .IN2(A[29]), .QN(n12) );
  OR2X1 U46 ( .IN1(n163), .IN2(n243), .Q(n13) );
  AND2X1 U47 ( .IN1(n335), .IN2(n71), .Q(n14) );
  AND2X4 U48 ( .IN1(n25), .IN2(n294), .Q(n15) );
  OR2X1 U49 ( .IN1(B[13]), .IN2(A[13]), .Q(n30) );
  NOR2X0 U50 ( .IN1(n123), .IN2(n120), .QN(n16) );
  OAI221X1 U51 ( .IN1(B[5]), .IN2(A[5]), .IN3(B[6]), .IN4(A[6]), .IN5(n22), 
        .QN(n57) );
  OR2X2 U52 ( .IN1(B[17]), .IN2(A[17]), .Q(n297) );
  NAND2X0 U53 ( .IN1(B[25]), .IN2(A[25]), .QN(n245) );
  INVX0 U54 ( .INP(n324), .ZN(n17) );
  INVX0 U55 ( .INP(n17), .ZN(n18) );
  OR2X1 U56 ( .IN1(B[10]), .IN2(A[10]), .Q(n324) );
  OR2X1 U57 ( .IN1(B[9]), .IN2(A[9]), .Q(n179) );
  NAND2X0 U58 ( .IN1(n313), .IN2(n325), .QN(n347) );
  NAND2X0 U59 ( .IN1(n353), .IN2(n18), .QN(n363) );
  AND2X1 U60 ( .IN1(n186), .IN2(n188), .Q(n19) );
  AND2X1 U61 ( .IN1(n299), .IN2(n297), .Q(n25) );
  INVX0 U62 ( .INP(n54), .ZN(n20) );
  XNOR3X1 U63 ( .IN1(n222), .IN2(A[30]), .IN3(n148), .Q(SUM[30]) );
  AND2X1 U64 ( .IN1(n106), .IN2(n270), .Q(n100) );
  NAND4X0 U65 ( .IN1(n352), .IN2(n351), .IN3(n353), .IN4(n180), .QN(n21) );
  AND2X1 U66 ( .IN1(B[4]), .IN2(A[4]), .Q(n22) );
  AND2X1 U67 ( .IN1(n205), .IN2(n368), .Q(n215) );
  AND2X1 U68 ( .IN1(n166), .IN2(n142), .Q(n143) );
  NOR2X0 U69 ( .IN1(B[13]), .IN2(A[13]), .QN(n23) );
  NAND2X0 U70 ( .IN1(n313), .IN2(n342), .QN(n24) );
  XNOR3X1 U71 ( .IN1(B[29]), .IN2(n227), .IN3(n225), .Q(SUM[29]) );
  NAND2X0 U72 ( .IN1(B[7]), .IN2(A[7]), .QN(n27) );
  OR2X1 U73 ( .IN1(n376), .IN2(n191), .Q(n29) );
  NAND4X0 U74 ( .IN1(n371), .IN2(n372), .IN3(n313), .IN4(n104), .QN(n333) );
  NAND2X0 U75 ( .IN1(n32), .IN2(n140), .QN(n31) );
  XOR2X1 U76 ( .IN1(n63), .IN2(n269), .Q(SUM[22]) );
  NOR2X0 U77 ( .IN1(n276), .IN2(n90), .QN(n32) );
  AND2X1 U78 ( .IN1(n224), .IN2(n220), .Q(n146) );
  AND4X1 U79 ( .IN1(n190), .IN2(n187), .IN3(n198), .IN4(n119), .Q(n65) );
  XOR3X1 U80 ( .IN1(A[13]), .IN2(n26), .IN3(n344), .Q(SUM[13]) );
  NAND2X0 U81 ( .IN1(n14), .IN2(n334), .QN(n332) );
  XOR3X1 U82 ( .IN1(A[25]), .IN2(B[25]), .IN3(n154), .Q(SUM[25]) );
  OA21X1 U83 ( .IN1(n193), .IN2(n194), .IN3(n28), .Q(n196) );
  AO21X1 U84 ( .IN1(n250), .IN2(n252), .IN3(n33), .Q(n256) );
  INVX0 U85 ( .INP(n255), .ZN(n33) );
  XOR3X1 U86 ( .IN1(A[15]), .IN2(B[15]), .IN3(n139), .Q(SUM[15]) );
  AO21X1 U87 ( .IN1(n280), .IN2(n9), .IN3(n34), .Q(n106) );
  INVX0 U88 ( .INP(n275), .ZN(n34) );
  AO22X2 U89 ( .IN1(B[25]), .IN2(A[25]), .IN3(B[24]), .IN4(A[24]), .Q(n122) );
  NAND4X0 U90 ( .IN1(n202), .IN2(n205), .IN3(n206), .IN4(n204), .QN(n183) );
  NAND2X0 U91 ( .IN1(n35), .IN2(n36), .QN(n56) );
  INVX0 U92 ( .INP(B[6]), .ZN(n35) );
  INVX0 U93 ( .INP(A[6]), .ZN(n36) );
  XOR3X1 U94 ( .IN1(A[26]), .IN2(B[26]), .IN3(n62), .Q(SUM[26]) );
  AO22X1 U95 ( .IN1(A[10]), .IN2(B[10]), .IN3(n359), .IN4(n18), .Q(n357) );
  AND3X1 U96 ( .IN1(n308), .IN2(n187), .IN3(n7), .Q(n171) );
  XOR3X1 U97 ( .IN1(A[14]), .IN2(B[14]), .IN3(n339), .Q(SUM[14]) );
  NAND2X0 U98 ( .IN1(n248), .IN2(n133), .QN(n154) );
  AND3X1 U99 ( .IN1(n240), .IN2(n157), .IN3(n13), .Q(n88) );
  AO21X1 U100 ( .IN1(n189), .IN2(n190), .IN3(n37), .Q(n184) );
  INVX0 U101 ( .INP(n188), .ZN(n37) );
  NAND3X0 U102 ( .IN1(n115), .IN2(n114), .IN3(n66), .QN(n160) );
  AO221X1 U103 ( .IN1(n91), .IN2(n277), .IN3(n264), .IN4(n124), .IN5(n38), .Q(
        n252) );
  INVX0 U104 ( .INP(n87), .ZN(n38) );
  AO222X1 U105 ( .IN1(n39), .IN2(n40), .IN3(n41), .IN4(n42), .IN5(n261), .IN6(
        n260), .Q(n249) );
  INVX0 U106 ( .INP(A[24]), .ZN(n39) );
  INVX0 U107 ( .INP(B[24]), .ZN(n40) );
  INVX0 U108 ( .INP(A[23]), .ZN(n41) );
  INVX0 U109 ( .INP(B[23]), .ZN(n42) );
  AO21X1 U110 ( .IN1(n343), .IN2(n108), .IN3(n43), .Q(n344) );
  INVX0 U111 ( .INP(n325), .ZN(n43) );
  AOI21X1 U112 ( .IN1(n44), .IN2(n264), .IN3(n283), .QN(n282) );
  INVX0 U113 ( .INP(n276), .ZN(n44) );
  AO21X1 U114 ( .IN1(n370), .IN2(n369), .IN3(n45), .Q(n200) );
  INVX0 U115 ( .INP(n205), .ZN(n45) );
  AO21X1 U116 ( .IN1(n249), .IN2(n248), .IN3(n46), .Q(n156) );
  INVX0 U117 ( .INP(n159), .ZN(n46) );
  AO22X2 U118 ( .IN1(n47), .IN2(n48), .IN3(n5), .IN4(n19), .Q(n109) );
  INVX0 U119 ( .INP(A[7]), .ZN(n47) );
  INVX0 U120 ( .INP(B[7]), .ZN(n48) );
  AO222X1 U121 ( .IN1(n227), .IN2(n226), .IN3(n239), .IN4(n238), .IN5(n96), 
        .IN6(n97), .Q(n151) );
  AO21X1 U122 ( .IN1(n85), .IN2(n61), .IN3(n138), .Q(n139) );
  MUX21X1 U123 ( .IN1(n241), .IN2(n79), .S(n170), .Q(SUM[27]) );
  AO22X1 U124 ( .IN1(n50), .IN2(n49), .IN3(n274), .IN4(n100), .Q(n63) );
  INVX0 U125 ( .INP(B[21]), .ZN(n49) );
  NAND2X0 U126 ( .IN1(n313), .IN2(n342), .QN(n107) );
  NAND2X0 U127 ( .IN1(n9), .IN2(n280), .QN(n277) );
  AOI21X1 U128 ( .IN1(n187), .IN2(n131), .IN3(n21), .QN(n345) );
  AOI21X1 U129 ( .IN1(n143), .IN2(n132), .IN3(n141), .QN(n77) );
  AO22X1 U130 ( .IN1(n49), .IN2(n50), .IN3(n51), .IN4(n52), .Q(n265) );
  INVX0 U131 ( .INP(A[21]), .ZN(n50) );
  INVX0 U132 ( .INP(B[22]), .ZN(n51) );
  INVX0 U133 ( .INP(A[22]), .ZN(n52) );
  AO221X1 U134 ( .IN1(n53), .IN2(n54), .IN3(n295), .IN4(n296), .IN5(n55), .Q(
        n128) );
  INVX0 U135 ( .INP(A[19]), .ZN(n53) );
  INVX0 U136 ( .INP(B[19]), .ZN(n54) );
  INVX0 U137 ( .INP(n294), .ZN(n55) );
  AND4X1 U138 ( .IN1(n318), .IN2(n306), .IN3(n307), .IN4(n319), .Q(n132) );
  AND2X1 U139 ( .IN1(n186), .IN2(n188), .Q(n373) );
  OA22X1 U140 ( .IN1(B[8]), .IN2(A[8]), .IN3(B[9]), .IN4(A[9]), .Q(n112) );
  AND3X1 U141 ( .IN1(n199), .IN2(n56), .IN3(n22), .Q(n374) );
  NAND3X0 U142 ( .IN1(n373), .IN2(n57), .IN3(n29), .QN(n78) );
  AOI21X1 U143 ( .IN1(n33), .IN2(n251), .IN3(n122), .QN(n137) );
  OA21X1 U144 ( .IN1(B[14]), .IN2(A[14]), .IN3(n314), .Q(n335) );
  NAND3X0 U145 ( .IN1(n58), .IN2(n59), .IN3(n364), .QN(n161) );
  INVX0 U146 ( .INP(n362), .ZN(n58) );
  AO21X1 U147 ( .IN1(n350), .IN2(n21), .IN3(n104), .Q(n342) );
  AND4X1 U148 ( .IN1(n318), .IN2(n307), .IN3(n306), .IN4(n319), .Q(n305) );
  AOI21X1 U149 ( .IN1(n64), .IN2(n15), .IN3(n284), .QN(n290) );
  NAND4X0 U150 ( .IN1(n320), .IN2(n317), .IN3(n321), .IN4(n118), .QN(n319) );
  INVX0 U151 ( .INP(n171), .ZN(n59) );
  NAND2X0 U152 ( .IN1(n88), .IN2(n156), .QN(n60) );
  OR2X1 U153 ( .IN1(n69), .IN2(n109), .Q(n68) );
  NAND2X0 U154 ( .IN1(n346), .IN2(n345), .QN(n61) );
  NAND2X0 U155 ( .IN1(n81), .IN2(n80), .QN(n62) );
  NAND2X0 U156 ( .IN1(n166), .IN2(n305), .QN(n64) );
  OR2X1 U157 ( .IN1(B[11]), .IN2(A[11]), .Q(n348) );
  AND2X1 U158 ( .IN1(B[8]), .IN2(A[8]), .Q(n354) );
  OR2X1 U159 ( .IN1(n3), .IN2(n247), .Q(n136) );
  NAND2X0 U160 ( .IN1(n21), .IN2(n350), .QN(n66) );
  AND2X1 U161 ( .IN1(n368), .IN2(n219), .Q(n369) );
  NAND2X0 U162 ( .IN1(n98), .IN2(n70), .QN(n67) );
  NAND2X0 U163 ( .IN1(n67), .IN2(n68), .QN(n177) );
  INVX0 U164 ( .INP(n6), .ZN(n69) );
  XOR2X1 U165 ( .IN1(n113), .IN2(n72), .Q(SUM[16]) );
  OR2X1 U166 ( .IN1(B[13]), .IN2(A[13]), .Q(n314) );
  OR2X1 U167 ( .IN1(n201), .IN2(n200), .Q(n73) );
  NAND2X0 U168 ( .IN1(n366), .IN2(n367), .QN(n74) );
  NOR2X0 U169 ( .IN1(n374), .IN2(n375), .QN(n75) );
  AND2X1 U170 ( .IN1(n10), .IN2(n136), .Q(n83) );
  NAND2X0 U171 ( .IN1(n93), .IN2(n92), .QN(n79) );
  NAND3X0 U172 ( .IN1(n135), .IN2(n342), .IN3(n8), .QN(n341) );
  OR2X1 U173 ( .IN1(B[12]), .IN2(A[12]), .Q(n313) );
  NAND2X0 U174 ( .IN1(n167), .IN2(n365), .QN(n98) );
  NAND2X0 U175 ( .IN1(n83), .IN2(n155), .QN(n80) );
  OR2X1 U176 ( .IN1(n137), .IN2(n82), .Q(n81) );
  INVX0 U177 ( .INP(n136), .ZN(n82) );
  NAND2X0 U178 ( .IN1(n366), .IN2(n367), .QN(n84) );
  NAND2X0 U179 ( .IN1(n366), .IN2(n367), .QN(n204) );
  NOR2X0 U180 ( .IN1(n107), .IN2(n337), .QN(n85) );
  AND2X1 U181 ( .IN1(n86), .IN2(n87), .Q(n260) );
  NAND2X0 U182 ( .IN1(n91), .IN2(n277), .QN(n86) );
  AND2X1 U183 ( .IN1(n266), .IN2(n267), .Q(n87) );
  AND2X1 U184 ( .IN1(n137), .IN2(n243), .Q(n95) );
  AND2X1 U185 ( .IN1(n198), .IN2(n119), .Q(n372) );
  NAND2X0 U186 ( .IN1(n88), .IN2(n156), .QN(n149) );
  AND2X1 U187 ( .IN1(n202), .IN2(n204), .Q(n167) );
  NOR2X0 U188 ( .IN1(n276), .IN2(n90), .QN(n89) );
  OR2X1 U189 ( .IN1(B[4]), .IN2(A[4]), .Q(n198) );
  INVX0 U190 ( .INP(n275), .ZN(n90) );
  NOR2X0 U191 ( .IN1(n265), .IN2(n34), .QN(n91) );
  NAND2X0 U192 ( .IN1(n95), .IN2(n133), .QN(n92) );
  AND2X1 U193 ( .IN1(n92), .IN2(n93), .Q(n241) );
  OR2X1 U194 ( .IN1(n94), .IN2(n110), .Q(n93) );
  NAND2X0 U195 ( .IN1(n159), .IN2(n246), .QN(n96) );
  AND2X1 U196 ( .IN1(n16), .IN2(n157), .Q(n97) );
  NAND3X0 U197 ( .IN1(n203), .IN2(n74), .IN3(n202), .QN(n201) );
  NAND2X0 U198 ( .IN1(n167), .IN2(n365), .QN(n99) );
  INVX0 U199 ( .INP(B[8]), .ZN(n101) );
  NAND2X0 U200 ( .IN1(n369), .IN2(n370), .QN(n102) );
  NAND2X0 U201 ( .IN1(n369), .IN2(n370), .QN(n206) );
  AND2X1 U202 ( .IN1(A[11]), .IN2(B[11]), .Q(n105) );
  AND3X1 U203 ( .IN1(n112), .IN2(n324), .IN3(n348), .Q(n104) );
  OR2X1 U204 ( .IN1(B[16]), .IN2(A[16]), .Q(n299) );
  INVX0 U205 ( .INP(n24), .ZN(n108) );
  NAND2X0 U206 ( .IN1(n299), .IN2(n297), .QN(n111) );
  NAND2X0 U207 ( .IN1(n166), .IN2(n132), .QN(n113) );
  NAND2X0 U208 ( .IN1(n98), .IN2(n116), .QN(n114) );
  OR2X1 U209 ( .IN1(n134), .IN2(n109), .Q(n115) );
  AND2X1 U210 ( .IN1(n65), .IN2(n117), .Q(n116) );
  INVX0 U211 ( .INP(n134), .ZN(n117) );
  NAND2X0 U212 ( .IN1(A[3]), .IN2(B[3]), .QN(n205) );
  AND3X1 U213 ( .IN1(n315), .IN2(n30), .IN3(n313), .Q(n118) );
  NAND2X0 U214 ( .IN1(n377), .IN2(n180), .QN(n362) );
  INVX0 U215 ( .INP(n240), .ZN(n120) );
  NOR2X0 U216 ( .IN1(B[14]), .IN2(A[14]), .QN(n121) );
  NOR2X0 U217 ( .IN1(n163), .IN2(n243), .QN(n123) );
  AND3X1 U218 ( .IN1(n89), .IN2(n262), .IN3(n263), .Q(n124) );
  AND2X1 U219 ( .IN1(n125), .IN2(n126), .Q(n318) );
  NAND2X0 U220 ( .IN1(n327), .IN2(n326), .QN(n125) );
  NAND2X0 U221 ( .IN1(n153), .IN2(n71), .QN(n126) );
  AND2X1 U222 ( .IN1(n234), .IN2(n127), .Q(n370) );
  AND2X1 U223 ( .IN1(B[0]), .IN2(A[0]), .Q(n127) );
  AND2X1 U224 ( .IN1(n129), .IN2(n128), .Q(n280) );
  OR2X1 U225 ( .IN1(n165), .IN2(n292), .Q(n129) );
  NAND2X0 U226 ( .IN1(n144), .IN2(n145), .QN(n130) );
  AND2X1 U227 ( .IN1(n206), .IN2(n205), .Q(n365) );
  NAND2X0 U228 ( .IN1(n19), .IN2(n5), .QN(n131) );
  NAND2X0 U229 ( .IN1(n19), .IN2(n75), .QN(n308) );
  NAND2X0 U230 ( .IN1(n10), .IN2(n252), .QN(n133) );
  INVX0 U231 ( .INP(n104), .ZN(n134) );
  NAND2X0 U232 ( .IN1(n345), .IN2(n178), .QN(n135) );
  NAND2X0 U233 ( .IN1(A[13]), .IN2(B[13]), .QN(n338) );
  NAND2X0 U234 ( .IN1(n336), .IN2(n331), .QN(n138) );
  NAND2X0 U235 ( .IN1(A[14]), .IN2(B[14]), .QN(n331) );
  AND2X1 U236 ( .IN1(n368), .IN2(n219), .Q(n366) );
  NAND2X0 U237 ( .IN1(n313), .IN2(n30), .QN(n312) );
  NAND2X0 U238 ( .IN1(n166), .IN2(n132), .QN(n140) );
  NAND2X0 U239 ( .IN1(n166), .IN2(n305), .QN(n264) );
  INVX0 U240 ( .INP(n293), .ZN(n142) );
  NAND2X0 U241 ( .IN1(n103), .IN2(n151), .QN(n144) );
  OR2X1 U242 ( .IN1(n11), .IN2(n221), .Q(n145) );
  AND2X1 U243 ( .IN1(n224), .IN2(n152), .Q(n147) );
  OR2X1 U244 ( .IN1(n12), .IN2(n235), .Q(n152) );
  OR2X4 U245 ( .IN1(B[6]), .IN2(A[6]), .Q(n190) );
  NAND2X0 U246 ( .IN1(n147), .IN2(n151), .QN(n148) );
  NOR3X0 U247 ( .IN1(n121), .IN2(n23), .IN3(n325), .QN(n153) );
  NAND2X0 U248 ( .IN1(n124), .IN2(n64), .QN(n261) );
  INVX0 U249 ( .INP(n119), .ZN(n209) );
  AND2X1 U250 ( .IN1(n247), .IN2(n164), .Q(n159) );
  OR2X1 U251 ( .IN1(n158), .IN2(n245), .Q(n157) );
  NAND2X0 U252 ( .IN1(n260), .IN2(n261), .QN(n155) );
  AND2X1 U253 ( .IN1(n242), .IN2(n244), .Q(n164) );
  OR2X1 U254 ( .IN1(B[14]), .IN2(A[14]), .Q(n315) );
  INVX0 U255 ( .INP(n164), .ZN(n158) );
  NAND2X0 U256 ( .IN1(n275), .IN2(n279), .QN(n281) );
  NAND2X0 U257 ( .IN1(n255), .IN2(n250), .QN(n259) );
  NAND2X0 U258 ( .IN1(n285), .IN2(n278), .QN(n289) );
  XNOR2X1 U259 ( .IN1(n161), .IN2(n363), .Q(SUM[10]) );
  NAND2X0 U260 ( .IN1(n198), .IN2(n119), .QN(n194) );
  NAND2X0 U261 ( .IN1(n222), .IN2(n223), .QN(n221) );
  NAND2X0 U262 ( .IN1(n20), .IN2(A[19]), .QN(n278) );
  NAND2X0 U263 ( .IN1(B[18]), .IN2(A[18]), .QN(n292) );
  NAND2X0 U264 ( .IN1(B[20]), .IN2(A[20]), .QN(n279) );
  NAND2X0 U265 ( .IN1(B[22]), .IN2(A[22]), .QN(n267) );
  NAND2X0 U266 ( .IN1(B[21]), .IN2(A[21]), .QN(n270) );
  NAND2X0 U267 ( .IN1(B[23]), .IN2(A[23]), .QN(n255) );
  AND2X1 U268 ( .IN1(n288), .IN2(n287), .Q(SUM[0]) );
  NAND2X0 U269 ( .IN1(B[27]), .IN2(A[27]), .QN(n240) );
  INVX0 U270 ( .INP(n242), .ZN(n163) );
  NOR2X0 U271 ( .IN1(B[19]), .IN2(A[19]), .QN(n165) );
  NAND2X0 U272 ( .IN1(n31), .IN2(n106), .QN(n271) );
  AND2X1 U273 ( .IN1(n7), .IN2(n65), .Q(n168) );
  INVX0 U274 ( .INP(n348), .ZN(n322) );
  INVX0 U275 ( .INP(n270), .ZN(n268) );
  NOR2X0 U276 ( .IN1(n356), .IN2(n322), .QN(n350) );
  AND2X1 U277 ( .IN1(n190), .IN2(n187), .Q(n371) );
  NAND2X0 U278 ( .IN1(n372), .IN2(n73), .QN(n192) );
  NOR2X0 U279 ( .IN1(n177), .IN2(n173), .QN(n176) );
  NOR2X0 U280 ( .IN1(n302), .IN2(n303), .QN(n301) );
  NOR2X0 U281 ( .IN1(n268), .IN2(n273), .QN(n272) );
  INVX0 U282 ( .INP(n263), .ZN(n273) );
  NOR2X0 U283 ( .IN1(n174), .IN2(n254), .QN(n257) );
  OR2X1 U284 ( .IN1(n169), .IN2(n337), .Q(n336) );
  AND2X1 U285 ( .IN1(n325), .IN2(n338), .Q(n169) );
  INVX0 U286 ( .INP(n198), .ZN(n213) );
  NAND2X0 U287 ( .IN1(n280), .IN2(n278), .QN(n283) );
  NOR2X0 U288 ( .IN1(n212), .IN2(n213), .QN(n211) );
  INVX0 U289 ( .INP(B[29]), .ZN(n226) );
  INVX0 U290 ( .INP(B[28]), .ZN(n238) );
  AND2X1 U291 ( .IN1(n338), .IN2(n172), .Q(n340) );
  OR2X1 U292 ( .IN1(n23), .IN2(n325), .Q(n172) );
  INVX0 U293 ( .INP(n287), .ZN(n233) );
  INVX0 U294 ( .INP(B[30]), .ZN(n222) );
  INVX0 U295 ( .INP(n297), .ZN(n303) );
  XNOR2X1 U296 ( .IN1(n286), .IN2(n233), .Q(SUM[1]) );
  NAND2X0 U297 ( .IN1(B[29]), .IN2(A[29]), .QN(n224) );
  NAND2X0 U298 ( .IN1(B[28]), .IN2(A[28]), .QN(n235) );
  NAND2X0 U299 ( .IN1(n238), .IN2(n239), .QN(n237) );
  OR2X1 U300 ( .IN1(B[5]), .IN2(A[5]), .Q(n199) );
  NAND2X0 U301 ( .IN1(B[30]), .IN2(A[30]), .QN(n220) );
  OR2X1 U302 ( .IN1(B[20]), .IN2(A[20]), .Q(n275) );
  OR2X1 U303 ( .IN1(B[24]), .IN2(A[24]), .Q(n251) );
  NAND2X0 U304 ( .IN1(A[11]), .IN2(B[11]), .QN(n352) );
  NAND2X1 U305 ( .IN1(B[12]), .IN2(A[12]), .QN(n325) );
  OR2X1 U306 ( .IN1(B[2]), .IN2(A[2]), .Q(n219) );
  NAND2X0 U307 ( .IN1(B[0]), .IN2(A[0]), .QN(n287) );
  OR2X1 U308 ( .IN1(B[21]), .IN2(A[21]), .Q(n263) );
  NAND2X0 U309 ( .IN1(B[10]), .IN2(A[10]), .QN(n353) );
  NAND2X1 U310 ( .IN1(B[26]), .IN2(A[26]), .QN(n243) );
  OR2X1 U311 ( .IN1(B[18]), .IN2(A[18]), .Q(n294) );
  OR2X1 U312 ( .IN1(B[25]), .IN2(A[25]), .Q(n247) );
  OR2X1 U313 ( .IN1(B[22]), .IN2(A[22]), .Q(n262) );
  OR2X1 U314 ( .IN1(B[1]), .IN2(A[1]), .Q(n234) );
  AND2X1 U315 ( .IN1(B[24]), .IN2(A[24]), .Q(n174) );
  OR2X1 U316 ( .IN1(B[27]), .IN2(A[27]), .Q(n242) );
  OR2X1 U317 ( .IN1(B[26]), .IN2(A[26]), .Q(n244) );
  OR2X1 U318 ( .IN1(B[23]), .IN2(A[23]), .Q(n250) );
  INVX0 U319 ( .INP(A[15]), .ZN(n328) );
  INVX0 U320 ( .INP(A[28]), .ZN(n239) );
  INVX0 U321 ( .INP(A[29]), .ZN(n227) );
  NAND2X0 U322 ( .IN1(n378), .IN2(n379), .QN(n288) );
  INVX0 U323 ( .INP(A[0]), .ZN(n379) );
  INVX0 U324 ( .INP(B[0]), .ZN(n378) );
  INVX0 U325 ( .INP(A[30]), .ZN(n223) );
  NAND2X0 U326 ( .IN1(n328), .IN2(n329), .QN(n327) );
  NAND2X0 U327 ( .IN1(n236), .IN2(n235), .QN(n225) );
  INVX0 U328 ( .INP(n155), .ZN(n258) );
  NAND2X0 U329 ( .IN1(n340), .IN2(n341), .QN(n339) );
  INVX0 U330 ( .INP(A[8]), .ZN(n355) );
  NAND2X0 U331 ( .IN1(B[9]), .IN2(A[9]), .QN(n180) );
  NAND2X0 U332 ( .IN1(A[17]), .IN2(B[17]), .QN(n296) );
  NAND2X0 U333 ( .IN1(A[1]), .IN2(B[1]), .QN(n231) );
  NAND2X0 U334 ( .IN1(B[16]), .IN2(A[16]), .QN(n298) );
  NAND2X0 U335 ( .IN1(B[7]), .IN2(A[7]), .QN(n186) );
  NAND2X0 U336 ( .IN1(n216), .IN2(n217), .QN(n214) );
  INVX0 U337 ( .INP(n216), .ZN(n229) );
  INVX0 U338 ( .INP(n338), .ZN(n316) );
  INVX0 U339 ( .INP(n296), .ZN(n302) );
  NAND2X0 U340 ( .IN1(n296), .IN2(n295), .QN(n293) );
  NAND2X0 U341 ( .IN1(n203), .IN2(n210), .QN(n207) );
  INVX0 U342 ( .INP(n203), .ZN(n212) );
  NAND2X0 U343 ( .IN1(n28), .IN2(n192), .QN(n189) );
  INVX0 U344 ( .INP(n28), .ZN(n197) );
  NOR2X0 U345 ( .IN1(n376), .IN2(n191), .QN(n375) );
  NAND2X0 U346 ( .IN1(n231), .IN2(n232), .QN(n218) );
  INVX0 U347 ( .INP(n231), .ZN(n367) );
  NAND2X0 U348 ( .IN1(n27), .IN2(n187), .QN(n185) );
  NAND2X0 U349 ( .IN1(n330), .IN2(n331), .QN(n326) );
  NAND2X0 U350 ( .IN1(A[15]), .IN2(B[15]), .QN(n330) );
  NAND2X0 U351 ( .IN1(n30), .IN2(n315), .QN(n337) );
  NAND2X0 U352 ( .IN1(n229), .IN2(n368), .QN(n202) );
  NAND2X0 U353 ( .IN1(n267), .IN2(n262), .QN(n269) );
  NAND2X0 U354 ( .IN1(n268), .IN2(n262), .QN(n266) );
  NAND2X0 U355 ( .IN1(n101), .IN2(n355), .QN(n349) );
  NAND2X0 U356 ( .IN1(n218), .IN2(n219), .QN(n217) );
  NAND2X0 U357 ( .IN1(A[4]), .IN2(B[4]), .QN(n203) );
  NAND2X0 U358 ( .IN1(n248), .IN2(n249), .QN(n246) );
  NOR2X0 U359 ( .IN1(n253), .IN2(n174), .QN(n248) );
  NAND2X0 U360 ( .IN1(n190), .IN2(n188), .QN(n195) );
  NAND2X0 U361 ( .IN1(A[6]), .IN2(B[6]), .QN(n188) );
  NOR2X0 U362 ( .IN1(B[6]), .IN2(A[6]), .QN(n376) );
  NOR2X0 U363 ( .IN1(n171), .IN2(n362), .QN(n360) );
  NOR2X0 U364 ( .IN1(n197), .IN2(n209), .QN(n208) );
  INVX0 U365 ( .INP(n219), .ZN(n230) );
  NAND2X0 U366 ( .IN1(n179), .IN2(n354), .QN(n351) );
  NAND2X0 U367 ( .IN1(n173), .IN2(n179), .QN(n377) );
  NAND2X0 U368 ( .IN1(n179), .IN2(n180), .QN(n175) );
  NAND2X0 U369 ( .IN1(n361), .IN2(n360), .QN(n359) );
  NAND2X0 U370 ( .IN1(n109), .IN2(n178), .QN(n181) );
  INVX0 U371 ( .INP(B[15]), .ZN(n329) );
  NAND4X0 U372 ( .IN1(n84), .IN2(n102), .IN3(n202), .IN4(n205), .QN(n334) );
  NOR2X0 U373 ( .IN1(n173), .IN2(n69), .QN(n182) );
  NAND2X1 U374 ( .IN1(n291), .IN2(n292), .QN(n284) );
  NOR2X0 U375 ( .IN1(n229), .IN2(n230), .QN(n228) );
  NAND2X0 U376 ( .IN1(A[2]), .IN2(B[2]), .QN(n216) );
  NAND2X0 U377 ( .IN1(n293), .IN2(n294), .QN(n291) );
  NAND2X0 U378 ( .IN1(n233), .IN2(n234), .QN(n232) );
  NAND2X0 U379 ( .IN1(n234), .IN2(n231), .QN(n286) );
  NOR2X0 U380 ( .IN1(n201), .IN2(n200), .QN(n193) );
  INVX0 U381 ( .INP(n251), .ZN(n254) );
  NOR2X0 U382 ( .IN1(n254), .IN2(n255), .QN(n253) );
  NOR2X0 U383 ( .IN1(n322), .IN2(n105), .QN(n358) );
  NOR2X0 U384 ( .IN1(n105), .IN2(n324), .QN(n356) );
  NOR2X0 U385 ( .IN1(n322), .IN2(n323), .QN(n320) );
  NOR2X0 U386 ( .IN1(n105), .IN2(n324), .QN(n323) );
  NAND2X0 U387 ( .IN1(n150), .IN2(n297), .QN(n295) );
  NAND2X0 U388 ( .IN1(n346), .IN2(n345), .QN(n343) );
  NAND2X0 U389 ( .IN1(n298), .IN2(n304), .QN(n300) );
  NAND2X0 U390 ( .IN1(n299), .IN2(n113), .QN(n304) );
  NAND2X0 U391 ( .IN1(n32), .IN2(n140), .QN(n274) );
  NOR2X0 U392 ( .IN1(n311), .IN2(n312), .QN(n309) );
  NAND2X0 U393 ( .IN1(n168), .IN2(n99), .QN(n364) );
  NAND2X0 U394 ( .IN1(n198), .IN2(n99), .QN(n210) );
  NAND2X0 U395 ( .IN1(n168), .IN2(n99), .QN(n361) );
  NAND2X0 U396 ( .IN1(n65), .IN2(n183), .QN(n178) );
  NAND2X0 U397 ( .IN1(n65), .IN2(n183), .QN(n346) );
  NAND2X0 U398 ( .IN1(n237), .IN2(n149), .QN(n236) );
  XOR2X1 U399 ( .IN1(n175), .IN2(n176), .Q(SUM[9]) );
  XOR2X1 U400 ( .IN1(n181), .IN2(n182), .Q(SUM[8]) );
  XOR2X1 U401 ( .IN1(n195), .IN2(n196), .Q(SUM[6]) );
  XOR2X1 U402 ( .IN1(n207), .IN2(n208), .Q(SUM[5]) );
  XOR2X1 U403 ( .IN1(n214), .IN2(n215), .Q(SUM[3]) );
  XOR2X1 U404 ( .IN1(n218), .IN2(n228), .Q(SUM[2]) );
  XOR2X1 U405 ( .IN1(n258), .IN2(n259), .Q(SUM[23]) );
  XOR2X1 U406 ( .IN1(n281), .IN2(n282), .Q(SUM[20]) );
  XOR2X1 U407 ( .IN1(n289), .IN2(n290), .Q(SUM[19]) );
  XOR2X1 U408 ( .IN1(n300), .IN2(n301), .Q(SUM[17]) );
  NAND4X0 U409 ( .IN1(n309), .IN2(n78), .IN3(n310), .IN4(n187), .QN(n307) );
  NAND3X0 U410 ( .IN1(n112), .IN2(n324), .IN3(n348), .QN(n311) );
  NAND4X0 U411 ( .IN1(n352), .IN2(n4), .IN3(n353), .IN4(n180), .QN(n321) );
endmodule


module SeqMult_DW01_sub_9 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115;

  OR2X4 U3 ( .IN1(n59), .IN2(n29), .Q(n58) );
  INVX0 U4 ( .INP(B[28]), .ZN(n81) );
  AND2X1 U5 ( .IN1(n90), .IN2(n91), .Q(n28) );
  NOR4X0 U6 ( .IN1(B[11]), .IN2(B[10]), .IN3(B[12]), .IN4(B[13]), .QN(n96) );
  AND2X1 U7 ( .IN1(n50), .IN2(n83), .Q(n49) );
  AND2X1 U8 ( .IN1(n41), .IN2(n87), .Q(n45) );
  NOR2X0 U9 ( .IN1(B[17]), .IN2(B[16]), .QN(n93) );
  AND2X1 U10 ( .IN1(n112), .IN2(n113), .Q(n38) );
  XOR2X1 U11 ( .IN1(n50), .IN2(n83), .Q(DIFF[26]) );
  XOR2X1 U12 ( .IN1(n45), .IN2(n86), .Q(DIFF[23]) );
  XOR2X1 U13 ( .IN1(n41), .IN2(n87), .Q(DIFF[22]) );
  XOR2X1 U14 ( .IN1(n43), .IN2(n88), .Q(DIFF[21]) );
  XOR2X1 U15 ( .IN1(n42), .IN2(n90), .Q(DIFF[18]) );
  NAND4X0 U16 ( .IN1(n3), .IN2(n11), .IN3(n57), .IN4(n24), .QN(n111) );
  AND2X1 U17 ( .IN1(n103), .IN2(n7), .Q(n24) );
  OR2X1 U18 ( .IN1(n53), .IN2(n29), .Q(n61) );
  NAND3X1 U19 ( .IN1(n16), .IN2(n74), .IN3(n15), .QN(n72) );
  XNOR2X1 U20 ( .IN1(n16), .IN2(DIFF[0]), .Q(DIFF[1]) );
  INVX0 U21 ( .INP(B[9]), .ZN(n1) );
  NOR2X0 U22 ( .IN1(n23), .IN2(B[25]), .QN(n2) );
  XOR2X1 U23 ( .IN1(n104), .IN2(n108), .Q(DIFF[12]) );
  AND2X1 U24 ( .IN1(n40), .IN2(n93), .Q(n42) );
  AND4X1 U25 ( .IN1(n14), .IN2(n74), .IN3(n15), .IN4(n73), .Q(n3) );
  XNOR2X1 U26 ( .IN1(n6), .IN2(n71), .Q(DIFF[4]) );
  INVX0 U27 ( .INP(n6), .ZN(n4) );
  INVX0 U28 ( .INP(n107), .ZN(n5) );
  INVX0 U29 ( .INP(n68), .ZN(n6) );
  INVX0 U30 ( .INP(B[9]), .ZN(n7) );
  INVX0 U31 ( .INP(n66), .ZN(n62) );
  INVX0 U32 ( .INP(n60), .ZN(n8) );
  INVX0 U33 ( .INP(n8), .ZN(n9) );
  INVX0 U34 ( .INP(B[6]), .ZN(n10) );
  NAND4X0 U35 ( .IN1(n104), .IN2(n5), .IN3(n38), .IN4(n18), .QN(n106) );
  INVX0 U36 ( .INP(n59), .ZN(n11) );
  INVX0 U37 ( .INP(B[8]), .ZN(n12) );
  AND3X1 U38 ( .IN1(n40), .IN2(n93), .IN3(n90), .Q(n13) );
  INVX0 U39 ( .INP(n13), .ZN(n92) );
  INVX0 U40 ( .INP(B[3]), .ZN(n14) );
  INVX0 U41 ( .INP(B[0]), .ZN(n15) );
  INVX0 U42 ( .INP(B[1]), .ZN(n16) );
  AND4X1 U43 ( .IN1(n39), .IN2(n65), .IN3(n60), .IN4(n10), .Q(n98) );
  AND4X1 U44 ( .IN1(n74), .IN2(n14), .IN3(n73), .IN4(n80), .Q(n99) );
  AND4X1 U45 ( .IN1(n1), .IN2(n57), .IN3(n100), .IN4(n101), .Q(n97) );
  OR2X1 U46 ( .IN1(n34), .IN2(n29), .Q(n56) );
  NAND2X0 U47 ( .IN1(n31), .IN2(n105), .QN(n19) );
  AND2X1 U48 ( .IN1(n41), .IN2(n17), .Q(n50) );
  AND2X1 U49 ( .IN1(n2), .IN2(n87), .Q(n17) );
  AND2X4 U50 ( .IN1(n105), .IN2(n100), .Q(n18) );
  XOR2X1 U51 ( .IN1(n103), .IN2(n47), .Q(DIFF[10]) );
  XOR2X1 U52 ( .IN1(B[14]), .IN2(n19), .Q(DIFF[14]) );
  AND3X1 U53 ( .IN1(n37), .IN2(n38), .IN3(n104), .Q(n20) );
  XOR2X1 U54 ( .IN1(n84), .IN2(n51), .Q(DIFF[25]) );
  AND4X1 U55 ( .IN1(n99), .IN2(n98), .IN3(n97), .IN4(n96), .Q(n35) );
  INVX0 U56 ( .INP(n80), .ZN(DIFF[0]) );
  NOR2X0 U57 ( .IN1(n22), .IN2(n23), .QN(n51) );
  NAND2X0 U58 ( .IN1(n41), .IN2(n87), .QN(n22) );
  NAND2X1 U59 ( .IN1(n85), .IN2(n86), .QN(n23) );
  XOR2X1 U60 ( .IN1(n20), .IN2(n105), .Q(DIFF[13]) );
  XOR2X1 U61 ( .IN1(n66), .IN2(n70), .Q(DIFF[5]) );
  XOR2X2 U62 ( .IN1(n35), .IN2(n94), .Q(DIFF[16]) );
  NAND2X1 U63 ( .IN1(n113), .IN2(n112), .QN(n29) );
  OR2X1 U64 ( .IN1(n52), .IN2(n29), .Q(n67) );
  AND2X1 U65 ( .IN1(n44), .IN2(n25), .Q(n41) );
  AND2X1 U66 ( .IN1(n89), .IN2(n88), .Q(n25) );
  AND2X1 U67 ( .IN1(n42), .IN2(n28), .Q(n44) );
  AND2X1 U68 ( .IN1(n26), .IN2(n27), .Q(n110) );
  NOR2X0 U69 ( .IN1(B[9]), .IN2(B[8]), .QN(n26) );
  NOR2X0 U70 ( .IN1(B[11]), .IN2(B[10]), .QN(n27) );
  NOR2X0 U71 ( .IN1(n59), .IN2(B[8]), .QN(n30) );
  AND3X1 U72 ( .IN1(n37), .IN2(n38), .IN3(n104), .Q(n31) );
  AND2X1 U73 ( .IN1(n49), .IN2(n82), .Q(n48) );
  AND2X1 U74 ( .IN1(n3), .IN2(n30), .Q(n32) );
  AND2X1 U75 ( .IN1(n50), .IN2(n83), .Q(n33) );
  NAND2X0 U76 ( .IN1(n12), .IN2(n36), .QN(n34) );
  NOR2X0 U77 ( .IN1(B[3]), .IN2(B[2]), .QN(n113) );
  AND2X1 U78 ( .IN1(n36), .IN2(n110), .Q(n37) );
  NOR2X0 U79 ( .IN1(B[5]), .IN2(B[6]), .QN(n115) );
  AND2X1 U80 ( .IN1(n114), .IN2(n115), .Q(n36) );
  INVX0 U81 ( .INP(B[5]), .ZN(n39) );
  XNOR2X1 U82 ( .IN1(n106), .IN2(n101), .Q(DIFF[15]) );
  XNOR2X1 U83 ( .IN1(n111), .IN2(n102), .Q(DIFF[11]) );
  XNOR2X1 U84 ( .IN1(n56), .IN2(n7), .Q(DIFF[9]) );
  XNOR2X1 U85 ( .IN1(n67), .IN2(n64), .Q(DIFF[6]) );
  XNOR2X1 U86 ( .IN1(n58), .IN2(n12), .Q(DIFF[8]) );
  XNOR2X1 U87 ( .IN1(n61), .IN2(n9), .Q(DIFF[7]) );
  XNOR2X1 U88 ( .IN1(n72), .IN2(n14), .Q(DIFF[3]) );
  AND4X1 U89 ( .IN1(n99), .IN2(n97), .IN3(n98), .IN4(n96), .Q(n40) );
  INVX0 U90 ( .INP(n38), .ZN(n109) );
  AND2X1 U91 ( .IN1(n44), .IN2(n89), .Q(n43) );
  XOR2X1 U92 ( .IN1(n46), .IN2(n85), .Q(DIFF[24]) );
  NOR2X0 U93 ( .IN1(n71), .IN2(n4), .QN(n70) );
  INVX0 U94 ( .INP(n74), .ZN(n78) );
  AND2X1 U95 ( .IN1(n45), .IN2(n86), .Q(n46) );
  AND2X1 U96 ( .IN1(n32), .IN2(n7), .Q(n47) );
  INVX0 U97 ( .INP(n65), .ZN(n68) );
  XOR2X1 U98 ( .IN1(B[19]), .IN2(n92), .Q(DIFF[19]) );
  XOR2X1 U99 ( .IN1(n79), .IN2(n78), .Q(DIFF[2]) );
  XOR2X1 U100 ( .IN1(B[17]), .IN2(n95), .Q(DIFF[17]) );
  XOR2X1 U101 ( .IN1(n89), .IN2(n44), .Q(DIFF[20]) );
  OR2X1 U102 ( .IN1(n68), .IN2(n69), .Q(n52) );
  OR2X1 U103 ( .IN1(n63), .IN2(n62), .Q(n53) );
  XOR2X1 U104 ( .IN1(n33), .IN2(n82), .Q(DIFF[27]) );
  INVX0 U105 ( .INP(B[5]), .ZN(n66) );
  INVX0 U106 ( .INP(B[1]), .ZN(n73) );
  INVX0 U107 ( .INP(B[6]), .ZN(n64) );
  INVX0 U108 ( .INP(B[7]), .ZN(n60) );
  INVX0 U109 ( .INP(B[2]), .ZN(n74) );
  INVX0 U110 ( .INP(B[0]), .ZN(n80) );
  INVX0 U111 ( .INP(B[12]), .ZN(n104) );
  AND2X1 U112 ( .IN1(n81), .IN2(n48), .Q(n54) );
  INVX0 U113 ( .INP(B[13]), .ZN(n105) );
  INVX0 U114 ( .INP(B[4]), .ZN(n65) );
  AND2X1 U115 ( .IN1(n77), .IN2(n54), .Q(n55) );
  INVX0 U116 ( .INP(B[16]), .ZN(n94) );
  INVX0 U117 ( .INP(B[8]), .ZN(n57) );
  INVX0 U118 ( .INP(B[10]), .ZN(n103) );
  INVX0 U119 ( .INP(B[18]), .ZN(n90) );
  INVX0 U120 ( .INP(B[29]), .ZN(n77) );
  XNOR2X1 U121 ( .IN1(n48), .IN2(B[28]), .Q(DIFF[28]) );
  XNOR2X1 U122 ( .IN1(n55), .IN2(B[30]), .Q(DIFF[30]) );
  INVX0 U123 ( .INP(B[11]), .ZN(n102) );
  XOR2X1 U124 ( .IN1(B[31]), .IN2(n75), .Q(DIFF[31]) );
  NAND2X0 U125 ( .IN1(n76), .IN2(n55), .QN(n75) );
  INVX0 U126 ( .INP(B[14]), .ZN(n100) );
  INVX0 U127 ( .INP(B[19]), .ZN(n91) );
  INVX0 U128 ( .INP(B[15]), .ZN(n101) );
  INVX0 U129 ( .INP(B[21]), .ZN(n88) );
  INVX0 U130 ( .INP(B[20]), .ZN(n89) );
  INVX0 U131 ( .INP(B[22]), .ZN(n87) );
  INVX0 U132 ( .INP(B[23]), .ZN(n86) );
  INVX0 U133 ( .INP(B[24]), .ZN(n85) );
  INVX0 U134 ( .INP(B[25]), .ZN(n84) );
  INVX0 U135 ( .INP(B[26]), .ZN(n83) );
  INVX0 U136 ( .INP(B[27]), .ZN(n82) );
  INVX0 U137 ( .INP(B[30]), .ZN(n76) );
  XOR2X1 U138 ( .IN1(n54), .IN2(n77), .Q(DIFF[29]) );
  INVX0 U139 ( .INP(n3), .ZN(n71) );
  NOR2X0 U140 ( .IN1(B[0]), .IN2(B[1]), .QN(n112) );
  NAND2X0 U141 ( .IN1(n114), .IN2(n115), .QN(n59) );
  NAND2X0 U142 ( .IN1(n35), .IN2(n94), .QN(n95) );
  NAND2X0 U143 ( .IN1(n15), .IN2(n16), .QN(n79) );
  NAND2X0 U144 ( .IN1(n64), .IN2(n65), .QN(n63) );
  NAND2X0 U145 ( .IN1(n110), .IN2(n36), .QN(n107) );
  NOR2X0 U146 ( .IN1(n109), .IN2(n107), .QN(n108) );
  NOR2X0 U147 ( .IN1(B[4]), .IN2(B[7]), .QN(n114) );
  INVX0 U148 ( .INP(n39), .ZN(n69) );
endmodule


module SeqMult ( clk, internalClk, rst, A, B, P );
  input [31:0] A;
  input [31:0] B;
  output [63:0] P;
  input clk, internalClk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N76, N77, N78, N79, N80, N81,
         N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95,
         N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107,
         N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151,
         N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162,
         N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261,
         N263, N264, N265, N266, N267, N268, N303, N304, N305, N306, N307,
         N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318,
         N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329,
         N330, N331, N332, N333, N334, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N465, N466, N467, N468, N469, N470, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483,
         N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494,
         N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505,
         N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516,
         N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527,
         N528, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542,
         N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553,
         N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564,
         N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575,
         N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586,
         N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N829,
         N831, N833, N835, N837, N839, N841, N843, N845, N847, N849, N851,
         N853, N855, N857, N859, N861, N863, N865, N867, N869, N871, N873,
         N875, N877, N879, N881, N883, N885, N887, N889, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n368,
         n370, n372, n376, n378, n380, n382, n384, n386, n388, n390, n392,
         n394, n396, n398, n399, n401, n402, n403, n404, n405, n406, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, N697, N696, N695, N694, N693, N692, N691, N690, N689,
         N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678,
         N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667,
         N666, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054;
  wire   [31:0] counter;
  wire   [31:0] A_reg;
  wire   [31:0] B_reg;
  wire   SYNOPSYS_UNCONNECTED__0;

  DFFX1 \A_reg_reg[31]  ( .D(N40), .CLK(clk), .Q(A_reg[31]), .QN(n399) );
  DFFX1 \A_reg_reg[30]  ( .D(N39), .CLK(clk), .Q(A_reg[30]) );
  DFFX1 \A_reg_reg[29]  ( .D(N38), .CLK(clk), .Q(A_reg[29]) );
  DFFX1 \A_reg_reg[28]  ( .D(N37), .CLK(clk), .Q(A_reg[28]) );
  DFFX1 \A_reg_reg[27]  ( .D(N36), .CLK(clk), .Q(A_reg[27]) );
  DFFX1 \A_reg_reg[26]  ( .D(N35), .CLK(clk), .Q(A_reg[26]) );
  DFFX1 \A_reg_reg[25]  ( .D(N34), .CLK(clk), .Q(A_reg[25]) );
  DFFX1 \A_reg_reg[24]  ( .D(N33), .CLK(clk), .Q(A_reg[24]) );
  DFFX1 \A_reg_reg[23]  ( .D(N32), .CLK(clk), .Q(A_reg[23]) );
  DFFX1 \A_reg_reg[22]  ( .D(N31), .CLK(clk), .Q(A_reg[22]) );
  DFFX1 \A_reg_reg[21]  ( .D(N30), .CLK(clk), .Q(A_reg[21]) );
  DFFX1 \A_reg_reg[20]  ( .D(N29), .CLK(clk), .Q(A_reg[20]) );
  DFFX1 \A_reg_reg[19]  ( .D(N28), .CLK(clk), .Q(A_reg[19]) );
  DFFX1 \A_reg_reg[18]  ( .D(N27), .CLK(clk), .Q(A_reg[18]) );
  DFFX1 \A_reg_reg[17]  ( .D(N26), .CLK(clk), .Q(A_reg[17]) );
  DFFX1 \A_reg_reg[16]  ( .D(N25), .CLK(clk), .Q(A_reg[16]) );
  DFFX1 \A_reg_reg[15]  ( .D(N24), .CLK(clk), .Q(A_reg[15]), .QN(n368) );
  DFFX1 \A_reg_reg[14]  ( .D(N23), .CLK(clk), .Q(A_reg[14]), .QN(n370) );
  DFFX1 \A_reg_reg[13]  ( .D(N22), .CLK(clk), .Q(A_reg[13]), .QN(n372) );
  DFFX1 \A_reg_reg[12]  ( .D(N21), .CLK(clk), .Q(A_reg[12]) );
  DFFX1 \A_reg_reg[11]  ( .D(N20), .CLK(clk), .Q(A_reg[11]), .QN(n376) );
  DFFX1 \A_reg_reg[10]  ( .D(N19), .CLK(clk), .Q(A_reg[10]), .QN(n378) );
  DFFX1 \A_reg_reg[9]  ( .D(N18), .CLK(clk), .Q(A_reg[9]), .QN(n380) );
  DFFX1 \A_reg_reg[8]  ( .D(N17), .CLK(clk), .Q(A_reg[8]), .QN(n382) );
  DFFX1 \A_reg_reg[7]  ( .D(N16), .CLK(clk), .Q(A_reg[7]), .QN(n384) );
  DFFX1 \A_reg_reg[6]  ( .D(N15), .CLK(clk), .Q(A_reg[6]), .QN(n386) );
  DFFX1 \A_reg_reg[5]  ( .D(N14), .CLK(clk), .Q(A_reg[5]), .QN(n388) );
  DFFX1 \A_reg_reg[4]  ( .D(N13), .CLK(clk), .Q(A_reg[4]), .QN(n390) );
  DFFX1 \A_reg_reg[3]  ( .D(N12), .CLK(clk), .Q(A_reg[3]), .QN(n392) );
  DFFX1 \A_reg_reg[2]  ( .D(N11), .CLK(clk), .Q(A_reg[2]), .QN(n394) );
  DFFX1 \A_reg_reg[1]  ( .D(N10), .CLK(clk), .Q(A_reg[1]), .QN(n396) );
  DFFX1 \A_reg_reg[0]  ( .D(N9), .CLK(clk), .Q(A_reg[0]), .QN(n398) );
  DFFX1 \B_reg_reg[30]  ( .D(N71), .CLK(clk), .Q(B_reg[30]) );
  DFFX1 \B_reg_reg[29]  ( .D(N70), .CLK(clk), .Q(B_reg[29]) );
  DFFX1 \B_reg_reg[28]  ( .D(N69), .CLK(clk), .Q(B_reg[28]) );
  DFFX1 \B_reg_reg[27]  ( .D(N68), .CLK(clk), .Q(B_reg[27]) );
  DFFX1 \B_reg_reg[26]  ( .D(N67), .CLK(clk), .Q(B_reg[26]) );
  DFFX1 \B_reg_reg[25]  ( .D(N66), .CLK(clk), .Q(B_reg[25]) );
  DFFX1 \B_reg_reg[24]  ( .D(N65), .CLK(clk), .Q(B_reg[24]) );
  DFFX1 \B_reg_reg[23]  ( .D(N64), .CLK(clk), .Q(B_reg[23]) );
  DFFX1 \B_reg_reg[22]  ( .D(N63), .CLK(clk), .Q(B_reg[22]) );
  DFFX1 \B_reg_reg[21]  ( .D(N62), .CLK(clk), .Q(B_reg[21]) );
  DFFX1 \B_reg_reg[20]  ( .D(N61), .CLK(clk), .Q(B_reg[20]) );
  DFFX1 \B_reg_reg[19]  ( .D(N60), .CLK(clk), .Q(B_reg[19]) );
  DFFX1 \B_reg_reg[18]  ( .D(N59), .CLK(clk), .Q(B_reg[18]) );
  DFFX1 \B_reg_reg[17]  ( .D(N58), .CLK(clk), .Q(B_reg[17]) );
  DFFX1 \B_reg_reg[16]  ( .D(N57), .CLK(clk), .Q(B_reg[16]) );
  DFFX1 \B_reg_reg[15]  ( .D(N56), .CLK(clk), .Q(B_reg[15]) );
  DFFX1 \B_reg_reg[14]  ( .D(N55), .CLK(clk), .Q(B_reg[14]) );
  DFFX1 \B_reg_reg[13]  ( .D(N54), .CLK(clk), .Q(B_reg[13]) );
  DFFX1 \B_reg_reg[12]  ( .D(N53), .CLK(clk), .Q(B_reg[12]) );
  DFFX1 \B_reg_reg[11]  ( .D(N52), .CLK(clk), .Q(B_reg[11]) );
  DFFX1 \B_reg_reg[10]  ( .D(N51), .CLK(clk), .Q(B_reg[10]) );
  DFFX1 \B_reg_reg[9]  ( .D(N50), .CLK(clk), .Q(B_reg[9]) );
  DFFX1 \B_reg_reg[8]  ( .D(N49), .CLK(clk), .Q(B_reg[8]) );
  DFFX1 \B_reg_reg[7]  ( .D(N48), .CLK(clk), .Q(B_reg[7]) );
  DFFX1 \B_reg_reg[6]  ( .D(N47), .CLK(clk), .Q(B_reg[6]) );
  DFFX1 \B_reg_reg[5]  ( .D(N46), .CLK(clk), .Q(B_reg[5]) );
  DFFX1 \B_reg_reg[4]  ( .D(N45), .CLK(clk), .Q(B_reg[4]) );
  DFFX1 \B_reg_reg[3]  ( .D(N44), .CLK(clk), .Q(B_reg[3]) );
  DFFX1 \B_reg_reg[2]  ( .D(N43), .CLK(clk), .Q(B_reg[2]) );
  DFFX1 \B_reg_reg[1]  ( .D(N42), .CLK(clk), .Q(B_reg[1]) );
  DFFX1 \B_reg_reg[0]  ( .D(N41), .CLK(clk), .Q(B_reg[0]) );
  DFFARX1 \counter_reg[0]  ( .D(N497), .CLK(internalClk), .RSTB(n973), .Q(
        counter[0]), .QN(n406) );
  DFFARX1 \counter_reg[1]  ( .D(N498), .CLK(internalClk), .RSTB(n976), .Q(
        counter[1]), .QN(n405) );
  DFFARX1 \counter_reg[2]  ( .D(N499), .CLK(internalClk), .RSTB(n975), .Q(
        counter[2]), .QN(n404) );
  DFFARX1 \counter_reg[3]  ( .D(N500), .CLK(internalClk), .RSTB(n976), .Q(
        counter[3]), .QN(n402) );
  DFFARX1 \counter_reg[4]  ( .D(N501), .CLK(internalClk), .RSTB(n972), .Q(
        counter[4]), .QN(n403) );
  DFFARX1 \counter_reg[5]  ( .D(N502), .CLK(internalClk), .RSTB(n975), .Q(
        counter[5]), .QN(n241) );
  DFFARX1 \counter_reg[6]  ( .D(N503), .CLK(internalClk), .RSTB(n975), .Q(n866), .QN(n885) );
  DFFARX1 \counter_reg[7]  ( .D(N504), .CLK(internalClk), .RSTB(n974), .Q(
        counter[7]), .QN(n886) );
  DFFARX1 \counter_reg[8]  ( .D(N505), .CLK(internalClk), .RSTB(n972), .Q(
        counter[8]), .QN(n233) );
  DFFARX1 \counter_reg[9]  ( .D(N506), .CLK(internalClk), .RSTB(n972), .Q(
        counter[9]), .QN(n234) );
  DFFARX1 \counter_reg[10]  ( .D(N507), .CLK(internalClk), .RSTB(n971), .Q(
        counter[10]), .QN(n236) );
  DFFARX1 \counter_reg[11]  ( .D(N508), .CLK(internalClk), .RSTB(n974), .Q(
        counter[11]), .QN(n897) );
  DFFARX1 \counter_reg[12]  ( .D(N509), .CLK(internalClk), .RSTB(n972), .Q(
        counter[12]), .QN(n235) );
  DFFARX1 \counter_reg[13]  ( .D(N510), .CLK(internalClk), .RSTB(n974), .Q(
        counter[13]), .QN(n888) );
  DFFARX1 \counter_reg[14]  ( .D(N511), .CLK(internalClk), .RSTB(n973), .Q(
        counter[14]), .QN(n893) );
  DFFARX1 \counter_reg[15]  ( .D(N512), .CLK(internalClk), .RSTB(n972), .Q(
        counter[15]), .QN(n894) );
  DFFARX1 \counter_reg[16]  ( .D(N513), .CLK(internalClk), .RSTB(n971), .Q(
        n869), .QN(n898) );
  DFFARX1 \counter_reg[17]  ( .D(N514), .CLK(internalClk), .RSTB(n971), .Q(
        counter[17]), .QN(n237) );
  DFFARX1 \counter_reg[18]  ( .D(N515), .CLK(internalClk), .RSTB(n973), .Q(
        counter[18]), .QN(n238) );
  DFFARX1 \counter_reg[19]  ( .D(N516), .CLK(internalClk), .RSTB(n971), .Q(
        counter[19]), .QN(n230) );
  DFFARX1 \counter_reg[20]  ( .D(N517), .CLK(internalClk), .RSTB(n975), .Q(
        n865), .QN(n892) );
  DFFARX1 \counter_reg[21]  ( .D(N518), .CLK(internalClk), .RSTB(n974), .Q(
        counter[21]), .QN(n228) );
  DFFARX1 \counter_reg[22]  ( .D(N519), .CLK(internalClk), .RSTB(n972), .Q(
        counter[22]), .QN(n229) );
  DFFARX1 \counter_reg[23]  ( .D(N520), .CLK(internalClk), .RSTB(n974), .Q(
        counter[23]), .QN(n239) );
  DFFARX1 \counter_reg[24]  ( .D(N521), .CLK(internalClk), .RSTB(n975), .Q(
        counter[24]), .QN(n914) );
  DFFARX1 \counter_reg[25]  ( .D(N522), .CLK(internalClk), .RSTB(n971), .Q(
        counter[25]), .QN(n889) );
  DFFARX1 \counter_reg[26]  ( .D(N523), .CLK(internalClk), .RSTB(n973), .Q(
        counter[26]), .QN(n231) );
  DFFARX1 \counter_reg[27]  ( .D(N524), .CLK(internalClk), .RSTB(n975), .Q(
        counter[27]), .QN(n232) );
  DFFARX1 \counter_reg[28]  ( .D(N525), .CLK(internalClk), .RSTB(n974), .Q(
        counter[28]), .QN(n895) );
  DFFARX1 \counter_reg[29]  ( .D(N526), .CLK(internalClk), .RSTB(n971), .Q(
        counter[29]), .QN(n890) );
  DFFARX1 \counter_reg[30]  ( .D(N527), .CLK(internalClk), .RSTB(n973), .Q(
        counter[30]), .QN(n242) );
  DFFARX1 \counter_reg[31]  ( .D(N528), .CLK(internalClk), .RSTB(n973), .Q(
        counter[31]), .QN(n240) );
  DFFX1 \P_reg[63]  ( .D(N596), .CLK(clk), .Q(P[63]) );
  DFFX1 \P_reg[62]  ( .D(N595), .CLK(clk), .Q(P[62]) );
  DFFX1 \P_reg[61]  ( .D(N594), .CLK(clk), .Q(P[61]) );
  DFFX1 \P_reg[60]  ( .D(N593), .CLK(clk), .Q(P[60]) );
  DFFX1 \P_reg[59]  ( .D(N592), .CLK(clk), .Q(P[59]) );
  DFFX1 \P_reg[58]  ( .D(N591), .CLK(clk), .Q(P[58]) );
  DFFX1 \P_reg[57]  ( .D(N590), .CLK(clk), .Q(P[57]) );
  DFFX1 \P_reg[56]  ( .D(N589), .CLK(clk), .Q(P[56]) );
  DFFX1 \P_reg[55]  ( .D(N588), .CLK(clk), .Q(P[55]) );
  DFFX1 \P_reg[54]  ( .D(N587), .CLK(clk), .Q(P[54]) );
  DFFX1 \P_reg[53]  ( .D(N586), .CLK(clk), .Q(P[53]) );
  DFFX1 \P_reg[52]  ( .D(N585), .CLK(clk), .Q(P[52]) );
  DFFX1 \P_reg[51]  ( .D(N584), .CLK(clk), .Q(P[51]) );
  DFFX1 \P_reg[50]  ( .D(N583), .CLK(clk), .Q(P[50]) );
  DFFX1 \P_reg[49]  ( .D(N582), .CLK(clk), .Q(P[49]) );
  DFFX1 \P_reg[48]  ( .D(N581), .CLK(clk), .Q(P[48]) );
  DFFX1 \P_reg[47]  ( .D(N580), .CLK(clk), .Q(P[47]) );
  DFFX1 \P_reg[46]  ( .D(N579), .CLK(clk), .Q(P[46]) );
  DFFX1 \P_reg[45]  ( .D(N578), .CLK(clk), .Q(P[45]) );
  DFFX1 \P_reg[44]  ( .D(N577), .CLK(clk), .Q(P[44]) );
  DFFX1 \P_reg[43]  ( .D(N576), .CLK(clk), .Q(P[43]) );
  DFFX1 \P_reg[42]  ( .D(N575), .CLK(clk), .Q(P[42]) );
  DFFX1 \P_reg[41]  ( .D(N574), .CLK(clk), .Q(P[41]) );
  DFFX1 \P_reg[40]  ( .D(N573), .CLK(clk), .Q(P[40]) );
  DFFX1 \P_reg[39]  ( .D(N572), .CLK(clk), .Q(P[39]) );
  DFFX1 \P_reg[38]  ( .D(N571), .CLK(clk), .Q(P[38]) );
  DFFX1 \P_reg[37]  ( .D(N570), .CLK(clk), .Q(P[37]) );
  DFFX1 \P_reg[36]  ( .D(N569), .CLK(clk), .Q(P[36]) );
  DFFX1 \P_reg[35]  ( .D(N568), .CLK(clk), .Q(P[35]) );
  DFFX1 \P_reg[34]  ( .D(N567), .CLK(clk), .Q(P[34]) );
  DFFX1 \P_reg[33]  ( .D(N566), .CLK(clk), .Q(P[33]) );
  DFFX1 \P_reg[32]  ( .D(N565), .CLK(clk), .Q(P[32]) );
  DFFX1 \P_reg[31]  ( .D(N564), .CLK(clk), .Q(P[31]) );
  DFFX1 \P_reg[30]  ( .D(N563), .CLK(clk), .Q(P[30]) );
  DFFX1 \P_reg[29]  ( .D(N562), .CLK(clk), .Q(P[29]) );
  DFFX1 \P_reg[28]  ( .D(N561), .CLK(clk), .Q(P[28]) );
  DFFX1 \P_reg[27]  ( .D(N560), .CLK(clk), .Q(P[27]) );
  DFFX1 \P_reg[26]  ( .D(N559), .CLK(clk), .Q(P[26]) );
  DFFX1 \P_reg[25]  ( .D(N558), .CLK(clk), .Q(P[25]) );
  DFFX1 \P_reg[24]  ( .D(N557), .CLK(clk), .Q(P[24]) );
  DFFX1 \P_reg[23]  ( .D(N556), .CLK(clk), .Q(P[23]) );
  DFFX1 \P_reg[22]  ( .D(N555), .CLK(clk), .Q(P[22]) );
  DFFX1 \P_reg[21]  ( .D(N554), .CLK(clk), .Q(P[21]) );
  DFFX1 \P_reg[20]  ( .D(N553), .CLK(clk), .Q(P[20]) );
  DFFX1 \P_reg[19]  ( .D(N552), .CLK(clk), .Q(P[19]) );
  DFFX1 \P_reg[18]  ( .D(N551), .CLK(clk), .Q(P[18]) );
  DFFX1 \P_reg[17]  ( .D(N550), .CLK(clk), .Q(P[17]) );
  DFFX1 \P_reg[16]  ( .D(N549), .CLK(clk), .Q(P[16]) );
  DFFX1 \P_reg[15]  ( .D(N548), .CLK(clk), .Q(P[15]) );
  DFFX1 \P_reg[14]  ( .D(N547), .CLK(clk), .Q(P[14]) );
  DFFX1 \P_reg[13]  ( .D(N546), .CLK(clk), .Q(P[13]) );
  DFFX1 \P_reg[12]  ( .D(N545), .CLK(clk), .Q(P[12]) );
  DFFX1 \P_reg[11]  ( .D(N544), .CLK(clk), .Q(P[11]) );
  DFFX1 \P_reg[10]  ( .D(N543), .CLK(clk), .Q(P[10]) );
  DFFX1 \P_reg[9]  ( .D(N542), .CLK(clk), .Q(P[9]) );
  DFFX1 \P_reg[8]  ( .D(N541), .CLK(clk), .Q(P[8]) );
  DFFX1 \P_reg[7]  ( .D(N540), .CLK(clk), .Q(P[7]) );
  DFFX1 \P_reg[6]  ( .D(N539), .CLK(clk), .Q(P[6]) );
  DFFX1 \P_reg[5]  ( .D(N538), .CLK(clk), .Q(P[5]) );
  DFFX1 \P_reg[4]  ( .D(N537), .CLK(clk), .Q(P[4]) );
  DFFX1 \P_reg[3]  ( .D(N536), .CLK(clk), .Q(P[3]) );
  DFFX1 \P_reg[2]  ( .D(N535), .CLK(clk), .Q(P[2]) );
  DFFX1 \P_reg[1]  ( .D(N534), .CLK(clk), .Q(P[1]) );
  DFFX1 \P_reg[0]  ( .D(N533), .CLK(clk), .Q(P[0]) );
  DFFX1 \multiplier_reg[31]  ( .D(n598), .CLK(internalClk), .Q(n661) );
  DFFX1 \Accumulator_reg[30]  ( .D(n597), .CLK(internalClk), .Q(n685), .QN(
        n438) );
  DFFX1 \Accumulator_reg[29]  ( .D(n596), .CLK(internalClk), .Q(n711), .QN(
        n437) );
  DFFX1 \Accumulator_reg[28]  ( .D(n595), .CLK(internalClk), .Q(n707), .QN(
        n436) );
  DFFX1 \Accumulator_reg[27]  ( .D(n594), .CLK(internalClk), .Q(n686), .QN(
        n435) );
  DFFX1 \Accumulator_reg[26]  ( .D(n593), .CLK(internalClk), .Q(n687), .QN(
        n434) );
  DFFX1 \Accumulator_reg[25]  ( .D(n592), .CLK(internalClk), .Q(n688), .QN(
        n433) );
  DFFX1 \Accumulator_reg[24]  ( .D(n591), .CLK(internalClk), .Q(n706), .QN(
        n432) );
  DFFX1 \Accumulator_reg[23]  ( .D(n590), .CLK(internalClk), .Q(n689), .QN(
        n431) );
  DFFX1 \Accumulator_reg[22]  ( .D(n589), .CLK(internalClk), .Q(n690), .QN(
        n430) );
  DFFX1 \Accumulator_reg[21]  ( .D(n588), .CLK(internalClk), .Q(n705), .QN(
        n429) );
  DFFX1 \Accumulator_reg[20]  ( .D(n587), .CLK(internalClk), .Q(n691), .QN(
        n428) );
  DFFX1 \Accumulator_reg[19]  ( .D(n586), .CLK(internalClk), .Q(n704), .QN(
        n427) );
  DFFX1 \Accumulator_reg[18]  ( .D(n585), .CLK(internalClk), .Q(n684), .QN(
        n426) );
  DFFX1 \Accumulator_reg[17]  ( .D(n584), .CLK(internalClk), .Q(n710), .QN(
        n425) );
  DFFX1 \Accumulator_reg[16]  ( .D(n583), .CLK(internalClk), .Q(n692), .QN(
        n424) );
  DFFX1 \Accumulator_reg[15]  ( .D(n582), .CLK(internalClk), .Q(n693), .QN(
        n423) );
  DFFX1 \Accumulator_reg[14]  ( .D(n581), .CLK(internalClk), .Q(n712), .QN(
        n422) );
  DFFX1 \Accumulator_reg[13]  ( .D(n580), .CLK(internalClk), .Q(n682), .QN(
        n421) );
  DFFX1 \Accumulator_reg[12]  ( .D(n579), .CLK(internalClk), .Q(n694), .QN(
        n420) );
  DFFX1 \Accumulator_reg[11]  ( .D(n578), .CLK(internalClk), .Q(n708), .QN(
        n419) );
  DFFX1 \Accumulator_reg[10]  ( .D(n577), .CLK(internalClk), .Q(n695), .QN(
        n418) );
  DFFX1 \Accumulator_reg[9]  ( .D(n576), .CLK(internalClk), .Q(n696), .QN(n417) );
  DFFX1 \Accumulator_reg[8]  ( .D(n575), .CLK(internalClk), .Q(n709), .QN(n416) );
  DFFX1 \Accumulator_reg[7]  ( .D(n574), .CLK(internalClk), .Q(n697), .QN(n415) );
  DFFX1 \Accumulator_reg[6]  ( .D(n573), .CLK(internalClk), .Q(n698), .QN(n414) );
  DFFX1 \Accumulator_reg[5]  ( .D(n572), .CLK(internalClk), .Q(n699), .QN(n413) );
  DFFX1 \Accumulator_reg[4]  ( .D(n571), .CLK(internalClk), .Q(n700), .QN(n412) );
  DFFX1 \Accumulator_reg[3]  ( .D(n570), .CLK(internalClk), .Q(n701), .QN(n411) );
  DFFX1 \Accumulator_reg[2]  ( .D(n569), .CLK(internalClk), .Q(n702), .QN(n410) );
  DFFX1 \Accumulator_reg[1]  ( .D(n568), .CLK(internalClk), .Q(n703), .QN(n409) );
  DFFX1 \Accumulator_reg[0]  ( .D(n567), .CLK(internalClk), .Q(n683), .QN(n408) );
  DFFX1 \multiplier_reg[30]  ( .D(n566), .CLK(internalClk), .Q(n659) );
  DFFX1 \multiplicand_reg[0]  ( .D(n565), .CLK(internalClk), .Q(n605) );
  DFFX1 \multiplicand_reg[1]  ( .D(n564), .CLK(internalClk), .Q(n612) );
  DFFX1 \multiplicand_reg[2]  ( .D(n563), .CLK(internalClk), .Q(n606) );
  DFFX1 \multiplicand_reg[3]  ( .D(n562), .CLK(internalClk), .Q(n607) );
  DFFX1 \multiplicand_reg[4]  ( .D(n561), .CLK(internalClk), .Q(n613) );
  DFFX1 \multiplicand_reg[5]  ( .D(n560), .CLK(internalClk), .Q(n614) );
  DFFX1 \multiplicand_reg[6]  ( .D(n559), .CLK(internalClk), .Q(n615) );
  DFFX1 \multiplicand_reg[7]  ( .D(n558), .CLK(internalClk), .Q(n608) );
  DFFX1 \multiplicand_reg[8]  ( .D(n557), .CLK(internalClk), .Q(n609) );
  DFFX1 \multiplicand_reg[9]  ( .D(n556), .CLK(internalClk), .Q(n610) );
  DFFX1 \multiplicand_reg[10]  ( .D(n555), .CLK(internalClk), .Q(n611) );
  DFFX1 \multiplicand_reg[11]  ( .D(n554), .CLK(internalClk), .Q(n603) );
  DFFX1 \multiplicand_reg[12]  ( .D(n553), .CLK(internalClk), .Q(n631) );
  DFFX1 \multiplicand_reg[13]  ( .D(n552), .CLK(internalClk), .Q(n616) );
  DFFX1 \multiplicand_reg[14]  ( .D(n551), .CLK(internalClk), .Q(n617) );
  DFFX1 \multiplicand_reg[15]  ( .D(n550), .CLK(internalClk), .Q(n618) );
  DFFX1 \multiplicand_reg[16]  ( .D(n549), .CLK(internalClk), .Q(n632) );
  DFFX1 \multiplicand_reg[17]  ( .D(n548), .CLK(internalClk), .Q(n619) );
  DFFX1 \multiplicand_reg[18]  ( .D(n547), .CLK(internalClk), .Q(n633) );
  DFFX1 \multiplicand_reg[19]  ( .D(n546), .CLK(internalClk), .Q(n634) );
  DFFX1 \multiplicand_reg[20]  ( .D(n545), .CLK(internalClk), .Q(n662) );
  DFFX1 \multiplicand_reg[21]  ( .D(n544), .CLK(internalClk), .Q(n663) );
  DFFX1 \multiplicand_reg[22]  ( .D(n543), .CLK(internalClk), .Q(n664) );
  DFFX1 \multiplicand_reg[23]  ( .D(n542), .CLK(internalClk), .Q(n665) );
  DFFX1 \multiplicand_reg[24]  ( .D(n541), .CLK(internalClk), .Q(n670) );
  DFFX1 \multiplicand_reg[25]  ( .D(n540), .CLK(internalClk), .Q(n666) );
  DFFX1 \multiplicand_reg[26]  ( .D(n539), .CLK(internalClk), .Q(n667) );
  DFFX1 \multiplicand_reg[27]  ( .D(n538), .CLK(internalClk), .Q(n671) );
  DFFX1 \multiplicand_reg[28]  ( .D(n537), .CLK(internalClk), .Q(n668) );
  DFFX1 \multiplicand_reg[29]  ( .D(n536), .CLK(internalClk), .Q(n669) );
  DFFX1 \multiplicand_reg[30]  ( .D(n535), .CLK(internalClk), .Q(n673) );
  DFFX1 \multiplicand_reg[31]  ( .D(n534), .CLK(internalClk), .Q(n674) );
  DFFX1 \multiplier_reg[29]  ( .D(n533), .CLK(internalClk), .Q(n672) );
  DFFX1 \multiplier_reg[28]  ( .D(n532), .CLK(internalClk), .Q(n643) );
  DFFX1 \multiplier_reg[27]  ( .D(n531), .CLK(internalClk), .Q(n644) );
  DFFX1 \multiplier_reg[26]  ( .D(n530), .CLK(internalClk), .Q(n645) );
  DFFX1 \multiplier_reg[25]  ( .D(n529), .CLK(internalClk), .Q(n646) );
  DFFX1 \multiplier_reg[24]  ( .D(n528), .CLK(internalClk), .Q(n623) );
  DFFX1 \multiplier_reg[23]  ( .D(n527), .CLK(internalClk), .Q(n647) );
  DFFX1 \multiplier_reg[22]  ( .D(n526), .CLK(internalClk), .Q(n648) );
  DFFX1 \multiplier_reg[21]  ( .D(n525), .CLK(internalClk), .Q(n649) );
  DFFX1 \multiplier_reg[20]  ( .D(n524), .CLK(internalClk), .Q(n624) );
  DFFX1 \multiplier_reg[19]  ( .D(n523), .CLK(internalClk), .Q(n650) );
  DFFX1 \multiplier_reg[18]  ( .D(n522), .CLK(internalClk), .Q(n651) );
  DFFX1 \multiplier_reg[17]  ( .D(n521), .CLK(internalClk), .Q(n790) );
  DFFX1 \multiplier_reg[16]  ( .D(n520), .CLK(internalClk), .Q(n625) );
  DFFX1 \multiplier_reg[15]  ( .D(n519), .CLK(internalClk), .Q(n652) );
  DFFX1 \multiplier_reg[14]  ( .D(n518), .CLK(internalClk), .Q(n653) );
  DFFX1 \multiplier_reg[13]  ( .D(n517), .CLK(internalClk), .Q(n654) );
  DFFX1 \multiplier_reg[12]  ( .D(n516), .CLK(internalClk), .Q(n626) );
  DFFX1 \multiplier_reg[11]  ( .D(n515), .CLK(internalClk), .Q(n655) );
  DFFX1 \multiplier_reg[10]  ( .D(n514), .CLK(internalClk), .Q(n656) );
  DFFX1 \multiplier_reg[9]  ( .D(n513), .CLK(internalClk), .Q(n660) );
  DFFX1 \multiplier_reg[8]  ( .D(n512), .CLK(internalClk), .Q(n627) );
  DFFX1 \multiplier_reg[7]  ( .D(n511), .CLK(internalClk), .Q(n657) );
  DFFX1 \multiplier_reg[6]  ( .D(n510), .CLK(internalClk), .Q(n789) );
  DFFX1 \multiplier_reg[5]  ( .D(n509), .CLK(internalClk), .Q(n628) );
  DFFX1 \multiplier_reg[4]  ( .D(n508), .CLK(internalClk), .Q(n604) );
  DFFX1 \multiplier_reg[3]  ( .D(n507), .CLK(internalClk), .Q(n658) );
  DFFX1 \multiplier_reg[2]  ( .D(n506), .CLK(internalClk), .Q(n629) );
  DFFX1 \multiplier_reg[1]  ( .D(n505), .CLK(internalClk), .Q(n630) );
  DFFX1 \multiplier_reg[0]  ( .D(n504), .CLK(internalClk), .Q(n792) );
  DFFX1 \P_reg_reg[0]  ( .D(n503), .CLK(internalClk), .Q(n713), .QN(n306) );
  DFFX1 \P_reg_reg[1]  ( .D(n502), .CLK(internalClk), .Q(n714), .QN(n305) );
  DFFX1 \P_reg_reg[2]  ( .D(n501), .CLK(internalClk), .Q(n715), .QN(n304) );
  DFFX1 \P_reg_reg[3]  ( .D(n500), .CLK(internalClk), .Q(n716), .QN(n303) );
  DFFX1 \P_reg_reg[4]  ( .D(n499), .CLK(internalClk), .Q(n717), .QN(n302) );
  DFFX1 \P_reg_reg[5]  ( .D(n498), .CLK(internalClk), .Q(n718), .QN(n301) );
  DFFX1 \P_reg_reg[6]  ( .D(n497), .CLK(internalClk), .Q(n719), .QN(n300) );
  DFFX1 \P_reg_reg[7]  ( .D(n496), .CLK(internalClk), .Q(n720), .QN(n299) );
  DFFX1 \P_reg_reg[8]  ( .D(n495), .CLK(internalClk), .Q(n721), .QN(n298) );
  DFFX1 \P_reg_reg[9]  ( .D(n494), .CLK(internalClk), .Q(n722), .QN(n297) );
  DFFX1 \P_reg_reg[10]  ( .D(n493), .CLK(internalClk), .Q(n723), .QN(n296) );
  DFFX1 \P_reg_reg[11]  ( .D(n492), .CLK(internalClk), .Q(n724), .QN(n295) );
  DFFX1 \P_reg_reg[12]  ( .D(n491), .CLK(internalClk), .Q(n725), .QN(n294) );
  DFFX1 \P_reg_reg[13]  ( .D(n490), .CLK(internalClk), .Q(n726), .QN(n293) );
  DFFX1 \P_reg_reg[14]  ( .D(n489), .CLK(internalClk), .Q(n727), .QN(n292) );
  DFFX1 \P_reg_reg[15]  ( .D(n488), .CLK(internalClk), .Q(n728), .QN(n291) );
  DFFX1 \P_reg_reg[16]  ( .D(n487), .CLK(internalClk), .Q(n729), .QN(n290) );
  DFFX1 \P_reg_reg[17]  ( .D(n486), .CLK(internalClk), .Q(n730), .QN(n289) );
  DFFX1 \P_reg_reg[18]  ( .D(n485), .CLK(internalClk), .Q(n731), .QN(n288) );
  DFFX1 \P_reg_reg[19]  ( .D(n484), .CLK(internalClk), .Q(n732), .QN(n287) );
  DFFX1 \P_reg_reg[20]  ( .D(n483), .CLK(internalClk), .Q(n733), .QN(n286) );
  DFFX1 \P_reg_reg[21]  ( .D(n482), .CLK(internalClk), .Q(n734), .QN(n285) );
  DFFX1 \P_reg_reg[22]  ( .D(n481), .CLK(internalClk), .Q(n735), .QN(n284) );
  DFFX1 \P_reg_reg[23]  ( .D(n480), .CLK(internalClk), .Q(n736), .QN(n283) );
  DFFX1 \P_reg_reg[24]  ( .D(n479), .CLK(internalClk), .Q(n737), .QN(n282) );
  DFFX1 \P_reg_reg[25]  ( .D(n478), .CLK(internalClk), .Q(n738), .QN(n281) );
  DFFX1 \P_reg_reg[26]  ( .D(n477), .CLK(internalClk), .Q(n739), .QN(n280) );
  DFFX1 \P_reg_reg[27]  ( .D(n476), .CLK(internalClk), .Q(n740), .QN(n279) );
  DFFX1 \P_reg_reg[28]  ( .D(n475), .CLK(internalClk), .Q(n741), .QN(n278) );
  DFFX1 \P_reg_reg[30]  ( .D(n474), .CLK(internalClk), .Q(n743), .QN(n277) );
  DFFX1 \P_reg_reg[31]  ( .D(n473), .CLK(internalClk), .Q(n744), .QN(n276) );
  DFFX1 \P_reg_reg[32]  ( .D(n472), .CLK(internalClk), .Q(n745), .QN(n275) );
  DFFX1 \P_reg_reg[33]  ( .D(n471), .CLK(internalClk), .Q(n746), .QN(n274) );
  DFFX1 \P_reg_reg[34]  ( .D(n470), .CLK(internalClk), .Q(n747), .QN(n273) );
  DFFX1 \P_reg_reg[35]  ( .D(n469), .CLK(internalClk), .Q(n748), .QN(n272) );
  DFFX1 \P_reg_reg[36]  ( .D(n468), .CLK(internalClk), .Q(n749), .QN(n271) );
  DFFX1 \P_reg_reg[37]  ( .D(n467), .CLK(internalClk), .Q(n750), .QN(n270) );
  DFFX1 \P_reg_reg[38]  ( .D(n466), .CLK(internalClk), .Q(n751), .QN(n269) );
  DFFX1 \P_reg_reg[39]  ( .D(n465), .CLK(internalClk), .Q(n752), .QN(n268) );
  DFFX1 \P_reg_reg[40]  ( .D(n464), .CLK(internalClk), .Q(n753), .QN(n267) );
  DFFX1 \P_reg_reg[41]  ( .D(n463), .CLK(internalClk), .Q(n754), .QN(n266) );
  DFFX1 \P_reg_reg[42]  ( .D(n462), .CLK(internalClk), .Q(n755), .QN(n265) );
  DFFX1 \P_reg_reg[43]  ( .D(n461), .CLK(internalClk), .Q(n756), .QN(n264) );
  DFFX1 \P_reg_reg[44]  ( .D(n460), .CLK(internalClk), .Q(n757), .QN(n263) );
  DFFX1 \P_reg_reg[45]  ( .D(n459), .CLK(internalClk), .Q(n758), .QN(n262) );
  DFFX1 \P_reg_reg[46]  ( .D(n458), .CLK(internalClk), .Q(n759), .QN(n261) );
  DFFX1 \P_reg_reg[47]  ( .D(n457), .CLK(internalClk), .Q(n675), .QN(n260) );
  DFFX1 \P_reg_reg[48]  ( .D(n456), .CLK(internalClk), .Q(n760), .QN(n259) );
  DFFX1 \P_reg_reg[49]  ( .D(n455), .CLK(internalClk), .Q(n761), .QN(n258) );
  DFFX1 \P_reg_reg[50]  ( .D(n454), .CLK(internalClk), .Q(n762), .QN(n257) );
  DFFX1 \P_reg_reg[51]  ( .D(n453), .CLK(internalClk), .Q(n763), .QN(n256) );
  DFFX1 \P_reg_reg[52]  ( .D(n452), .CLK(internalClk), .Q(n764), .QN(n255) );
  DFFX1 \P_reg_reg[53]  ( .D(n451), .CLK(internalClk), .Q(n765), .QN(n254) );
  DFFX1 \P_reg_reg[54]  ( .D(n450), .CLK(internalClk), .Q(n766), .QN(n253) );
  DFFX1 \P_reg_reg[55]  ( .D(n449), .CLK(internalClk), .Q(n680), .QN(n252) );
  DFFX1 \P_reg_reg[56]  ( .D(n448), .CLK(internalClk), .Q(n679), .QN(n251) );
  DFFX1 \P_reg_reg[57]  ( .D(n447), .CLK(internalClk), .Q(n677), .QN(n250) );
  DFFX1 \P_reg_reg[58]  ( .D(n446), .CLK(internalClk), .Q(n769), .QN(n249) );
  DFFX1 \P_reg_reg[59]  ( .D(n445), .CLK(internalClk), .Q(n678), .QN(n248) );
  DFFX1 \P_reg_reg[60]  ( .D(n444), .CLK(internalClk), .Q(n676), .QN(n247) );
  DFFX1 \P_reg_reg[61]  ( .D(n443), .CLK(internalClk), .Q(n681), .QN(n246) );
  DFFX1 \P_reg_reg[62]  ( .D(n442), .CLK(internalClk), .Q(n768), .QN(n245) );
  DFFX1 \P_reg_reg[63]  ( .D(n441), .CLK(internalClk), .Q(n767), .QN(n244) );
  DFFX1 \P_reg_reg[29]  ( .D(n440), .CLK(internalClk), .Q(n742), .QN(n243) );
  SeqMult_DW02_mult_0 mult_add_51_S2_aco ( .A({N205, N206, N207, N208, N209, 
        N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, 
        N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, 
        N234, N235, N236}), .B(N268), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, N697, N696, N695, N694, N693, N692, N691, 
        N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, 
        N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, 
        N666}) );
  SeqMult_DW01_sub_4 sub_46_S2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B(B_reg), .CI(1'b0), .DIFF({N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, 
        N143, N142, N141}) );
  SeqMult_DW01_inc_1 add_60 ( .A({counter[31:29], n896, counter[27:21], n865, 
        counter[19:17], n869, counter[15:7], n866, counter[5:0]}), .SUM({N496, 
        N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, 
        N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, 
        N471, N470, N469, N468, N467, N466, N465}) );
  SeqMult_DW01_sub_8 sub_59_S2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, N334, 
        N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, 
        N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, 
        N309, N308, N307, N306, N305, N304, N303, N237, N238, N239, N240, N241, 
        N242, N243, N244, N245, N246, N247, N248, N249, N250, n602, N252, N253, 
        N254, N255, N256, N257, N258, N259, N260, N261, n601, N263, N264, N265, 
        N266, N267}), .CI(1'b0), .DIFF({N400, N399, N398, N397, N396, N395, 
        N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, 
        N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, 
        N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, 
        N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, 
        N346, N345, N344, N343, N342, N341, N340, N339, N338, N337}) );
  SeqMult_DW01_add_3 add_51_S2_aco ( .A({1'b0, N829, N831, N833, N835, N837, 
        N839, N841, N843, N845, N847, N849, N851, N853, N855, N857, N859, N861, 
        N863, N865, N867, N869, N871, N873, N875, N877, N879, N881, N883, N885, 
        N887, N889}), .B({N697, N696, N695, N694, N693, N692, N691, N690, N689, 
        N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, 
        N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666}), 
        .CI(1'b0), .SUM({N334, N333, N332, N331, N330, N329, N328, N327, N326, 
        N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, 
        N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303}) );
  SeqMult_DW01_sub_9 sub_43_S2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B(A_reg), .CI(1'b0), .DIFF({N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76})
         );
  DFFX1 \B_reg_reg[31]  ( .D(N72), .CLK(clk), .Q(B_reg[31]), .QN(n401) );
  OR2X1 U641 ( .IN1(n1035), .IN2(n372), .Q(n837) );
  NOR2X0 U642 ( .IN1(n421), .IN2(n936), .QN(N863) );
  AND2X1 U643 ( .IN1(n943), .IN2(B_reg[31]), .Q(n903) );
  AND3X1 U644 ( .IN1(counter[2]), .IN2(counter[1]), .IN3(counter[0]), .Q(n999)
         );
  INVX0 U645 ( .INP(n1053), .ZN(n1052) );
  NBUFFX2 U646 ( .INP(n904), .Z(n959) );
  NBUFFX2 U647 ( .INP(N329), .Z(n845) );
  DELLN1X2 U648 ( .INP(n998), .Z(n600) );
  NOR2X0 U649 ( .IN1(n408), .IN2(n932), .QN(N889) );
  NBUFFX2 U650 ( .INP(N315), .Z(n871) );
  NBUFFX2 U651 ( .INP(N322), .Z(n870) );
  NBUFFX2 U652 ( .INP(N323), .Z(n803) );
  NBUFFX2 U653 ( .INP(N333), .Z(n770) );
  NAND2X1 U654 ( .IN1(n954), .IN2(n676), .QN(n819) );
  NAND2X1 U655 ( .IN1(n954), .IN2(n678), .QN(n849) );
  NAND2X1 U656 ( .IN1(n952), .IN2(n677), .QN(n825) );
  NAND2X1 U657 ( .IN1(n953), .IN2(n679), .QN(n852) );
  MUX21X1 U658 ( .IN1(N258), .IN2(n660), .S(n967), .Q(n513) );
  MUX21X1 U659 ( .IN1(N238), .IN2(n672), .S(n966), .Q(n533) );
  MUX21X1 U660 ( .IN1(N237), .IN2(n659), .S(n965), .Q(n566) );
  MUX21X1 U661 ( .IN1(n807), .IN2(n709), .S(n965), .Q(n575) );
  MUX21X1 U662 ( .IN1(n871), .IN2(n708), .S(n964), .Q(n578) );
  MUX21X1 U663 ( .IN1(n881), .IN2(n712), .S(n964), .Q(n581) );
  MUX21X1 U664 ( .IN1(N321), .IN2(n710), .S(n965), .Q(n584) );
  MUX21X1 U665 ( .IN1(n803), .IN2(n704), .S(n964), .Q(n586) );
  MUX21X1 U666 ( .IN1(n794), .IN2(n705), .S(n967), .Q(n588) );
  MUX21X1 U667 ( .IN1(n800), .IN2(n706), .S(n964), .Q(n591) );
  MUX21X1 U668 ( .IN1(n864), .IN2(n707), .S(n964), .Q(n595) );
  MUX21X1 U669 ( .IN1(n770), .IN2(n711), .S(n964), .Q(n596) );
  INVX0 U670 ( .INP(n955), .ZN(n954) );
  AO222X1 U671 ( .IN1(N147), .IN2(n903), .IN3(B_reg[6]), .IN4(n907), .IN5(n780), .IN6(n789), .Q(n601) );
  AO222X1 U672 ( .IN1(N158), .IN2(n903), .IN3(B_reg[17]), .IN4(n907), .IN5(
        n779), .IN6(n790), .Q(n602) );
  AND2X1 U673 ( .IN1(n954), .IN2(n675), .Q(n620) );
  AND2X1 U674 ( .IN1(n822), .IN2(n821), .Q(n621) );
  AND2X1 U675 ( .IN1(n889), .IN2(n914), .Q(n622) );
  AND4X1 U676 ( .IN1(n236), .IN2(n241), .IN3(n233), .IN4(n234), .Q(n635) );
  OR2X1 U677 ( .IN1(n1035), .IN2(n396), .Q(n636) );
  AND2X1 U678 ( .IN1(n844), .IN2(n843), .Q(n637) );
  AND2X1 U679 ( .IN1(n621), .IN2(n1018), .Q(n638) );
  AND2X1 U680 ( .IN1(n815), .IN2(n816), .Q(n639) );
  AND2X1 U681 ( .IN1(n854), .IN2(n855), .Q(n640) );
  AND2X1 U682 ( .IN1(n857), .IN2(n858), .Q(n641) );
  NOR2X0 U683 ( .IN1(n891), .IN2(counter[28]), .QN(n642) );
  AND4X1 U684 ( .IN1(n1016), .IN2(n1022), .IN3(counter[3]), .IN4(n999), .Q(
        n909) );
  INVX0 U685 ( .INP(n796), .ZN(n797) );
  NAND2X0 U686 ( .IN1(n232), .IN2(n231), .QN(n1003) );
  NOR4X0 U687 ( .IN1(n1031), .IN2(n1033), .IN3(n1032), .IN4(counter[31]), .QN(
        n771) );
  INVX0 U688 ( .INP(n1035), .ZN(n772) );
  NAND4X0 U689 ( .IN1(n1008), .IN2(n1007), .IN3(n1006), .IN4(n1005), .QN(n773)
         );
  INVX0 U690 ( .INP(n882), .ZN(n774) );
  INVX0 U691 ( .INP(n882), .ZN(n775) );
  INVX0 U692 ( .INP(n774), .ZN(n776) );
  INVX0 U693 ( .INP(n774), .ZN(n777) );
  INVX0 U694 ( .INP(n774), .ZN(n778) );
  INVX0 U695 ( .INP(n775), .ZN(n779) );
  INVX0 U696 ( .INP(n775), .ZN(n780) );
  INVX0 U697 ( .INP(n775), .ZN(n781) );
  INVX0 U698 ( .INP(n775), .ZN(n782) );
  INVX0 U699 ( .INP(n775), .ZN(n783) );
  INVX0 U700 ( .INP(n775), .ZN(n784) );
  INVX0 U701 ( .INP(n775), .ZN(n785) );
  INVX0 U702 ( .INP(n775), .ZN(n786) );
  INVX0 U703 ( .INP(n775), .ZN(n787) );
  INVX0 U704 ( .INP(n775), .ZN(n788) );
  OR2X1 U705 ( .IN1(n1013), .IN2(n1012), .Q(n882) );
  AO221X1 U706 ( .IN1(N319), .IN2(n905), .IN3(N384), .IN4(n904), .IN5(n620), 
        .Q(n457) );
  AND2X2 U707 ( .IN1(n401), .IN2(n942), .Q(n916) );
  AND3X1 U708 ( .IN1(n399), .IN2(n771), .IN3(n901), .Q(n911) );
  AND2X2 U709 ( .IN1(n943), .IN2(B_reg[31]), .Q(n918) );
  NAND4X0 U710 ( .IN1(n1007), .IN2(n1006), .IN3(n862), .IN4(n1005), .QN(n1013)
         );
  AO222X1 U711 ( .IN1(n868), .IN2(n611), .IN3(n912), .IN4(n1046), .IN5(N86), 
        .IN6(n902), .Q(N226) );
  AND3X1 U712 ( .IN1(n908), .IN2(n901), .IN3(A_reg[31]), .Q(n902) );
  OR2X2 U713 ( .IN1(n887), .IN2(n846), .Q(n868) );
  AND4X1 U714 ( .IN1(n239), .IN2(n229), .IN3(n231), .IN4(n228), .Q(n791) );
  INVX0 U715 ( .INP(n791), .ZN(n1032) );
  AND4X1 U716 ( .IN1(n821), .IN2(n822), .IN3(n890), .IN4(n895), .Q(n793) );
  AO22X1 U717 ( .IN1(n1050), .IN2(n792), .IN3(n1017), .IN4(n638), .Q(N268) );
  DELLN1X2 U718 ( .INP(N325), .Z(n794) );
  OR2X4 U719 ( .IN1(n1013), .IN2(n846), .Q(n884) );
  DELLN1X2 U720 ( .INP(N317), .Z(n829) );
  AND3X1 U721 ( .IN1(n908), .IN2(n901), .IN3(A_reg[31]), .Q(n826) );
  NAND4X0 U722 ( .IN1(n228), .IN2(n230), .IN3(n239), .IN4(n229), .QN(n795) );
  INVX0 U723 ( .INP(n899), .ZN(n796) );
  AND3X1 U724 ( .IN1(n399), .IN2(n771), .IN3(n901), .Q(n899) );
  INVX0 U725 ( .INP(N316), .ZN(n798) );
  INVX0 U726 ( .INP(n798), .ZN(n799) );
  DELLN1X2 U727 ( .INP(N328), .Z(n800) );
  INVX0 U728 ( .INP(N310), .ZN(n801) );
  INVX0 U729 ( .INP(n801), .ZN(n802) );
  INVX0 U730 ( .INP(N314), .ZN(n804) );
  INVX0 U731 ( .INP(n804), .ZN(n805) );
  INVX0 U732 ( .INP(N312), .ZN(n806) );
  INVX0 U733 ( .INP(n806), .ZN(n807) );
  NAND2X0 U734 ( .IN1(n814), .IN2(n639), .QN(n446) );
  NAND2X0 U735 ( .IN1(N100), .IN2(n883), .QN(n808) );
  NAND2X0 U736 ( .IN1(n797), .IN2(A_reg[24]), .QN(n809) );
  NAND2X0 U737 ( .IN1(n784), .IN2(n670), .QN(n810) );
  NAND3X0 U738 ( .IN1(n808), .IN2(n809), .IN3(n810), .QN(N212) );
  INVX0 U739 ( .INP(N330), .ZN(n811) );
  INVX0 U740 ( .INP(n811), .ZN(n812) );
  NAND2X0 U741 ( .IN1(n237), .IN2(n236), .QN(n1000) );
  AND2X1 U742 ( .IN1(n832), .IN2(n831), .Q(n813) );
  NAND2X0 U743 ( .IN1(n960), .IN2(N395), .QN(n814) );
  NAND2X0 U744 ( .IN1(n812), .IN2(n951), .QN(n815) );
  NAND2X0 U745 ( .IN1(n952), .IN2(n769), .QN(n816) );
  NAND2X0 U746 ( .IN1(n960), .IN2(N397), .QN(n817) );
  NAND2X0 U747 ( .IN1(n864), .IN2(n951), .QN(n818) );
  NAND3X0 U748 ( .IN1(n817), .IN2(n818), .IN3(n819), .QN(n444) );
  NBUFFX2 U749 ( .INP(n904), .Z(n960) );
  NAND3X0 U750 ( .IN1(n771), .IN2(n399), .IN3(n901), .QN(n1035) );
  DELLN2X2 U751 ( .INP(n997), .Z(n820) );
  NAND2X0 U752 ( .IN1(n813), .IN2(n830), .QN(N222) );
  NAND2X0 U753 ( .IN1(n842), .IN2(n637), .QN(N221) );
  AND2X1 U754 ( .IN1(n406), .IN2(n405), .Q(n821) );
  AND2X1 U755 ( .IN1(n402), .IN2(n404), .Q(n822) );
  NAND2X0 U756 ( .IN1(n960), .IN2(N394), .QN(n823) );
  NAND2X0 U757 ( .IN1(n845), .IN2(n951), .QN(n824) );
  NAND3X0 U758 ( .IN1(n823), .IN2(n824), .IN3(n825), .QN(n447) );
  NAND2X0 U759 ( .IN1(N77), .IN2(n902), .QN(n827) );
  NAND2X0 U760 ( .IN1(n884), .IN2(n612), .QN(n828) );
  NAND3X0 U761 ( .IN1(n827), .IN2(n636), .IN3(n828), .QN(N235) );
  NBUFFX2 U762 ( .INP(n868), .Z(n929) );
  NAND2X0 U763 ( .IN1(n902), .IN2(N90), .QN(n830) );
  NAND2X0 U764 ( .IN1(n899), .IN2(n1048), .QN(n831) );
  NAND2X0 U765 ( .IN1(n884), .IN2(n617), .QN(n832) );
  NAND2X0 U766 ( .IN1(N93), .IN2(n902), .QN(n833) );
  NAND2X0 U767 ( .IN1(n912), .IN2(A_reg[17]), .QN(n834) );
  NAND2X0 U768 ( .IN1(n884), .IN2(n619), .QN(n835) );
  NAND3X0 U769 ( .IN1(n835), .IN2(n834), .IN3(n833), .QN(N219) );
  NAND2X0 U770 ( .IN1(N89), .IN2(n902), .QN(n836) );
  NAND2X0 U771 ( .IN1(n929), .IN2(n616), .QN(n838) );
  NAND3X0 U772 ( .IN1(n836), .IN2(n837), .IN3(n838), .QN(N223) );
  NBUFFX2 U773 ( .INP(n868), .Z(n931) );
  NBUFFX2 U774 ( .INP(n868), .Z(n930) );
  NAND2X0 U775 ( .IN1(N80), .IN2(n826), .QN(n839) );
  NAND2X0 U776 ( .IN1(n899), .IN2(n1040), .QN(n840) );
  NAND2X0 U777 ( .IN1(n884), .IN2(n613), .QN(n841) );
  NAND3X0 U778 ( .IN1(n839), .IN2(n840), .IN3(n841), .QN(N232) );
  NAND2X0 U779 ( .IN1(n826), .IN2(N91), .QN(n842) );
  NAND2X0 U780 ( .IN1(n899), .IN2(n1049), .QN(n843) );
  NAND2X0 U781 ( .IN1(n884), .IN2(n618), .QN(n844) );
  NAND4X0 U782 ( .IN1(n793), .IN2(n1009), .IN3(n1010), .IN4(n1011), .QN(n846)
         );
  NAND2X0 U783 ( .IN1(N396), .IN2(n960), .QN(n847) );
  NAND2X0 U784 ( .IN1(N331), .IN2(n951), .QN(n848) );
  NAND3X0 U785 ( .IN1(n847), .IN2(n848), .IN3(n849), .QN(n445) );
  NAND2X0 U786 ( .IN1(n853), .IN2(n640), .QN(n449) );
  NAND2X1 U787 ( .IN1(n953), .IN2(n680), .QN(n855) );
  NAND2X0 U788 ( .IN1(n960), .IN2(N393), .QN(n850) );
  NAND2X0 U789 ( .IN1(n800), .IN2(n951), .QN(n851) );
  NAND3X0 U790 ( .IN1(n850), .IN2(n851), .IN3(n852), .QN(n448) );
  DELLN1X2 U791 ( .INP(N318), .Z(n881) );
  NAND2X0 U792 ( .IN1(n856), .IN2(n641), .QN(n443) );
  NAND2X1 U793 ( .IN1(n954), .IN2(n681), .QN(n858) );
  NAND2X0 U794 ( .IN1(N392), .IN2(n960), .QN(n853) );
  NAND2X0 U795 ( .IN1(N327), .IN2(n951), .QN(n854) );
  NAND2X0 U796 ( .IN1(n960), .IN2(N398), .QN(n856) );
  NAND2X0 U797 ( .IN1(n770), .IN2(n951), .QN(n857) );
  NAND2X0 U798 ( .IN1(N95), .IN2(n826), .QN(n859) );
  NAND2X0 U799 ( .IN1(n772), .IN2(A_reg[19]), .QN(n860) );
  NAND2X0 U800 ( .IN1(n777), .IN2(n634), .QN(n861) );
  NAND3X0 U801 ( .IN1(n859), .IN2(n860), .IN3(n861), .QN(N217) );
  NAND2X0 U802 ( .IN1(n235), .IN2(n237), .QN(n1029) );
  NOR2X0 U803 ( .IN1(n1000), .IN2(n1001), .QN(n862) );
  INVX0 U804 ( .INP(N332), .ZN(n863) );
  INVX0 U805 ( .INP(n863), .ZN(n864) );
  NOR4X0 U806 ( .IN1(counter[3]), .IN2(counter[2]), .IN3(n1022), .IN4(n1021), 
        .QN(n1028) );
  NAND2X0 U807 ( .IN1(n892), .IN2(n898), .QN(n1023) );
  NAND2X0 U808 ( .IN1(n885), .IN2(n886), .QN(n1025) );
  NOR2X0 U809 ( .IN1(n998), .IN2(n867), .QN(n1017) );
  OR2X1 U810 ( .IN1(n997), .IN2(counter[4]), .Q(n867) );
  OR2X1 U811 ( .IN1(n773), .IN2(n1012), .Q(n1050) );
  NAND2X0 U812 ( .IN1(n888), .IN2(n897), .QN(n1026) );
  AO22X1 U813 ( .IN1(N107), .IN2(n944), .IN3(n787), .IN4(n674), .Q(N205) );
  NBUFFX2 U814 ( .INP(n902), .Z(n883) );
  NAND2X0 U815 ( .IN1(N81), .IN2(n826), .QN(n872) );
  NAND2X0 U816 ( .IN1(n911), .IN2(n1041), .QN(n873) );
  NAND2X0 U817 ( .IN1(n929), .IN2(n614), .QN(n874) );
  NAND3X0 U818 ( .IN1(n874), .IN2(n873), .IN3(n872), .QN(N231) );
  NAND2X1 U819 ( .IN1(n894), .IN2(n893), .QN(n1024) );
  NAND2X0 U820 ( .IN1(N82), .IN2(n826), .QN(n875) );
  NAND2X0 U821 ( .IN1(n899), .IN2(n1042), .QN(n876) );
  NAND2X0 U822 ( .IN1(n884), .IN2(n615), .QN(n877) );
  NAND3X0 U823 ( .IN1(n875), .IN2(n876), .IN3(n877), .QN(N230) );
  NAND2X0 U824 ( .IN1(n883), .IN2(N103), .QN(n878) );
  NAND2X0 U825 ( .IN1(n797), .IN2(A_reg[27]), .QN(n879) );
  NAND2X0 U826 ( .IN1(n785), .IN2(n671), .QN(n880) );
  NAND3X0 U827 ( .IN1(n878), .IN2(n879), .IN3(n880), .QN(N209) );
  NAND4X0 U828 ( .IN1(n1008), .IN2(n1007), .IN3(n1006), .IN4(n1005), .QN(n887)
         );
  INVX0 U829 ( .INP(n890), .ZN(n891) );
  INVX0 U830 ( .INP(n895), .ZN(n896) );
  NAND2X0 U831 ( .IN1(n889), .IN2(n914), .QN(n1020) );
  INVX0 U832 ( .INP(n955), .ZN(n953) );
  INVX0 U833 ( .INP(n955), .ZN(n952) );
  INVX0 U834 ( .INP(n900), .ZN(n924) );
  NBUFFX2 U835 ( .INP(n903), .Z(n920) );
  NBUFFX2 U836 ( .INP(n906), .Z(n928) );
  AND2X1 U837 ( .IN1(n943), .IN2(n977), .Q(n900) );
  INVX0 U838 ( .INP(n977), .ZN(n966) );
  INVX0 U839 ( .INP(n978), .ZN(n965) );
  INVX0 U840 ( .INP(n977), .ZN(n967) );
  INVX0 U841 ( .INP(n977), .ZN(n964) );
  INVX0 U842 ( .INP(n977), .ZN(n969) );
  INVX0 U843 ( .INP(n976), .ZN(n968) );
  INVX0 U844 ( .INP(n977), .ZN(n963) );
  NOR2X0 U845 ( .IN1(counter[5]), .IN2(n1022), .QN(n1011) );
  NOR2X0 U846 ( .IN1(counter[8]), .IN2(counter[9]), .QN(n1006) );
  NOR2X0 U847 ( .IN1(n1000), .IN2(n1001), .QN(n1008) );
  AND4X1 U848 ( .IN1(n1027), .IN2(n1028), .IN3(n642), .IN4(n622), .Q(n901) );
  NOR2X0 U849 ( .IN1(n1002), .IN2(n1003), .QN(n996) );
  NBUFFX2 U850 ( .INP(n907), .Z(n917) );
  AND2X1 U851 ( .IN1(n955), .IN2(n1052), .Q(n904) );
  INVX0 U852 ( .INP(n909), .ZN(n946) );
  INVX0 U853 ( .INP(n909), .ZN(n945) );
  INVX0 U854 ( .INP(n961), .ZN(n977) );
  AND2X1 U855 ( .IN1(n955), .IN2(n1053), .Q(n905) );
  NBUFFX2 U856 ( .INP(n910), .Z(n923) );
  AND2X1 U857 ( .IN1(n900), .IN2(A_reg[31]), .Q(n906) );
  INVX0 U858 ( .INP(n961), .ZN(n976) );
  INVX0 U859 ( .INP(n962), .ZN(n978) );
  NOR2X0 U860 ( .IN1(n970), .IN2(n1051), .QN(N72) );
  INVX0 U861 ( .INP(n962), .ZN(n984) );
  INVX0 U862 ( .INP(n962), .ZN(n985) );
  INVX0 U863 ( .INP(n962), .ZN(n986) );
  INVX0 U864 ( .INP(n962), .ZN(n983) );
  INVX0 U865 ( .INP(n962), .ZN(n979) );
  INVX0 U866 ( .INP(n962), .ZN(n980) );
  INVX0 U867 ( .INP(n962), .ZN(n981) );
  INVX0 U868 ( .INP(n962), .ZN(n982) );
  INVX0 U869 ( .INP(n962), .ZN(n987) );
  INVX0 U870 ( .INP(n961), .ZN(n974) );
  INVX0 U871 ( .INP(n961), .ZN(n975) );
  INVX0 U872 ( .INP(n961), .ZN(n973) );
  INVX0 U873 ( .INP(n961), .ZN(n971) );
  INVX0 U874 ( .INP(n961), .ZN(n972) );
  NOR2X0 U875 ( .IN1(n428), .IN2(n938), .QN(N849) );
  NOR2X0 U876 ( .IN1(n429), .IN2(n938), .QN(N847) );
  NOR2X0 U877 ( .IN1(n414), .IN2(n934), .QN(N877) );
  NOR2X0 U878 ( .IN1(n1015), .IN2(n1014), .QN(n1018) );
  NOR2X0 U879 ( .IN1(n430), .IN2(n939), .QN(N845) );
  NOR2X0 U880 ( .IN1(n427), .IN2(n937), .QN(N851) );
  NOR2X0 U881 ( .IN1(n434), .IN2(n941), .QN(N837) );
  NOR2X0 U882 ( .IN1(n420), .IN2(n935), .QN(N865) );
  NOR2X0 U883 ( .IN1(n426), .IN2(n937), .QN(N853) );
  NOR2X0 U884 ( .IN1(n433), .IN2(n940), .QN(N839) );
  NOR2X0 U885 ( .IN1(n419), .IN2(n935), .QN(N867) );
  NOR2X0 U886 ( .IN1(n418), .IN2(n935), .QN(N869) );
  NOR2X0 U887 ( .IN1(n431), .IN2(n939), .QN(N843) );
  NOR2X0 U888 ( .IN1(n432), .IN2(n940), .QN(N841) );
  NOR2X0 U889 ( .IN1(n412), .IN2(n934), .QN(N881) );
  NOR2X0 U890 ( .IN1(n422), .IN2(n936), .QN(N861) );
  NOR2X0 U891 ( .IN1(n411), .IN2(n933), .QN(N883) );
  NOR2X0 U892 ( .IN1(n413), .IN2(n940), .QN(N879) );
  NOR2X0 U893 ( .IN1(n410), .IN2(n933), .QN(N885) );
  NOR2X0 U894 ( .IN1(n409), .IN2(n932), .QN(N887) );
  NOR2X0 U895 ( .IN1(n415), .IN2(n937), .QN(N875) );
  NOR2X0 U896 ( .IN1(n425), .IN2(n939), .QN(N855) );
  NOR2X0 U897 ( .IN1(n424), .IN2(n938), .QN(N857) );
  NOR2X0 U898 ( .IN1(n423), .IN2(n939), .QN(N859) );
  NOR2X0 U899 ( .IN1(n417), .IN2(n936), .QN(N871) );
  NOR2X0 U900 ( .IN1(n416), .IN2(n935), .QN(N873) );
  NOR2X0 U901 ( .IN1(n600), .IN2(n820), .QN(n1016) );
  NAND2X0 U902 ( .IN1(n989), .IN2(n988), .QN(n990) );
  NAND2X0 U903 ( .IN1(n238), .IN2(n235), .QN(n1001) );
  AND2X1 U904 ( .IN1(n401), .IN2(n942), .Q(n907) );
  NOR2X0 U905 ( .IN1(n1029), .IN2(counter[18]), .QN(n995) );
  INVX0 U906 ( .INP(n240), .ZN(n1034) );
  NAND2X0 U907 ( .IN1(n240), .IN2(n242), .QN(n1004) );
  INVX0 U908 ( .INP(n403), .ZN(n1022) );
  NOR4X0 U909 ( .IN1(n1031), .IN2(n1033), .IN3(n1032), .IN4(counter[31]), .QN(
        n908) );
  INVX0 U910 ( .INP(n1029), .ZN(n1030) );
  NOR2X0 U911 ( .IN1(n436), .IN2(n941), .QN(N833) );
  NOR2X0 U912 ( .IN1(n437), .IN2(n941), .QN(N831) );
  NOR2X0 U913 ( .IN1(n438), .IN2(n942), .QN(N829) );
  NOR2X0 U914 ( .IN1(n435), .IN2(n941), .QN(N835) );
  MUX21X1 U915 ( .IN1(n870), .IN2(n684), .S(n965), .Q(n585) );
  INVX0 U916 ( .INP(n394), .ZN(n1038) );
  INVX0 U917 ( .INP(n390), .ZN(n1040) );
  INVX0 U918 ( .INP(n398), .ZN(n1036) );
  INVX0 U919 ( .INP(n370), .ZN(n1048) );
  INVX0 U920 ( .INP(n396), .ZN(n1037) );
  INVX0 U921 ( .INP(n392), .ZN(n1039) );
  INVX0 U922 ( .INP(n386), .ZN(n1042) );
  INVX0 U923 ( .INP(n384), .ZN(n1043) );
  INVX0 U924 ( .INP(n388), .ZN(n1041) );
  INVX0 U925 ( .INP(n382), .ZN(n1044) );
  INVX0 U926 ( .INP(n380), .ZN(n1045) );
  INVX0 U927 ( .INP(n376), .ZN(n1047) );
  INVX0 U928 ( .INP(n368), .ZN(n1049) );
  INVX0 U929 ( .INP(n378), .ZN(n1046) );
  NBUFFX2 U930 ( .INP(rst), .Z(n961) );
  AND2X1 U931 ( .IN1(n399), .IN2(n900), .Q(n910) );
  NBUFFX2 U932 ( .INP(rst), .Z(n962) );
  INVX0 U933 ( .INP(B[31]), .ZN(n1051) );
  NOR2X0 U934 ( .IN1(n292), .IN2(n969), .QN(N547) );
  NOR2X0 U935 ( .IN1(n291), .IN2(n969), .QN(N548) );
  NOR2X0 U936 ( .IN1(n290), .IN2(n969), .QN(N549) );
  NOR2X0 U937 ( .IN1(n289), .IN2(n969), .QN(N550) );
  NOR2X0 U938 ( .IN1(n288), .IN2(n969), .QN(N551) );
  NOR2X0 U939 ( .IN1(n287), .IN2(n969), .QN(N552) );
  NOR2X0 U940 ( .IN1(n286), .IN2(n969), .QN(N553) );
  NOR2X0 U941 ( .IN1(n285), .IN2(n969), .QN(N554) );
  NOR2X0 U942 ( .IN1(n284), .IN2(n969), .QN(N555) );
  NOR2X0 U943 ( .IN1(n283), .IN2(n969), .QN(N556) );
  NOR2X0 U944 ( .IN1(n282), .IN2(n969), .QN(N557) );
  NOR2X0 U945 ( .IN1(n281), .IN2(n969), .QN(N558) );
  NOR2X0 U946 ( .IN1(n280), .IN2(n969), .QN(N559) );
  NOR2X0 U947 ( .IN1(n279), .IN2(n969), .QN(N560) );
  NOR2X0 U948 ( .IN1(n278), .IN2(n969), .QN(N561) );
  NOR2X0 U949 ( .IN1(n243), .IN2(n969), .QN(N562) );
  NOR2X0 U950 ( .IN1(n277), .IN2(n969), .QN(N563) );
  NOR2X0 U951 ( .IN1(n276), .IN2(n969), .QN(N564) );
  NOR2X0 U952 ( .IN1(n275), .IN2(n969), .QN(N565) );
  NOR2X0 U953 ( .IN1(n274), .IN2(n969), .QN(N566) );
  NOR2X0 U954 ( .IN1(n273), .IN2(n969), .QN(N567) );
  NOR2X0 U955 ( .IN1(n272), .IN2(n968), .QN(N568) );
  NOR2X0 U956 ( .IN1(n271), .IN2(n968), .QN(N569) );
  NOR2X0 U957 ( .IN1(n270), .IN2(n968), .QN(N570) );
  NOR2X0 U958 ( .IN1(n269), .IN2(n968), .QN(N571) );
  NOR2X0 U959 ( .IN1(n268), .IN2(n968), .QN(N572) );
  NOR2X0 U960 ( .IN1(n267), .IN2(n968), .QN(N573) );
  NOR2X0 U961 ( .IN1(n266), .IN2(n968), .QN(N574) );
  NOR2X0 U962 ( .IN1(n265), .IN2(n968), .QN(N575) );
  NOR2X0 U963 ( .IN1(n264), .IN2(n968), .QN(N576) );
  NOR2X0 U964 ( .IN1(n263), .IN2(n968), .QN(N577) );
  NOR2X0 U965 ( .IN1(n262), .IN2(n968), .QN(N578) );
  NOR2X0 U966 ( .IN1(n261), .IN2(n968), .QN(N579) );
  NOR2X0 U967 ( .IN1(n260), .IN2(n968), .QN(N580) );
  NOR2X0 U968 ( .IN1(n259), .IN2(n968), .QN(N581) );
  NOR2X0 U969 ( .IN1(n258), .IN2(n968), .QN(N582) );
  NOR2X0 U970 ( .IN1(n257), .IN2(n968), .QN(N583) );
  NOR2X0 U971 ( .IN1(n256), .IN2(n968), .QN(N584) );
  NOR2X0 U972 ( .IN1(n255), .IN2(n968), .QN(N585) );
  NOR2X0 U973 ( .IN1(n254), .IN2(n968), .QN(N586) );
  NOR2X0 U974 ( .IN1(n253), .IN2(n968), .QN(N587) );
  NOR2X0 U975 ( .IN1(n244), .IN2(n968), .QN(N596) );
  NOR2X0 U976 ( .IN1(n252), .IN2(n967), .QN(N588) );
  NOR2X0 U977 ( .IN1(n251), .IN2(n967), .QN(N589) );
  NOR2X0 U978 ( .IN1(n250), .IN2(n967), .QN(N590) );
  NOR2X0 U979 ( .IN1(n249), .IN2(n967), .QN(N591) );
  NOR2X0 U980 ( .IN1(n248), .IN2(n967), .QN(N592) );
  NOR2X0 U981 ( .IN1(n247), .IN2(n967), .QN(N593) );
  NOR2X0 U982 ( .IN1(n246), .IN2(n967), .QN(N594) );
  NOR2X0 U983 ( .IN1(n245), .IN2(n967), .QN(N595) );
  NOR2X0 U984 ( .IN1(n964), .IN2(n294), .QN(N545) );
  NOR2X0 U985 ( .IN1(n963), .IN2(n306), .QN(N533) );
  NOR2X0 U986 ( .IN1(n963), .IN2(n305), .QN(N534) );
  NOR2X0 U987 ( .IN1(n963), .IN2(n304), .QN(N535) );
  NOR2X0 U988 ( .IN1(n963), .IN2(n303), .QN(N536) );
  NOR2X0 U989 ( .IN1(n963), .IN2(n302), .QN(N537) );
  NOR2X0 U990 ( .IN1(n963), .IN2(n301), .QN(N538) );
  NOR2X0 U991 ( .IN1(n963), .IN2(n300), .QN(N539) );
  NOR2X0 U992 ( .IN1(n963), .IN2(n299), .QN(N540) );
  NOR2X0 U993 ( .IN1(n963), .IN2(n298), .QN(N541) );
  NOR2X0 U994 ( .IN1(n963), .IN2(n297), .QN(N542) );
  NOR2X0 U995 ( .IN1(n963), .IN2(n296), .QN(N543) );
  NOR2X0 U996 ( .IN1(n963), .IN2(n295), .QN(N544) );
  NOR2X0 U997 ( .IN1(n293), .IN2(n970), .QN(N546) );
  NOR2X0 U998 ( .IN1(n970), .IN2(n1019), .QN(N40) );
  INVX0 U999 ( .INP(A[31]), .ZN(n1019) );
  INVX0 U1000 ( .INP(n1035), .ZN(n912) );
  NOR4X0 U1001 ( .IN1(n1023), .IN2(n1025), .IN3(n1024), .IN4(n1026), .QN(n1027) );
  AND4X1 U1002 ( .IN1(n233), .IN2(n241), .IN3(n234), .IN4(n236), .Q(n913) );
  INVX0 U1003 ( .INP(n1025), .ZN(n1007) );
  NAND2X0 U1004 ( .IN1(n406), .IN2(n405), .QN(n1021) );
  NOR2X0 U1005 ( .IN1(counter[25]), .IN2(counter[28]), .QN(n988) );
  NOR2X0 U1006 ( .IN1(counter[29]), .IN2(n1034), .QN(n989) );
  NOR2X0 U1007 ( .IN1(n990), .IN2(n869), .QN(n993) );
  NOR2X0 U1008 ( .IN1(n865), .IN2(counter[24]), .QN(n994) );
  NOR2X0 U1009 ( .IN1(n1023), .IN2(n1020), .QN(n1010) );
  NOR2X0 U1010 ( .IN1(B_reg[31]), .IN2(B_reg[0]), .QN(n1015) );
  NOR2X0 U1011 ( .IN1(n401), .IN2(N141), .QN(n1014) );
  NOR2X0 U1012 ( .IN1(counter[13]), .IN2(n1024), .QN(n991) );
  NOR2X0 U1013 ( .IN1(n1026), .IN2(n1024), .QN(n1009) );
  NBUFFX2 U1014 ( .INP(n907), .Z(n915) );
  NBUFFX2 U1015 ( .INP(n903), .Z(n919) );
  NBUFFX2 U1016 ( .INP(n910), .Z(n921) );
  NBUFFX2 U1017 ( .INP(n910), .Z(n922) );
  NBUFFX2 U1018 ( .INP(n906), .Z(n926) );
  NBUFFX2 U1019 ( .INP(n906), .Z(n927) );
  NBUFFX2 U1020 ( .INP(n902), .Z(n944) );
  NBUFFX2 U1021 ( .INP(n905), .Z(n947) );
  NBUFFX2 U1022 ( .INP(n905), .Z(n948) );
  NBUFFX2 U1023 ( .INP(n905), .Z(n949) );
  NBUFFX2 U1024 ( .INP(n905), .Z(n950) );
  NBUFFX2 U1025 ( .INP(n905), .Z(n951) );
  NBUFFX2 U1026 ( .INP(n904), .Z(n956) );
  NBUFFX2 U1027 ( .INP(n904), .Z(n957) );
  NBUFFX2 U1028 ( .INP(n904), .Z(n958) );
  INVX0 U1029 ( .INP(n900), .ZN(n925) );
  INVX0 U1030 ( .INP(n930), .ZN(n932) );
  INVX0 U1031 ( .INP(n930), .ZN(n933) );
  INVX0 U1032 ( .INP(n930), .ZN(n934) );
  INVX0 U1033 ( .INP(n931), .ZN(n935) );
  INVX0 U1034 ( .INP(n931), .ZN(n936) );
  INVX0 U1035 ( .INP(n931), .ZN(n937) );
  INVX0 U1036 ( .INP(n930), .ZN(n938) );
  INVX0 U1037 ( .INP(n930), .ZN(n939) );
  INVX0 U1038 ( .INP(n930), .ZN(n940) );
  INVX0 U1039 ( .INP(n931), .ZN(n941) );
  INVX0 U1040 ( .INP(n929), .ZN(n942) );
  INVX0 U1041 ( .INP(n929), .ZN(n943) );
  INVX0 U1042 ( .INP(n1054), .ZN(n955) );
  INVX0 U1043 ( .INP(n978), .ZN(n970) );
  NOR3X0 U1044 ( .IN1(counter[11]), .IN2(n866), .IN3(counter[7]), .QN(n992) );
  NAND4X0 U1045 ( .IN1(n993), .IN2(n994), .IN3(n992), .IN4(n991), .QN(n998) );
  NAND4X0 U1046 ( .IN1(n228), .IN2(n230), .IN3(n239), .IN4(n229), .QN(n1002)
         );
  NAND4X0 U1047 ( .IN1(n996), .IN2(n242), .IN3(n635), .IN4(n995), .QN(n997) );
  AND2X1 U1048 ( .IN1(N470), .IN2(n945), .Q(N502) );
  AND2X1 U1049 ( .IN1(N473), .IN2(n945), .Q(N505) );
  AND2X1 U1050 ( .IN1(N474), .IN2(n945), .Q(N506) );
  AND2X1 U1051 ( .IN1(N475), .IN2(n945), .Q(N507) );
  AND2X1 U1052 ( .IN1(N477), .IN2(n945), .Q(N509) );
  AND2X1 U1053 ( .IN1(N482), .IN2(n945), .Q(N514) );
  AND2X1 U1054 ( .IN1(N483), .IN2(n945), .Q(N515) );
  AND2X1 U1055 ( .IN1(N484), .IN2(n945), .Q(N516) );
  AND2X1 U1056 ( .IN1(N486), .IN2(n945), .Q(N518) );
  AND2X1 U1057 ( .IN1(N487), .IN2(n945), .Q(N519) );
  AND2X1 U1058 ( .IN1(N488), .IN2(n945), .Q(N520) );
  AND2X1 U1059 ( .IN1(N491), .IN2(n945), .Q(N523) );
  AND2X1 U1060 ( .IN1(N492), .IN2(n946), .Q(N524) );
  AND2X1 U1061 ( .IN1(N495), .IN2(n946), .Q(N527) );
  AND2X1 U1062 ( .IN1(N494), .IN2(n946), .Q(N526) );
  AND2X1 U1063 ( .IN1(N493), .IN2(n946), .Q(N525) );
  AND2X1 U1064 ( .IN1(N490), .IN2(n946), .Q(N522) );
  AND2X1 U1065 ( .IN1(N489), .IN2(n946), .Q(N521) );
  AND2X1 U1066 ( .IN1(N485), .IN2(n946), .Q(N517) );
  AND2X1 U1067 ( .IN1(N481), .IN2(n946), .Q(N513) );
  AND2X1 U1068 ( .IN1(N480), .IN2(n946), .Q(N512) );
  AND2X1 U1069 ( .IN1(N479), .IN2(n946), .Q(N511) );
  AND2X1 U1070 ( .IN1(N478), .IN2(n946), .Q(N510) );
  AND2X1 U1071 ( .IN1(N476), .IN2(n946), .Q(N508) );
  AND2X1 U1072 ( .IN1(N472), .IN2(n945), .Q(N504) );
  AND2X1 U1073 ( .IN1(N471), .IN2(n946), .Q(N503) );
  AND2X1 U1074 ( .IN1(N469), .IN2(n945), .Q(N501) );
  AND2X1 U1075 ( .IN1(N468), .IN2(n946), .Q(N500) );
  AND2X1 U1076 ( .IN1(N467), .IN2(n945), .Q(N499) );
  AND2X1 U1077 ( .IN1(N466), .IN2(n946), .Q(N498) );
  AND2X1 U1078 ( .IN1(N496), .IN2(n945), .Q(N528) );
  AND2X1 U1079 ( .IN1(N465), .IN2(n946), .Q(N497) );
  AND2X1 U1080 ( .IN1(B[1]), .IN2(n978), .Q(N42) );
  AND2X1 U1081 ( .IN1(B[30]), .IN2(n987), .Q(N71) );
  AND2X1 U1082 ( .IN1(B[29]), .IN2(n987), .Q(N70) );
  AND2X1 U1083 ( .IN1(B[28]), .IN2(n986), .Q(N69) );
  AND2X1 U1084 ( .IN1(B[27]), .IN2(n986), .Q(N68) );
  AND2X1 U1085 ( .IN1(B[26]), .IN2(n986), .Q(N67) );
  AND2X1 U1086 ( .IN1(B[25]), .IN2(n986), .Q(N66) );
  AND2X1 U1087 ( .IN1(B[24]), .IN2(n986), .Q(N65) );
  AND2X1 U1088 ( .IN1(B[23]), .IN2(n986), .Q(N64) );
  AND2X1 U1089 ( .IN1(B[22]), .IN2(n986), .Q(N63) );
  AND2X1 U1090 ( .IN1(B[21]), .IN2(n985), .Q(N62) );
  AND2X1 U1091 ( .IN1(B[20]), .IN2(n985), .Q(N61) );
  AND2X1 U1092 ( .IN1(B[19]), .IN2(n985), .Q(N60) );
  AND2X1 U1093 ( .IN1(B[18]), .IN2(n985), .Q(N59) );
  AND2X1 U1094 ( .IN1(B[17]), .IN2(n985), .Q(N58) );
  AND2X1 U1095 ( .IN1(B[16]), .IN2(n985), .Q(N57) );
  AND2X1 U1096 ( .IN1(B[15]), .IN2(n985), .Q(N56) );
  AND2X1 U1097 ( .IN1(B[14]), .IN2(n984), .Q(N55) );
  AND2X1 U1098 ( .IN1(B[13]), .IN2(n980), .Q(N54) );
  AND2X1 U1099 ( .IN1(B[12]), .IN2(n984), .Q(N53) );
  AND2X1 U1100 ( .IN1(B[11]), .IN2(n984), .Q(N52) );
  AND2X1 U1101 ( .IN1(B[10]), .IN2(n984), .Q(N51) );
  AND2X1 U1102 ( .IN1(B[9]), .IN2(n984), .Q(N50) );
  AND2X1 U1103 ( .IN1(B[8]), .IN2(n984), .Q(N49) );
  AND2X1 U1104 ( .IN1(B[7]), .IN2(n984), .Q(N48) );
  AND2X1 U1105 ( .IN1(B[6]), .IN2(n983), .Q(N47) );
  AND2X1 U1106 ( .IN1(B[5]), .IN2(n983), .Q(N46) );
  AND2X1 U1107 ( .IN1(B[4]), .IN2(n983), .Q(N45) );
  AND2X1 U1108 ( .IN1(B[3]), .IN2(n983), .Q(N44) );
  AND2X1 U1109 ( .IN1(B[2]), .IN2(n983), .Q(N43) );
  AND2X1 U1110 ( .IN1(B[0]), .IN2(n983), .Q(N41) );
  MUX21X1 U1111 ( .IN1(N334), .IN2(n685), .S(n964), .Q(n597) );
  NOR3X0 U1112 ( .IN1(n795), .IN2(n1003), .IN3(n1004), .QN(n1005) );
  NAND4X0 U1113 ( .IN1(n793), .IN2(n1009), .IN3(n1010), .IN4(n1011), .QN(n1012) );
  MUX21X1 U1114 ( .IN1(N331), .IN2(n686), .S(n964), .Q(n594) );
  MUX21X1 U1115 ( .IN1(n812), .IN2(n687), .S(n964), .Q(n593) );
  MUX21X1 U1116 ( .IN1(n845), .IN2(n688), .S(n964), .Q(n592) );
  MUX21X1 U1117 ( .IN1(N327), .IN2(n689), .S(n964), .Q(n590) );
  MUX21X1 U1118 ( .IN1(N326), .IN2(n690), .S(n964), .Q(n589) );
  MUX21X1 U1119 ( .IN1(N324), .IN2(n691), .S(n964), .Q(n587) );
  MUX21X1 U1120 ( .IN1(N320), .IN2(n692), .S(n964), .Q(n583) );
  MUX21X1 U1121 ( .IN1(N319), .IN2(n693), .S(n965), .Q(n582) );
  MUX21X1 U1122 ( .IN1(n829), .IN2(n682), .S(n964), .Q(n580) );
  MUX21X1 U1123 ( .IN1(n799), .IN2(n694), .S(n965), .Q(n579) );
  MUX21X1 U1124 ( .IN1(n805), .IN2(n695), .S(n964), .Q(n577) );
  MUX21X1 U1125 ( .IN1(N313), .IN2(n696), .S(n965), .Q(n576) );
  MUX21X1 U1126 ( .IN1(N311), .IN2(n697), .S(n965), .Q(n574) );
  MUX21X1 U1127 ( .IN1(n802), .IN2(n698), .S(n965), .Q(n573) );
  MUX21X1 U1128 ( .IN1(N309), .IN2(n699), .S(n965), .Q(n572) );
  MUX21X1 U1129 ( .IN1(N308), .IN2(n700), .S(n965), .Q(n571) );
  MUX21X1 U1130 ( .IN1(N307), .IN2(n701), .S(n965), .Q(n570) );
  MUX21X1 U1131 ( .IN1(N306), .IN2(n702), .S(n965), .Q(n569) );
  MUX21X1 U1132 ( .IN1(N305), .IN2(n703), .S(n965), .Q(n568) );
  MUX21X1 U1133 ( .IN1(N304), .IN2(n683), .S(n966), .Q(n567) );
  MUX21X1 U1134 ( .IN1(N303), .IN2(n661), .S(n965), .Q(n598) );
  AO22X1 U1135 ( .IN1(n783), .IN2(n661), .IN3(N172), .IN4(n918), .Q(N237) );
  AO222X1 U1136 ( .IN1(N171), .IN2(n918), .IN3(B_reg[30]), .IN4(n917), .IN5(
        n782), .IN6(n659), .Q(N238) );
  AO222X1 U1137 ( .IN1(N170), .IN2(n918), .IN3(B_reg[29]), .IN4(n917), .IN5(
        n785), .IN6(n672), .Q(N239) );
  MUX21X1 U1138 ( .IN1(N239), .IN2(n643), .S(n965), .Q(n532) );
  AO222X1 U1139 ( .IN1(N169), .IN2(n918), .IN3(B_reg[28]), .IN4(n917), .IN5(
        n781), .IN6(n643), .Q(N240) );
  MUX21X1 U1140 ( .IN1(N240), .IN2(n644), .S(n965), .Q(n531) );
  AO222X1 U1141 ( .IN1(N168), .IN2(n918), .IN3(B_reg[27]), .IN4(n917), .IN5(
        n779), .IN6(n644), .Q(N241) );
  MUX21X1 U1142 ( .IN1(N241), .IN2(n645), .S(n966), .Q(n530) );
  AO222X1 U1143 ( .IN1(N167), .IN2(n918), .IN3(B_reg[26]), .IN4(n917), .IN5(
        n786), .IN6(n645), .Q(N242) );
  MUX21X1 U1144 ( .IN1(N242), .IN2(n646), .S(n966), .Q(n529) );
  AO222X1 U1145 ( .IN1(N166), .IN2(n918), .IN3(B_reg[25]), .IN4(n917), .IN5(
        n777), .IN6(n646), .Q(N243) );
  MUX21X1 U1146 ( .IN1(N243), .IN2(n623), .S(n965), .Q(n528) );
  AO222X1 U1147 ( .IN1(N165), .IN2(n918), .IN3(B_reg[24]), .IN4(n916), .IN5(
        n776), .IN6(n623), .Q(N244) );
  MUX21X1 U1148 ( .IN1(N244), .IN2(n647), .S(n966), .Q(n527) );
  AO222X1 U1149 ( .IN1(N164), .IN2(n918), .IN3(B_reg[23]), .IN4(n916), .IN5(
        n788), .IN6(n647), .Q(N245) );
  MUX21X1 U1150 ( .IN1(N245), .IN2(n648), .S(n966), .Q(n526) );
  AO222X1 U1151 ( .IN1(N163), .IN2(n918), .IN3(B_reg[22]), .IN4(n916), .IN5(
        n778), .IN6(n648), .Q(N246) );
  MUX21X1 U1152 ( .IN1(N246), .IN2(n649), .S(n966), .Q(n525) );
  AO222X1 U1153 ( .IN1(N162), .IN2(n918), .IN3(B_reg[21]), .IN4(n916), .IN5(
        n788), .IN6(n649), .Q(N247) );
  MUX21X1 U1154 ( .IN1(N247), .IN2(n624), .S(n966), .Q(n524) );
  AO222X1 U1155 ( .IN1(N161), .IN2(n918), .IN3(B_reg[20]), .IN4(n916), .IN5(
        n780), .IN6(n624), .Q(N248) );
  MUX21X1 U1156 ( .IN1(N248), .IN2(n650), .S(n966), .Q(n523) );
  AO222X1 U1157 ( .IN1(N160), .IN2(n918), .IN3(B_reg[19]), .IN4(n916), .IN5(
        n782), .IN6(n650), .Q(N249) );
  MUX21X1 U1158 ( .IN1(N249), .IN2(n651), .S(n966), .Q(n522) );
  AO222X1 U1159 ( .IN1(N159), .IN2(n919), .IN3(B_reg[18]), .IN4(n916), .IN5(
        n783), .IN6(n651), .Q(N250) );
  MUX21X1 U1160 ( .IN1(N250), .IN2(n790), .S(n966), .Q(n521) );
  MUX21X1 U1161 ( .IN1(n602), .IN2(n625), .S(n966), .Q(n520) );
  AO222X1 U1162 ( .IN1(N157), .IN2(n919), .IN3(B_reg[16]), .IN4(n916), .IN5(
        n782), .IN6(n625), .Q(N252) );
  MUX21X1 U1163 ( .IN1(N252), .IN2(n652), .S(n966), .Q(n519) );
  AO222X1 U1164 ( .IN1(N156), .IN2(n919), .IN3(B_reg[15]), .IN4(n916), .IN5(
        n778), .IN6(n652), .Q(N253) );
  MUX21X1 U1165 ( .IN1(N253), .IN2(n653), .S(n967), .Q(n518) );
  AO222X1 U1166 ( .IN1(N155), .IN2(n919), .IN3(B_reg[14]), .IN4(n916), .IN5(
        n786), .IN6(n653), .Q(N254) );
  MUX21X1 U1167 ( .IN1(N254), .IN2(n654), .S(n966), .Q(n517) );
  AO222X1 U1168 ( .IN1(N154), .IN2(n919), .IN3(B_reg[13]), .IN4(n916), .IN5(
        n785), .IN6(n654), .Q(N255) );
  MUX21X1 U1169 ( .IN1(N255), .IN2(n626), .S(n966), .Q(n516) );
  AO222X1 U1170 ( .IN1(N153), .IN2(n919), .IN3(B_reg[12]), .IN4(n915), .IN5(
        n784), .IN6(n626), .Q(N256) );
  MUX21X1 U1171 ( .IN1(N256), .IN2(n655), .S(n967), .Q(n515) );
  AO222X1 U1172 ( .IN1(N152), .IN2(n919), .IN3(B_reg[11]), .IN4(n915), .IN5(
        n780), .IN6(n655), .Q(N257) );
  MUX21X1 U1173 ( .IN1(N257), .IN2(n656), .S(n966), .Q(n514) );
  AO222X1 U1174 ( .IN1(N151), .IN2(n919), .IN3(B_reg[10]), .IN4(n915), .IN5(
        n787), .IN6(n656), .Q(N258) );
  AO222X1 U1175 ( .IN1(N150), .IN2(n919), .IN3(B_reg[9]), .IN4(n915), .IN5(
        n782), .IN6(n660), .Q(N259) );
  MUX21X1 U1176 ( .IN1(N259), .IN2(n627), .S(n967), .Q(n512) );
  AO222X1 U1177 ( .IN1(N149), .IN2(n919), .IN3(B_reg[8]), .IN4(n915), .IN5(
        n777), .IN6(n627), .Q(N260) );
  MUX21X1 U1178 ( .IN1(N260), .IN2(n657), .S(n966), .Q(n511) );
  AO222X1 U1179 ( .IN1(N148), .IN2(n919), .IN3(B_reg[7]), .IN4(n915), .IN5(
        n781), .IN6(n657), .Q(N261) );
  MUX21X1 U1180 ( .IN1(N261), .IN2(n789), .S(n966), .Q(n510) );
  MUX21X1 U1181 ( .IN1(n601), .IN2(n628), .S(n967), .Q(n509) );
  AO222X1 U1182 ( .IN1(N146), .IN2(n920), .IN3(B_reg[5]), .IN4(n915), .IN5(
        n788), .IN6(n628), .Q(N263) );
  MUX21X1 U1183 ( .IN1(N263), .IN2(n604), .S(n967), .Q(n508) );
  AO222X1 U1184 ( .IN1(N145), .IN2(n920), .IN3(B_reg[4]), .IN4(n915), .IN5(
        n776), .IN6(n604), .Q(N264) );
  MUX21X1 U1185 ( .IN1(N264), .IN2(n658), .S(n967), .Q(n507) );
  AO222X1 U1186 ( .IN1(N144), .IN2(n920), .IN3(B_reg[3]), .IN4(n915), .IN5(
        n779), .IN6(n658), .Q(N265) );
  MUX21X1 U1187 ( .IN1(N265), .IN2(n629), .S(n967), .Q(n506) );
  AO222X1 U1188 ( .IN1(N143), .IN2(n920), .IN3(B_reg[2]), .IN4(n915), .IN5(
        n784), .IN6(n629), .Q(N266) );
  MUX21X1 U1189 ( .IN1(N266), .IN2(n630), .S(n967), .Q(n505) );
  AO222X1 U1190 ( .IN1(N142), .IN2(n920), .IN3(B_reg[1]), .IN4(n915), .IN5(
        n783), .IN6(n630), .Q(N267) );
  MUX21X1 U1191 ( .IN1(N267), .IN2(n792), .S(n967), .Q(n504) );
  AND2X1 U1192 ( .IN1(A[0]), .IN2(n983), .Q(N9) );
  AND2X1 U1193 ( .IN1(A[30]), .IN2(n982), .Q(N39) );
  AND2X1 U1194 ( .IN1(A[29]), .IN2(n982), .Q(N38) );
  AND2X1 U1195 ( .IN1(A[28]), .IN2(n982), .Q(N37) );
  AND2X1 U1196 ( .IN1(A[27]), .IN2(n982), .Q(N36) );
  AND2X1 U1197 ( .IN1(A[26]), .IN2(n982), .Q(N35) );
  AND2X1 U1198 ( .IN1(A[25]), .IN2(n982), .Q(N34) );
  AND2X1 U1199 ( .IN1(A[24]), .IN2(n982), .Q(N33) );
  AND2X1 U1200 ( .IN1(A[23]), .IN2(n981), .Q(N32) );
  AND2X1 U1201 ( .IN1(A[22]), .IN2(n981), .Q(N31) );
  AND2X1 U1202 ( .IN1(A[21]), .IN2(n981), .Q(N30) );
  AND2X1 U1203 ( .IN1(A[20]), .IN2(n981), .Q(N29) );
  AND2X1 U1204 ( .IN1(A[19]), .IN2(n981), .Q(N28) );
  AND2X1 U1205 ( .IN1(A[18]), .IN2(n981), .Q(N27) );
  AND2X1 U1206 ( .IN1(A[17]), .IN2(n981), .Q(N26) );
  AND2X1 U1207 ( .IN1(A[16]), .IN2(n980), .Q(N25) );
  AND2X1 U1208 ( .IN1(A[15]), .IN2(n980), .Q(N24) );
  AND2X1 U1209 ( .IN1(A[14]), .IN2(n980), .Q(N23) );
  AND2X1 U1210 ( .IN1(A[13]), .IN2(n980), .Q(N22) );
  AND2X1 U1211 ( .IN1(A[12]), .IN2(n980), .Q(N21) );
  AND2X1 U1212 ( .IN1(A[11]), .IN2(n980), .Q(N20) );
  AND2X1 U1213 ( .IN1(A[10]), .IN2(n979), .Q(N19) );
  AND2X1 U1214 ( .IN1(A[9]), .IN2(n979), .Q(N18) );
  AND2X1 U1215 ( .IN1(A[8]), .IN2(n979), .Q(N17) );
  AND2X1 U1216 ( .IN1(A[7]), .IN2(n979), .Q(N16) );
  AND2X1 U1217 ( .IN1(A[6]), .IN2(n979), .Q(N15) );
  AND2X1 U1218 ( .IN1(A[5]), .IN2(n979), .Q(N14) );
  AND2X1 U1219 ( .IN1(A[4]), .IN2(n979), .Q(N13) );
  AND2X1 U1220 ( .IN1(A[3]), .IN2(n978), .Q(N12) );
  AND2X1 U1221 ( .IN1(A[2]), .IN2(n978), .Q(N11) );
  AND2X1 U1222 ( .IN1(A[1]), .IN2(n978), .Q(N10) );
  AO222X1 U1223 ( .IN1(N76), .IN2(n926), .IN3(n923), .IN4(n1036), .IN5(n924), 
        .IN6(n605), .Q(n565) );
  NAND2X1 U1224 ( .IN1(n242), .IN2(n232), .QN(n1033) );
  NAND4X0 U1225 ( .IN1(n1030), .IN2(n913), .IN3(n230), .IN4(n238), .QN(n1031)
         );
  AO222X1 U1226 ( .IN1(N76), .IN2(n902), .IN3(n911), .IN4(n1036), .IN5(n930), 
        .IN6(n605), .Q(N236) );
  AO222X1 U1227 ( .IN1(N77), .IN2(n926), .IN3(n923), .IN4(n1037), .IN5(n925), 
        .IN6(n612), .Q(n564) );
  AO222X1 U1228 ( .IN1(N78), .IN2(n926), .IN3(n923), .IN4(n1038), .IN5(n924), 
        .IN6(n606), .Q(n563) );
  AO222X1 U1229 ( .IN1(N78), .IN2(n826), .IN3(n911), .IN4(n1038), .IN5(n929), 
        .IN6(n606), .Q(N234) );
  AO222X1 U1230 ( .IN1(N79), .IN2(n926), .IN3(n923), .IN4(n1039), .IN5(n925), 
        .IN6(n607), .Q(n562) );
  AO222X1 U1231 ( .IN1(N79), .IN2(n826), .IN3(n899), .IN4(n1039), .IN5(n884), 
        .IN6(n607), .Q(N233) );
  AO222X1 U1232 ( .IN1(N80), .IN2(n926), .IN3(n923), .IN4(n1040), .IN5(n924), 
        .IN6(n613), .Q(n561) );
  AO222X1 U1233 ( .IN1(N81), .IN2(n926), .IN3(n923), .IN4(n1041), .IN5(n925), 
        .IN6(n614), .Q(n560) );
  AO222X1 U1234 ( .IN1(N82), .IN2(n926), .IN3(n923), .IN4(n1042), .IN5(n925), 
        .IN6(n615), .Q(n559) );
  AO222X1 U1235 ( .IN1(N83), .IN2(n926), .IN3(n922), .IN4(n1043), .IN5(n924), 
        .IN6(n608), .Q(n558) );
  AO222X1 U1236 ( .IN1(N83), .IN2(n902), .IN3(n911), .IN4(n1043), .IN5(n884), 
        .IN6(n608), .Q(N229) );
  AO222X1 U1237 ( .IN1(N84), .IN2(n926), .IN3(n922), .IN4(n1044), .IN5(n925), 
        .IN6(n609), .Q(n557) );
  AO222X1 U1238 ( .IN1(N84), .IN2(n902), .IN3(n912), .IN4(n1044), .IN5(n931), 
        .IN6(n609), .Q(N228) );
  AO222X1 U1239 ( .IN1(n926), .IN2(N85), .IN3(n922), .IN4(n1045), .IN5(n925), 
        .IN6(n610), .Q(n556) );
  AO222X1 U1240 ( .IN1(N85), .IN2(n826), .IN3(n911), .IN4(n1045), .IN5(n931), 
        .IN6(n610), .Q(N227) );
  AO222X1 U1241 ( .IN1(N86), .IN2(n926), .IN3(n922), .IN4(n1046), .IN5(n925), 
        .IN6(n611), .Q(n555) );
  AO222X1 U1242 ( .IN1(N87), .IN2(n926), .IN3(n922), .IN4(n1047), .IN5(n925), 
        .IN6(n603), .Q(n554) );
  AO222X1 U1243 ( .IN1(N87), .IN2(n902), .IN3(n899), .IN4(n1047), .IN5(n776), 
        .IN6(n603), .Q(N225) );
  AO222X1 U1244 ( .IN1(N88), .IN2(n927), .IN3(n922), .IN4(A_reg[12]), .IN5(
        n924), .IN6(n631), .Q(n553) );
  AO222X1 U1245 ( .IN1(N88), .IN2(n902), .IN3(n772), .IN4(A_reg[12]), .IN5(
        n884), .IN6(n631), .Q(N224) );
  AO222X1 U1246 ( .IN1(N89), .IN2(n927), .IN3(n922), .IN4(A_reg[13]), .IN5(
        n924), .IN6(n616), .Q(n552) );
  AO222X1 U1247 ( .IN1(N90), .IN2(n927), .IN3(n922), .IN4(n1048), .IN5(n924), 
        .IN6(n617), .Q(n551) );
  AO222X1 U1248 ( .IN1(N91), .IN2(n927), .IN3(n922), .IN4(n1049), .IN5(n924), 
        .IN6(n618), .Q(n550) );
  AO222X1 U1249 ( .IN1(N92), .IN2(n927), .IN3(n922), .IN4(A_reg[16]), .IN5(
        n924), .IN6(n632), .Q(n549) );
  AO222X1 U1250 ( .IN1(N92), .IN2(n826), .IN3(n911), .IN4(A_reg[16]), .IN5(
        n931), .IN6(n632), .Q(N220) );
  AO222X1 U1251 ( .IN1(N93), .IN2(n927), .IN3(n922), .IN4(A_reg[17]), .IN5(
        n924), .IN6(n619), .Q(n548) );
  AO222X1 U1252 ( .IN1(N94), .IN2(n927), .IN3(n922), .IN4(A_reg[18]), .IN5(
        n924), .IN6(n633), .Q(n547) );
  AO222X1 U1253 ( .IN1(N94), .IN2(n826), .IN3(n772), .IN4(A_reg[18]), .IN5(
        n778), .IN6(n633), .Q(N218) );
  AO222X1 U1254 ( .IN1(N95), .IN2(n927), .IN3(n921), .IN4(A_reg[19]), .IN5(
        n924), .IN6(n634), .Q(n546) );
  AO222X1 U1255 ( .IN1(N96), .IN2(n927), .IN3(n921), .IN4(A_reg[20]), .IN5(
        n924), .IN6(n662), .Q(n545) );
  AO222X1 U1256 ( .IN1(N96), .IN2(n944), .IN3(n797), .IN4(A_reg[20]), .IN5(
        n930), .IN6(n662), .Q(N216) );
  AO222X1 U1257 ( .IN1(N97), .IN2(n927), .IN3(n921), .IN4(A_reg[21]), .IN5(
        n924), .IN6(n663), .Q(n544) );
  AO222X1 U1258 ( .IN1(N97), .IN2(n883), .IN3(n797), .IN4(A_reg[21]), .IN5(
        n781), .IN6(n663), .Q(N215) );
  AO222X1 U1259 ( .IN1(N98), .IN2(n927), .IN3(n921), .IN4(A_reg[22]), .IN5(
        n924), .IN6(n664), .Q(n543) );
  AO222X1 U1260 ( .IN1(N98), .IN2(n944), .IN3(n797), .IN4(A_reg[22]), .IN5(
        n931), .IN6(n664), .Q(N214) );
  AO222X1 U1261 ( .IN1(N99), .IN2(n927), .IN3(n921), .IN4(A_reg[23]), .IN5(
        n924), .IN6(n665), .Q(n542) );
  AO222X1 U1262 ( .IN1(N99), .IN2(n883), .IN3(n797), .IN4(A_reg[23]), .IN5(
        n786), .IN6(n665), .Q(N213) );
  AO222X1 U1263 ( .IN1(N100), .IN2(n928), .IN3(n921), .IN4(A_reg[24]), .IN5(
        n925), .IN6(n670), .Q(n541) );
  AO222X1 U1264 ( .IN1(N101), .IN2(n928), .IN3(n921), .IN4(A_reg[25]), .IN5(
        n925), .IN6(n666), .Q(n540) );
  AO222X1 U1265 ( .IN1(N101), .IN2(n883), .IN3(n797), .IN4(A_reg[25]), .IN5(
        n931), .IN6(n666), .Q(N211) );
  AO222X1 U1266 ( .IN1(N102), .IN2(n928), .IN3(n921), .IN4(A_reg[26]), .IN5(
        n925), .IN6(n667), .Q(n539) );
  AO222X1 U1267 ( .IN1(N102), .IN2(n883), .IN3(n797), .IN4(A_reg[26]), .IN5(
        n787), .IN6(n667), .Q(N210) );
  AO222X1 U1268 ( .IN1(N103), .IN2(n928), .IN3(n921), .IN4(A_reg[27]), .IN5(
        n925), .IN6(n671), .Q(n538) );
  AO222X1 U1269 ( .IN1(N104), .IN2(n928), .IN3(n921), .IN4(A_reg[28]), .IN5(
        n925), .IN6(n668), .Q(n537) );
  AO222X1 U1270 ( .IN1(N104), .IN2(n944), .IN3(n797), .IN4(A_reg[28]), .IN5(
        n784), .IN6(n668), .Q(N208) );
  AO222X1 U1271 ( .IN1(N105), .IN2(n928), .IN3(n921), .IN4(A_reg[29]), .IN5(
        n925), .IN6(n669), .Q(n536) );
  AO222X1 U1272 ( .IN1(N105), .IN2(n883), .IN3(n797), .IN4(A_reg[29]), .IN5(
        n930), .IN6(n669), .Q(N207) );
  AO222X1 U1273 ( .IN1(N106), .IN2(n928), .IN3(n921), .IN4(A_reg[30]), .IN5(
        n925), .IN6(n673), .Q(n535) );
  AO222X1 U1274 ( .IN1(N106), .IN2(n883), .IN3(n797), .IN4(A_reg[30]), .IN5(
        n786), .IN6(n673), .Q(N206) );
  AO22X1 U1275 ( .IN1(n928), .IN2(N107), .IN3(n925), .IN4(n674), .Q(n534) );
  NAND2X1 U1276 ( .IN1(n909), .IN2(n976), .QN(n1054) );
  XOR2X1 U1277 ( .IN1(n1051), .IN2(A[31]), .Q(n1053) );
  AO222X1 U1278 ( .IN1(N337), .IN2(n958), .IN3(n947), .IN4(N267), .IN5(n952), 
        .IN6(n713), .Q(n503) );
  AO222X1 U1279 ( .IN1(N338), .IN2(n956), .IN3(n947), .IN4(N266), .IN5(n952), 
        .IN6(n714), .Q(n502) );
  AO222X1 U1280 ( .IN1(N339), .IN2(n956), .IN3(n947), .IN4(N265), .IN5(n952), 
        .IN6(n715), .Q(n501) );
  AO222X1 U1281 ( .IN1(N340), .IN2(n956), .IN3(n947), .IN4(N264), .IN5(n952), 
        .IN6(n716), .Q(n500) );
  AO222X1 U1282 ( .IN1(N341), .IN2(n956), .IN3(n947), .IN4(N263), .IN5(n952), 
        .IN6(n717), .Q(n499) );
  AO222X1 U1283 ( .IN1(N342), .IN2(n956), .IN3(n947), .IN4(n601), .IN5(n952), 
        .IN6(n718), .Q(n498) );
  AO222X1 U1284 ( .IN1(N343), .IN2(n956), .IN3(n947), .IN4(N261), .IN5(n952), 
        .IN6(n719), .Q(n497) );
  AO222X1 U1285 ( .IN1(N344), .IN2(n956), .IN3(n947), .IN4(N260), .IN5(n952), 
        .IN6(n720), .Q(n496) );
  AO222X1 U1286 ( .IN1(N345), .IN2(n956), .IN3(n947), .IN4(N259), .IN5(n952), 
        .IN6(n721), .Q(n495) );
  AO222X1 U1287 ( .IN1(N346), .IN2(n956), .IN3(n947), .IN4(N258), .IN5(n952), 
        .IN6(n722), .Q(n494) );
  AO222X1 U1288 ( .IN1(N347), .IN2(n956), .IN3(n947), .IN4(N257), .IN5(n952), 
        .IN6(n723), .Q(n493) );
  AO222X1 U1289 ( .IN1(N348), .IN2(n956), .IN3(n947), .IN4(N256), .IN5(n952), 
        .IN6(n724), .Q(n492) );
  AO222X1 U1290 ( .IN1(N349), .IN2(n956), .IN3(n948), .IN4(N255), .IN5(n953), 
        .IN6(n725), .Q(n491) );
  AO222X1 U1291 ( .IN1(N350), .IN2(n956), .IN3(n948), .IN4(N254), .IN5(n953), 
        .IN6(n726), .Q(n490) );
  AO222X1 U1292 ( .IN1(N351), .IN2(n957), .IN3(n948), .IN4(N253), .IN5(n953), 
        .IN6(n727), .Q(n489) );
  AO222X1 U1293 ( .IN1(N352), .IN2(n957), .IN3(n948), .IN4(N252), .IN5(n953), 
        .IN6(n728), .Q(n488) );
  AO222X1 U1294 ( .IN1(N353), .IN2(n957), .IN3(n948), .IN4(n602), .IN5(n953), 
        .IN6(n729), .Q(n487) );
  AO222X1 U1295 ( .IN1(N354), .IN2(n957), .IN3(n948), .IN4(N250), .IN5(n953), 
        .IN6(n730), .Q(n486) );
  AO222X1 U1296 ( .IN1(N355), .IN2(n957), .IN3(n948), .IN4(N249), .IN5(n953), 
        .IN6(n731), .Q(n485) );
  AO222X1 U1297 ( .IN1(N356), .IN2(n957), .IN3(n948), .IN4(N248), .IN5(n953), 
        .IN6(n732), .Q(n484) );
  AO222X1 U1298 ( .IN1(N357), .IN2(n957), .IN3(n948), .IN4(N247), .IN5(n953), 
        .IN6(n733), .Q(n483) );
  AO222X1 U1299 ( .IN1(N358), .IN2(n957), .IN3(n948), .IN4(N246), .IN5(n953), 
        .IN6(n734), .Q(n482) );
  AO222X1 U1300 ( .IN1(N359), .IN2(n957), .IN3(n948), .IN4(N245), .IN5(n953), 
        .IN6(n735), .Q(n481) );
  AO222X1 U1301 ( .IN1(N360), .IN2(n957), .IN3(n948), .IN4(N244), .IN5(n953), 
        .IN6(n736), .Q(n480) );
  AO222X1 U1302 ( .IN1(N361), .IN2(n957), .IN3(n949), .IN4(N243), .IN5(n1054), 
        .IN6(n737), .Q(n479) );
  AO222X1 U1303 ( .IN1(N362), .IN2(n957), .IN3(n949), .IN4(N242), .IN5(n1054), 
        .IN6(n738), .Q(n478) );
  AO222X1 U1304 ( .IN1(N363), .IN2(n957), .IN3(n949), .IN4(N241), .IN5(n1054), 
        .IN6(n739), .Q(n477) );
  AO222X1 U1305 ( .IN1(N364), .IN2(n957), .IN3(n949), .IN4(N240), .IN5(n1054), 
        .IN6(n740), .Q(n476) );
  AO222X1 U1306 ( .IN1(N365), .IN2(n958), .IN3(n949), .IN4(N239), .IN5(n1054), 
        .IN6(n741), .Q(n475) );
  AO222X1 U1307 ( .IN1(N366), .IN2(n958), .IN3(n949), .IN4(N238), .IN5(n1054), 
        .IN6(n742), .Q(n440) );
  AO222X1 U1308 ( .IN1(N367), .IN2(n958), .IN3(n949), .IN4(N237), .IN5(n1054), 
        .IN6(n743), .Q(n474) );
  AO222X1 U1309 ( .IN1(N368), .IN2(n958), .IN3(N303), .IN4(n949), .IN5(n1054), 
        .IN6(n744), .Q(n473) );
  AO222X1 U1310 ( .IN1(N369), .IN2(n958), .IN3(N304), .IN4(n949), .IN5(n952), 
        .IN6(n745), .Q(n472) );
  AO222X1 U1311 ( .IN1(N370), .IN2(n958), .IN3(N305), .IN4(n949), .IN5(n954), 
        .IN6(n746), .Q(n471) );
  AO222X1 U1312 ( .IN1(N371), .IN2(n958), .IN3(N306), .IN4(n949), .IN5(n954), 
        .IN6(n747), .Q(n470) );
  AO222X1 U1313 ( .IN1(N372), .IN2(n958), .IN3(N307), .IN4(n949), .IN5(n954), 
        .IN6(n748), .Q(n469) );
  AO222X1 U1314 ( .IN1(N373), .IN2(n958), .IN3(N308), .IN4(n949), .IN5(n1054), 
        .IN6(n749), .Q(n468) );
  AO222X1 U1315 ( .IN1(N374), .IN2(n958), .IN3(N309), .IN4(n950), .IN5(n1054), 
        .IN6(n750), .Q(n467) );
  AO222X1 U1316 ( .IN1(N375), .IN2(n958), .IN3(n802), .IN4(n950), .IN5(n1054), 
        .IN6(n751), .Q(n466) );
  AO222X1 U1317 ( .IN1(N376), .IN2(n958), .IN3(N311), .IN4(n950), .IN5(n1054), 
        .IN6(n752), .Q(n465) );
  AO222X1 U1318 ( .IN1(N377), .IN2(n958), .IN3(n807), .IN4(n950), .IN5(n953), 
        .IN6(n753), .Q(n464) );
  AO222X1 U1319 ( .IN1(N378), .IN2(n959), .IN3(N313), .IN4(n950), .IN5(n954), 
        .IN6(n754), .Q(n463) );
  AO222X1 U1320 ( .IN1(N379), .IN2(n959), .IN3(n805), .IN4(n950), .IN5(n954), 
        .IN6(n755), .Q(n462) );
  AO222X1 U1321 ( .IN1(N380), .IN2(n959), .IN3(n871), .IN4(n950), .IN5(n954), 
        .IN6(n756), .Q(n461) );
  AO222X1 U1322 ( .IN1(N381), .IN2(n959), .IN3(n799), .IN4(n950), .IN5(n954), 
        .IN6(n757), .Q(n460) );
  AO222X1 U1323 ( .IN1(N382), .IN2(n959), .IN3(n829), .IN4(n950), .IN5(n954), 
        .IN6(n758), .Q(n459) );
  AO222X1 U1324 ( .IN1(N383), .IN2(n959), .IN3(n881), .IN4(n950), .IN5(n954), 
        .IN6(n759), .Q(n458) );
  AO222X1 U1325 ( .IN1(N385), .IN2(n959), .IN3(N320), .IN4(n950), .IN5(n953), 
        .IN6(n760), .Q(n456) );
  AO222X1 U1326 ( .IN1(N386), .IN2(n959), .IN3(N321), .IN4(n950), .IN5(n952), 
        .IN6(n761), .Q(n455) );
  AO222X1 U1327 ( .IN1(N387), .IN2(n959), .IN3(n870), .IN4(n951), .IN5(n954), 
        .IN6(n762), .Q(n454) );
  AO222X1 U1328 ( .IN1(N388), .IN2(n959), .IN3(n803), .IN4(n951), .IN5(n953), 
        .IN6(n763), .Q(n453) );
  AO222X1 U1329 ( .IN1(N389), .IN2(n959), .IN3(N324), .IN4(n951), .IN5(n952), 
        .IN6(n764), .Q(n452) );
  AO222X1 U1330 ( .IN1(N390), .IN2(n959), .IN3(n794), .IN4(n951), .IN5(n953), 
        .IN6(n765), .Q(n451) );
  AO222X1 U1331 ( .IN1(N391), .IN2(n959), .IN3(N326), .IN4(n951), .IN5(n952), 
        .IN6(n766), .Q(n450) );
  AO222X1 U1332 ( .IN1(n954), .IN2(n768), .IN3(N334), .IN4(n951), .IN5(n956), 
        .IN6(N399), .Q(n442) );
  AO22X1 U1333 ( .IN1(n960), .IN2(N400), .IN3(n954), .IN4(n767), .Q(n441) );
endmodule

