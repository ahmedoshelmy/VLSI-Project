
module WallaceTreeMultiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119;
  wire   [63:1] carry;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  FADDX1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  FADDX1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  FADDX1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  FADDX1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  FADDX1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  FADDX1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  FADDX1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  FADDX1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  FADDX1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  FADDX1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  FADDX1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(n24), .B(n39), .CI(carry[14]), .CO(carry[15]), .S(SUM[14])
         );
  FADDX1 U1_13 ( .A(A[13]), .B(n119), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  XOR3X1 U1_63 ( .IN1(A[63]), .IN2(B[63]), .IN3(carry[63]), .Q(SUM[63]) );
  XOR3X2 U1 ( .IN1(A[24]), .IN2(B[24]), .IN3(carry[24]), .Q(SUM[24]) );
  XOR3X2 U2 ( .IN1(A[30]), .IN2(B[30]), .IN3(carry[30]), .Q(SUM[30]) );
  XOR3X2 U3 ( .IN1(A[48]), .IN2(B[48]), .IN3(carry[48]), .Q(SUM[48]) );
  XOR3X2 U4 ( .IN1(A[51]), .IN2(B[51]), .IN3(carry[51]), .Q(SUM[51]) );
  XOR3X2 U5 ( .IN1(A[61]), .IN2(B[61]), .IN3(carry[61]), .Q(SUM[61]) );
  XOR3X2 U6 ( .IN1(A[36]), .IN2(B[36]), .IN3(carry[36]), .Q(SUM[36]) );
  XOR3X2 U7 ( .IN1(A[54]), .IN2(B[54]), .IN3(carry[54]), .Q(SUM[54]) );
  XOR3X2 U8 ( .IN1(A[40]), .IN2(B[40]), .IN3(carry[40]), .Q(SUM[40]) );
  XOR3X2 U9 ( .IN1(A[58]), .IN2(B[58]), .IN3(carry[58]), .Q(SUM[58]) );
  XOR3X2 U10 ( .IN1(A[26]), .IN2(B[26]), .IN3(carry[26]), .Q(SUM[26]) );
  XOR3X2 U11 ( .IN1(A[42]), .IN2(B[42]), .IN3(carry[42]), .Q(SUM[42]) );
  XOR3X2 U12 ( .IN1(A[18]), .IN2(B[18]), .IN3(carry[18]), .Q(SUM[18]) );
  XOR3X1 U13 ( .IN1(A[10]), .IN2(B[10]), .IN3(carry[10]), .Q(SUM[10]) );
  XOR3X1 U14 ( .IN1(B[16]), .IN2(A[16]), .IN3(carry[16]), .Q(SUM[16]) );
  XOR2X1 U15 ( .IN1(A[53]), .IN2(B[53]), .Q(n58) );
  XOR2X1 U16 ( .IN1(A[57]), .IN2(B[57]), .Q(n47) );
  AND2X1 U17 ( .IN1(B[1]), .IN2(A[1]), .Q(n1) );
  NAND2X1 U18 ( .IN1(A[24]), .IN2(B[24]), .QN(n2) );
  NAND2X0 U19 ( .IN1(A[24]), .IN2(carry[24]), .QN(n3) );
  NAND2X0 U20 ( .IN1(B[24]), .IN2(carry[24]), .QN(n4) );
  NAND3X0 U21 ( .IN1(n2), .IN2(n3), .IN3(n4), .QN(carry[25]) );
  XOR2X1 U22 ( .IN1(A[25]), .IN2(B[25]), .Q(n5) );
  XOR2X1 U23 ( .IN1(n5), .IN2(carry[25]), .Q(SUM[25]) );
  NAND2X1 U24 ( .IN1(A[25]), .IN2(B[25]), .QN(n6) );
  NAND2X0 U25 ( .IN1(A[25]), .IN2(carry[25]), .QN(n7) );
  NAND2X0 U26 ( .IN1(B[25]), .IN2(carry[25]), .QN(n8) );
  NAND3X0 U27 ( .IN1(n6), .IN2(n7), .IN3(n8), .QN(carry[26]) );
  NAND2X1 U28 ( .IN1(B[16]), .IN2(A[16]), .QN(n9) );
  NAND2X0 U29 ( .IN1(B[16]), .IN2(carry[16]), .QN(n10) );
  NAND2X0 U30 ( .IN1(A[16]), .IN2(carry[16]), .QN(n11) );
  NAND3X0 U31 ( .IN1(n9), .IN2(n10), .IN3(n11), .QN(carry[17]) );
  XOR2X1 U32 ( .IN1(B[17]), .IN2(A[17]), .Q(n12) );
  XOR2X1 U33 ( .IN1(n12), .IN2(carry[17]), .Q(SUM[17]) );
  NAND2X1 U34 ( .IN1(B[17]), .IN2(A[17]), .QN(n13) );
  NAND2X0 U35 ( .IN1(B[17]), .IN2(carry[17]), .QN(n14) );
  NAND2X0 U36 ( .IN1(A[17]), .IN2(carry[17]), .QN(n15) );
  NAND3X0 U37 ( .IN1(n13), .IN2(n14), .IN3(n15), .QN(carry[18]) );
  NAND2X1 U38 ( .IN1(A[42]), .IN2(B[42]), .QN(n16) );
  NAND2X0 U39 ( .IN1(A[42]), .IN2(carry[42]), .QN(n17) );
  NAND2X0 U40 ( .IN1(B[42]), .IN2(carry[42]), .QN(n18) );
  NAND3X0 U41 ( .IN1(n16), .IN2(n17), .IN3(n18), .QN(carry[43]) );
  XOR2X1 U42 ( .IN1(A[43]), .IN2(B[43]), .Q(n19) );
  XOR2X1 U43 ( .IN1(n19), .IN2(carry[43]), .Q(SUM[43]) );
  NAND2X1 U44 ( .IN1(A[43]), .IN2(B[43]), .QN(n20) );
  NAND2X0 U45 ( .IN1(A[43]), .IN2(carry[43]), .QN(n21) );
  NAND2X0 U46 ( .IN1(B[43]), .IN2(carry[43]), .QN(n22) );
  NAND3X0 U47 ( .IN1(n20), .IN2(n21), .IN3(n22), .QN(carry[44]) );
  INVX0 U48 ( .INP(A[14]), .ZN(n23) );
  INVX0 U49 ( .INP(n23), .ZN(n24) );
  XOR3X1 U50 ( .IN1(carry[35]), .IN2(A[35]), .IN3(B[35]), .Q(SUM[35]) );
  NAND2X0 U51 ( .IN1(carry[35]), .IN2(B[35]), .QN(n25) );
  NAND2X0 U52 ( .IN1(carry[35]), .IN2(A[35]), .QN(n26) );
  NAND2X0 U53 ( .IN1(B[35]), .IN2(A[35]), .QN(n27) );
  NAND3X0 U54 ( .IN1(n25), .IN2(n26), .IN3(n27), .QN(carry[36]) );
  XOR3X1 U55 ( .IN1(carry[39]), .IN2(A[39]), .IN3(B[39]), .Q(SUM[39]) );
  NAND2X0 U56 ( .IN1(carry[39]), .IN2(B[39]), .QN(n28) );
  NAND2X0 U57 ( .IN1(carry[39]), .IN2(A[39]), .QN(n29) );
  NAND2X0 U58 ( .IN1(B[39]), .IN2(A[39]), .QN(n30) );
  NAND3X0 U59 ( .IN1(n28), .IN2(n30), .IN3(n29), .QN(carry[40]) );
  NAND2X1 U60 ( .IN1(A[40]), .IN2(B[40]), .QN(n31) );
  NAND2X0 U61 ( .IN1(A[40]), .IN2(carry[40]), .QN(n32) );
  NAND2X0 U62 ( .IN1(B[40]), .IN2(carry[40]), .QN(n33) );
  NAND3X0 U63 ( .IN1(n31), .IN2(n32), .IN3(n33), .QN(carry[41]) );
  XOR2X1 U64 ( .IN1(A[41]), .IN2(B[41]), .Q(n34) );
  XOR2X1 U65 ( .IN1(n34), .IN2(carry[41]), .Q(SUM[41]) );
  NAND2X1 U66 ( .IN1(A[41]), .IN2(B[41]), .QN(n35) );
  NAND2X0 U67 ( .IN1(A[41]), .IN2(carry[41]), .QN(n36) );
  NAND2X0 U68 ( .IN1(B[41]), .IN2(carry[41]), .QN(n37) );
  NAND3X0 U69 ( .IN1(n35), .IN2(n36), .IN3(n37), .QN(carry[42]) );
  INVX0 U70 ( .INP(B[14]), .ZN(n38) );
  INVX0 U71 ( .INP(n38), .ZN(n39) );
  NAND2X1 U72 ( .IN1(A[10]), .IN2(B[10]), .QN(n40) );
  NAND2X0 U73 ( .IN1(A[10]), .IN2(carry[10]), .QN(n41) );
  NAND2X0 U74 ( .IN1(B[10]), .IN2(carry[10]), .QN(n42) );
  NAND3X0 U75 ( .IN1(n41), .IN2(n40), .IN3(n42), .QN(carry[11]) );
  XOR2X1 U76 ( .IN1(B[11]), .IN2(A[11]), .Q(n43) );
  XOR2X1 U77 ( .IN1(n43), .IN2(carry[11]), .Q(SUM[11]) );
  NAND2X1 U78 ( .IN1(B[11]), .IN2(A[11]), .QN(n44) );
  NAND2X0 U79 ( .IN1(B[11]), .IN2(carry[11]), .QN(n45) );
  NAND2X0 U80 ( .IN1(A[11]), .IN2(carry[11]), .QN(n46) );
  NAND3X0 U81 ( .IN1(n44), .IN2(n45), .IN3(n46), .QN(carry[12]) );
  XOR2X1 U82 ( .IN1(n47), .IN2(carry[57]), .Q(SUM[57]) );
  NAND2X0 U83 ( .IN1(carry[57]), .IN2(B[57]), .QN(n48) );
  NAND2X0 U84 ( .IN1(carry[57]), .IN2(A[57]), .QN(n49) );
  NAND2X0 U85 ( .IN1(B[57]), .IN2(A[57]), .QN(n50) );
  NAND3X0 U86 ( .IN1(n48), .IN2(n50), .IN3(n49), .QN(carry[58]) );
  NAND2X1 U87 ( .IN1(A[30]), .IN2(B[30]), .QN(n51) );
  NAND2X0 U88 ( .IN1(A[30]), .IN2(carry[30]), .QN(n52) );
  NAND2X0 U89 ( .IN1(B[30]), .IN2(carry[30]), .QN(n53) );
  NAND3X0 U90 ( .IN1(n51), .IN2(n52), .IN3(n53), .QN(carry[31]) );
  XOR2X1 U91 ( .IN1(A[31]), .IN2(B[31]), .Q(n54) );
  XOR2X1 U92 ( .IN1(n54), .IN2(carry[31]), .Q(SUM[31]) );
  NAND2X1 U93 ( .IN1(A[31]), .IN2(B[31]), .QN(n55) );
  NAND2X0 U94 ( .IN1(A[31]), .IN2(carry[31]), .QN(n56) );
  NAND2X0 U95 ( .IN1(B[31]), .IN2(carry[31]), .QN(n57) );
  NAND3X0 U96 ( .IN1(n55), .IN2(n56), .IN3(n57), .QN(carry[32]) );
  XOR2X1 U97 ( .IN1(n58), .IN2(carry[53]), .Q(SUM[53]) );
  NAND2X0 U98 ( .IN1(carry[53]), .IN2(B[53]), .QN(n59) );
  NAND2X0 U99 ( .IN1(carry[53]), .IN2(A[53]), .QN(n60) );
  NAND2X0 U100 ( .IN1(B[53]), .IN2(A[53]), .QN(n61) );
  NAND3X0 U101 ( .IN1(n59), .IN2(n60), .IN3(n61), .QN(carry[54]) );
  NAND2X1 U102 ( .IN1(A[48]), .IN2(B[48]), .QN(n62) );
  NAND2X0 U103 ( .IN1(A[48]), .IN2(carry[48]), .QN(n63) );
  NAND2X0 U104 ( .IN1(B[48]), .IN2(carry[48]), .QN(n64) );
  NAND3X0 U105 ( .IN1(n63), .IN2(n62), .IN3(n64), .QN(carry[49]) );
  XOR2X1 U106 ( .IN1(A[49]), .IN2(B[49]), .Q(n65) );
  XOR2X1 U107 ( .IN1(n65), .IN2(carry[49]), .Q(SUM[49]) );
  NAND2X1 U108 ( .IN1(A[49]), .IN2(B[49]), .QN(n66) );
  NAND2X0 U109 ( .IN1(A[49]), .IN2(carry[49]), .QN(n67) );
  NAND2X0 U110 ( .IN1(B[49]), .IN2(carry[49]), .QN(n68) );
  NAND3X0 U111 ( .IN1(n66), .IN2(n67), .IN3(n68), .QN(carry[50]) );
  NAND2X1 U112 ( .IN1(A[26]), .IN2(B[26]), .QN(n69) );
  NAND2X0 U113 ( .IN1(A[26]), .IN2(carry[26]), .QN(n70) );
  NAND2X0 U114 ( .IN1(B[26]), .IN2(carry[26]), .QN(n71) );
  NAND3X0 U115 ( .IN1(n70), .IN2(n69), .IN3(n71), .QN(carry[27]) );
  XOR2X1 U116 ( .IN1(A[27]), .IN2(B[27]), .Q(n72) );
  XOR2X1 U117 ( .IN1(n72), .IN2(carry[27]), .Q(SUM[27]) );
  NAND2X1 U118 ( .IN1(A[27]), .IN2(B[27]), .QN(n73) );
  NAND2X0 U119 ( .IN1(A[27]), .IN2(carry[27]), .QN(n74) );
  NAND2X0 U120 ( .IN1(B[27]), .IN2(carry[27]), .QN(n75) );
  NAND3X0 U121 ( .IN1(n73), .IN2(n74), .IN3(n75), .QN(carry[28]) );
  NAND2X1 U122 ( .IN1(A[51]), .IN2(B[51]), .QN(n76) );
  NAND2X0 U123 ( .IN1(A[51]), .IN2(carry[51]), .QN(n77) );
  NAND2X0 U124 ( .IN1(B[51]), .IN2(carry[51]), .QN(n78) );
  NAND3X0 U125 ( .IN1(n76), .IN2(n77), .IN3(n78), .QN(carry[52]) );
  XOR2X1 U126 ( .IN1(A[52]), .IN2(B[52]), .Q(n79) );
  XOR2X1 U127 ( .IN1(n79), .IN2(carry[52]), .Q(SUM[52]) );
  NAND2X1 U128 ( .IN1(A[52]), .IN2(B[52]), .QN(n80) );
  NAND2X0 U129 ( .IN1(A[52]), .IN2(carry[52]), .QN(n81) );
  NAND2X0 U130 ( .IN1(B[52]), .IN2(carry[52]), .QN(n82) );
  NAND3X0 U131 ( .IN1(n80), .IN2(n81), .IN3(n82), .QN(carry[53]) );
  NAND2X1 U132 ( .IN1(A[36]), .IN2(B[36]), .QN(n83) );
  NAND2X0 U133 ( .IN1(A[36]), .IN2(carry[36]), .QN(n84) );
  NAND2X0 U134 ( .IN1(B[36]), .IN2(carry[36]), .QN(n85) );
  NAND3X0 U135 ( .IN1(n83), .IN2(n84), .IN3(n85), .QN(carry[37]) );
  XOR2X1 U136 ( .IN1(A[37]), .IN2(B[37]), .Q(n86) );
  XOR2X1 U137 ( .IN1(n86), .IN2(carry[37]), .Q(SUM[37]) );
  NAND2X1 U138 ( .IN1(A[37]), .IN2(B[37]), .QN(n87) );
  NAND2X0 U139 ( .IN1(A[37]), .IN2(carry[37]), .QN(n88) );
  NAND2X0 U140 ( .IN1(B[37]), .IN2(carry[37]), .QN(n89) );
  NAND3X0 U141 ( .IN1(n87), .IN2(n88), .IN3(n89), .QN(carry[38]) );
  NAND2X1 U142 ( .IN1(A[18]), .IN2(B[18]), .QN(n90) );
  NAND2X0 U143 ( .IN1(A[18]), .IN2(carry[18]), .QN(n91) );
  NAND2X0 U144 ( .IN1(B[18]), .IN2(carry[18]), .QN(n92) );
  NAND3X0 U145 ( .IN1(n90), .IN2(n91), .IN3(n92), .QN(carry[19]) );
  XOR2X1 U146 ( .IN1(A[19]), .IN2(B[19]), .Q(n93) );
  XOR2X1 U147 ( .IN1(n93), .IN2(carry[19]), .Q(SUM[19]) );
  NAND2X1 U148 ( .IN1(A[19]), .IN2(B[19]), .QN(n94) );
  NAND2X0 U149 ( .IN1(A[19]), .IN2(carry[19]), .QN(n95) );
  NAND2X0 U150 ( .IN1(B[19]), .IN2(carry[19]), .QN(n96) );
  NAND3X0 U151 ( .IN1(n94), .IN2(n95), .IN3(n96), .QN(carry[20]) );
  NAND2X1 U152 ( .IN1(A[54]), .IN2(B[54]), .QN(n97) );
  NAND2X0 U153 ( .IN1(A[54]), .IN2(carry[54]), .QN(n98) );
  NAND2X0 U154 ( .IN1(B[54]), .IN2(carry[54]), .QN(n99) );
  NAND3X0 U155 ( .IN1(n97), .IN2(n98), .IN3(n99), .QN(carry[55]) );
  XOR2X1 U156 ( .IN1(A[55]), .IN2(B[55]), .Q(n100) );
  XOR2X1 U157 ( .IN1(n100), .IN2(carry[55]), .Q(SUM[55]) );
  NAND2X1 U158 ( .IN1(A[55]), .IN2(B[55]), .QN(n101) );
  NAND2X0 U159 ( .IN1(A[55]), .IN2(carry[55]), .QN(n102) );
  NAND2X0 U160 ( .IN1(B[55]), .IN2(carry[55]), .QN(n103) );
  NAND3X0 U161 ( .IN1(n101), .IN2(n102), .IN3(n103), .QN(carry[56]) );
  NAND2X1 U162 ( .IN1(A[58]), .IN2(B[58]), .QN(n104) );
  NAND2X0 U163 ( .IN1(A[58]), .IN2(carry[58]), .QN(n105) );
  NAND2X0 U164 ( .IN1(B[58]), .IN2(carry[58]), .QN(n106) );
  NAND3X0 U165 ( .IN1(n104), .IN2(n105), .IN3(n106), .QN(carry[59]) );
  XOR2X1 U166 ( .IN1(A[59]), .IN2(B[59]), .Q(n107) );
  XOR2X1 U167 ( .IN1(n107), .IN2(carry[59]), .Q(SUM[59]) );
  NAND2X1 U168 ( .IN1(A[59]), .IN2(B[59]), .QN(n108) );
  NAND2X0 U169 ( .IN1(A[59]), .IN2(carry[59]), .QN(n109) );
  NAND2X0 U170 ( .IN1(B[59]), .IN2(carry[59]), .QN(n110) );
  NAND3X0 U171 ( .IN1(n108), .IN2(n109), .IN3(n110), .QN(carry[60]) );
  NAND2X1 U172 ( .IN1(A[61]), .IN2(B[61]), .QN(n111) );
  NAND2X0 U173 ( .IN1(A[61]), .IN2(carry[61]), .QN(n112) );
  NAND2X0 U174 ( .IN1(B[61]), .IN2(carry[61]), .QN(n113) );
  NAND3X0 U175 ( .IN1(n112), .IN2(n111), .IN3(n113), .QN(carry[62]) );
  XOR2X1 U176 ( .IN1(A[62]), .IN2(B[62]), .Q(n114) );
  XOR2X1 U177 ( .IN1(n114), .IN2(carry[62]), .Q(SUM[62]) );
  NAND2X1 U178 ( .IN1(A[62]), .IN2(B[62]), .QN(n115) );
  NAND2X0 U179 ( .IN1(A[62]), .IN2(carry[62]), .QN(n116) );
  NAND2X0 U180 ( .IN1(B[62]), .IN2(carry[62]), .QN(n117) );
  NAND3X0 U181 ( .IN1(n115), .IN2(n116), .IN3(n117), .QN(carry[63]) );
  XOR2X1 U182 ( .IN1(B[1]), .IN2(A[1]), .Q(SUM[1]) );
  INVX0 U183 ( .INP(B[13]), .ZN(n118) );
  INVX0 U184 ( .INP(n118), .ZN(n119) );
endmodule


module WallaceTreeMultiplier ( A, B, out, clk, rst );
  input [31:0] A;
  input [31:0] B;
  output [63:0] out;
  input clk, rst;
  wire   N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, \p[7][63] , \p[7][37] ,
         \p[7][36] , \p[7][35] , \p[7][34] , \p[7][33] , \p[7][32] ,
         \p[7][31] , \p[7][30] , \p[7][29] , \p[7][28] , \p[7][27] ,
         \p[7][26] , \p[7][25] , \p[7][24] , \p[7][23] , \p[7][22] ,
         \p[7][21] , \p[7][20] , \p[7][19] , \p[7][18] , \p[7][17] ,
         \p[7][16] , \p[7][15] , \p[7][14] , \p[7][13] , \p[7][12] ,
         \p[7][11] , \p[7][10] , \p[7][9] , \p[7][8] , \p[7][7] , \p[6][63] ,
         \p[6][36] , \p[6][35] , \p[6][34] , \p[6][33] , \p[6][32] ,
         \p[6][31] , \p[6][30] , \p[6][29] , \p[6][28] , \p[6][27] ,
         \p[6][26] , \p[6][25] , \p[6][24] , \p[6][23] , \p[6][22] ,
         \p[6][21] , \p[6][20] , \p[6][19] , \p[6][18] , \p[6][17] ,
         \p[6][16] , \p[6][15] , \p[6][14] , \p[6][13] , \p[6][12] ,
         \p[6][11] , \p[6][10] , \p[6][9] , \p[6][8] , \p[6][7] , \p[6][6] ,
         \p[5][63] , \p[5][35] , \p[5][34] , \p[5][33] , \p[5][32] ,
         \p[5][31] , \p[5][30] , \p[5][29] , \p[5][28] , \p[5][27] ,
         \p[5][26] , \p[5][25] , \p[5][24] , \p[5][23] , \p[5][22] ,
         \p[5][21] , \p[5][20] , \p[5][19] , \p[5][18] , \p[5][17] ,
         \p[5][16] , \p[5][15] , \p[5][14] , \p[5][13] , \p[5][12] ,
         \p[5][11] , \p[5][10] , \p[5][9] , \p[5][8] , \p[5][7] , \p[5][6] ,
         \p[5][5] , \p[4][63] , \p[4][34] , \p[4][33] , \p[4][32] , \p[4][31] ,
         \p[4][30] , \p[4][29] , \p[4][28] , \p[4][27] , \p[4][26] ,
         \p[4][25] , \p[4][24] , \p[4][23] , \p[4][22] , \p[4][21] ,
         \p[4][20] , \p[4][19] , \p[4][18] , \p[4][17] , \p[4][16] ,
         \p[4][15] , \p[4][14] , \p[4][13] , \p[4][12] , \p[4][11] ,
         \p[4][10] , \p[4][9] , \p[4][8] , \p[4][7] , \p[4][6] , \p[4][5] ,
         \p[4][4] , \p[3][63] , \p[3][33] , \p[3][32] , \p[3][31] , \p[3][30] ,
         \p[3][29] , \p[3][28] , \p[3][27] , \p[3][26] , \p[3][25] ,
         \p[3][24] , \p[3][23] , \p[3][22] , \p[3][21] , \p[3][20] ,
         \p[3][19] , \p[3][18] , \p[3][17] , \p[3][16] , \p[3][15] ,
         \p[3][14] , \p[3][13] , \p[3][12] , \p[3][11] , \p[3][10] , \p[3][9] ,
         \p[3][8] , \p[3][7] , \p[3][6] , \p[3][5] , \p[3][4] , \p[3][3] ,
         \p[2][63] , \p[2][32] , \p[2][31] , \p[2][30] , \p[2][29] ,
         \p[2][28] , \p[2][27] , \p[2][26] , \p[2][25] , \p[2][24] ,
         \p[2][23] , \p[2][22] , \p[2][21] , \p[2][20] , \p[2][19] ,
         \p[2][18] , \p[2][17] , \p[2][16] , \p[2][15] , \p[2][14] ,
         \p[2][13] , \p[2][12] , \p[2][11] , \p[2][10] , \p[2][9] , \p[2][8] ,
         \p[2][7] , \p[2][6] , \p[2][5] , \p[2][4] , \p[2][3] , \p[2][2] ,
         \p[1][63] , \p[1][31] , \p[1][30] , \p[1][29] , \p[1][28] ,
         \p[1][27] , \p[1][26] , \p[1][25] , \p[1][24] , \p[1][23] ,
         \p[1][22] , \p[1][21] , \p[1][20] , \p[1][19] , \p[1][18] ,
         \p[1][17] , \p[1][16] , \p[1][15] , \p[1][14] , \p[1][13] ,
         \p[1][12] , \p[1][11] , \p[1][10] , \p[1][9] , \p[1][8] , \p[1][7] ,
         \p[1][6] , \p[1][5] , \p[1][4] , \p[1][3] , \p[1][2] , \p[1][1] ,
         \p[0][63] , \p[0][30] , \p[0][29] , \p[0][28] , \p[0][27] ,
         \p[0][26] , \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] ,
         \p[0][21] , \p[0][20] , \p[0][19] , \p[0][18] , \p[0][17] ,
         \p[0][16] , \p[0][15] , \p[0][14] , \p[0][13] , \p[0][12] ,
         \p[0][11] , \p[0][10] , \p[0][9] , \p[0][8] , \p[0][7] , \p[0][6] ,
         \p[0][5] , \p[0][4] , \p[0][3] , \p[0][2] , \p[0][1] , \p[0][0] ,
         \p[63][63] , \p[62][63] , \p[61][63] , \p[60][63] , \p[59][63] ,
         \p[58][63] , \p[57][63] , \p[56][63] , \p[55][63] , \p[54][63] ,
         \p[53][63] , \p[52][63] , \p[51][63] , \p[50][63] , \p[49][63] ,
         \p[48][63] , \p[47][63] , \p[46][63] , \p[45][63] , \p[44][63] ,
         \p[43][63] , \p[42][63] , \p[41][63] , \p[40][63] , \p[39][63] ,
         \p[38][63] , \p[37][63] , \p[36][63] , \p[35][63] , \p[34][63] ,
         \p[33][63] , \p[32][63] , \p[30][63] , \p[30][60] , \p[30][59] ,
         \p[30][58] , \p[30][57] , \p[30][56] , \p[30][55] , \p[30][54] ,
         \p[30][53] , \p[30][52] , \p[30][51] , \p[30][50] , \p[30][49] ,
         \p[30][48] , \p[30][47] , \p[30][46] , \p[30][45] , \p[30][44] ,
         \p[30][43] , \p[30][42] , \p[30][41] , \p[30][40] , \p[30][39] ,
         \p[30][38] , \p[30][37] , \p[30][36] , \p[30][35] , \p[30][34] ,
         \p[30][33] , \p[30][32] , \p[30][31] , \p[30][30] , \p[29][63] ,
         \p[29][59] , \p[29][58] , \p[29][57] , \p[29][56] , \p[29][55] ,
         \p[29][54] , \p[29][53] , \p[29][52] , \p[29][51] , \p[29][50] ,
         \p[29][49] , \p[29][48] , \p[29][47] , \p[29][46] , \p[29][45] ,
         \p[29][44] , \p[29][43] , \p[29][42] , \p[29][41] , \p[29][40] ,
         \p[29][39] , \p[29][38] , \p[29][37] , \p[29][36] , \p[29][35] ,
         \p[29][34] , \p[29][33] , \p[29][32] , \p[29][31] , \p[29][30] ,
         \p[29][29] , \p[28][63] , \p[28][58] , \p[28][57] , \p[28][56] ,
         \p[28][55] , \p[28][54] , \p[28][53] , \p[28][52] , \p[28][51] ,
         \p[28][50] , \p[28][49] , \p[28][48] , \p[28][47] , \p[28][46] ,
         \p[28][45] , \p[28][44] , \p[28][43] , \p[28][42] , \p[28][41] ,
         \p[28][40] , \p[28][39] , \p[28][38] , \p[28][37] , \p[28][36] ,
         \p[28][35] , \p[28][34] , \p[28][33] , \p[28][32] , \p[28][31] ,
         \p[28][30] , \p[28][29] , \p[28][28] , \p[27][63] , \p[27][57] ,
         \p[27][56] , \p[27][55] , \p[27][54] , \p[27][53] , \p[27][52] ,
         \p[27][51] , \p[27][50] , \p[27][49] , \p[27][48] , \p[27][47] ,
         \p[27][46] , \p[27][45] , \p[27][44] , \p[27][43] , \p[27][42] ,
         \p[27][41] , \p[27][40] , \p[27][39] , \p[27][38] , \p[27][37] ,
         \p[27][36] , \p[27][35] , \p[27][34] , \p[27][33] , \p[27][32] ,
         \p[27][31] , \p[27][30] , \p[27][29] , \p[27][28] , \p[27][27] ,
         \p[26][63] , \p[26][56] , \p[26][55] , \p[26][54] , \p[26][53] ,
         \p[26][52] , \p[26][51] , \p[26][50] , \p[26][49] , \p[26][48] ,
         \p[26][47] , \p[26][46] , \p[26][45] , \p[26][44] , \p[26][43] ,
         \p[26][42] , \p[26][41] , \p[26][40] , \p[26][39] , \p[26][38] ,
         \p[26][37] , \p[26][36] , \p[26][35] , \p[26][34] , \p[26][33] ,
         \p[26][32] , \p[26][31] , \p[26][30] , \p[26][29] , \p[26][28] ,
         \p[26][27] , \p[26][26] , \p[25][63] , \p[25][55] , \p[25][54] ,
         \p[25][53] , \p[25][52] , \p[25][51] , \p[25][50] , \p[25][49] ,
         \p[25][48] , \p[25][47] , \p[25][46] , \p[25][45] , \p[25][44] ,
         \p[25][43] , \p[25][42] , \p[25][41] , \p[25][40] , \p[25][39] ,
         \p[25][38] , \p[25][37] , \p[25][36] , \p[25][35] , \p[25][34] ,
         \p[25][33] , \p[25][32] , \p[25][31] , \p[25][30] , \p[25][29] ,
         \p[25][28] , \p[25][27] , \p[25][26] , \p[25][25] , \p[24][63] ,
         \p[24][54] , \p[24][53] , \p[24][52] , \p[24][51] , \p[24][50] ,
         \p[24][49] , \p[24][48] , \p[24][47] , \p[24][46] , \p[24][45] ,
         \p[24][44] , \p[24][43] , \p[24][42] , \p[24][41] , \p[24][40] ,
         \p[24][39] , \p[24][38] , \p[24][37] , \p[24][36] , \p[24][35] ,
         \p[24][34] , \p[24][33] , \p[24][32] , \p[24][31] , \p[24][30] ,
         \p[24][29] , \p[24][28] , \p[24][27] , \p[24][26] , \p[24][25] ,
         \p[24][24] , \p[23][63] , \p[23][53] , \p[23][52] , \p[23][51] ,
         \p[23][50] , \p[23][49] , \p[23][48] , \p[23][47] , \p[23][46] ,
         \p[23][45] , \p[23][44] , \p[23][43] , \p[23][42] , \p[23][41] ,
         \p[23][40] , \p[23][39] , \p[23][38] , \p[23][37] , \p[23][36] ,
         \p[23][35] , \p[23][34] , \p[23][33] , \p[23][32] , \p[23][31] ,
         \p[23][30] , \p[23][29] , \p[23][28] , \p[23][27] , \p[23][26] ,
         \p[23][25] , \p[23][24] , \p[23][23] , \p[22][63] , \p[22][52] ,
         \p[22][51] , \p[22][50] , \p[22][49] , \p[22][48] , \p[22][47] ,
         \p[22][46] , \p[22][45] , \p[22][44] , \p[22][43] , \p[22][42] ,
         \p[22][41] , \p[22][40] , \p[22][39] , \p[22][38] , \p[22][37] ,
         \p[22][36] , \p[22][35] , \p[22][34] , \p[22][33] , \p[22][32] ,
         \p[22][31] , \p[22][30] , \p[22][29] , \p[22][28] , \p[22][27] ,
         \p[22][26] , \p[22][25] , \p[22][24] , \p[22][23] , \p[22][22] ,
         \p[21][63] , \p[21][51] , \p[21][50] , \p[21][49] , \p[21][48] ,
         \p[21][47] , \p[21][46] , \p[21][45] , \p[21][44] , \p[21][43] ,
         \p[21][42] , \p[21][41] , \p[21][40] , \p[21][39] , \p[21][38] ,
         \p[21][37] , \p[21][36] , \p[21][35] , \p[21][34] , \p[21][33] ,
         \p[21][32] , \p[21][31] , \p[21][30] , \p[21][29] , \p[21][28] ,
         \p[21][27] , \p[21][26] , \p[21][25] , \p[21][24] , \p[21][23] ,
         \p[21][22] , \p[21][21] , \p[20][63] , \p[20][50] , \p[20][49] ,
         \p[20][48] , \p[20][47] , \p[20][46] , \p[20][45] , \p[20][44] ,
         \p[20][43] , \p[20][42] , \p[20][41] , \p[20][40] , \p[20][39] ,
         \p[20][38] , \p[20][37] , \p[20][36] , \p[20][35] , \p[20][34] ,
         \p[20][33] , \p[20][32] , \p[20][31] , \p[20][30] , \p[20][29] ,
         \p[20][28] , \p[20][27] , \p[20][26] , \p[20][25] , \p[20][24] ,
         \p[20][23] , \p[20][22] , \p[20][21] , \p[20][20] , \p[19][63] ,
         \p[19][49] , \p[19][48] , \p[19][47] , \p[19][46] , \p[19][45] ,
         \p[19][44] , \p[19][43] , \p[19][42] , \p[19][41] , \p[19][40] ,
         \p[19][39] , \p[19][38] , \p[19][37] , \p[19][36] , \p[19][35] ,
         \p[19][34] , \p[19][33] , \p[19][32] , \p[19][31] , \p[19][30] ,
         \p[19][29] , \p[19][28] , \p[19][27] , \p[19][26] , \p[19][25] ,
         \p[19][24] , \p[19][23] , \p[19][22] , \p[19][21] , \p[19][20] ,
         \p[19][19] , \p[18][63] , \p[18][48] , \p[18][47] , \p[18][46] ,
         \p[18][45] , \p[18][44] , \p[18][43] , \p[18][42] , \p[18][41] ,
         \p[18][40] , \p[18][39] , \p[18][38] , \p[18][37] , \p[18][36] ,
         \p[18][35] , \p[18][34] , \p[18][33] , \p[18][32] , \p[18][31] ,
         \p[18][30] , \p[18][29] , \p[18][28] , \p[18][27] , \p[18][26] ,
         \p[18][25] , \p[18][24] , \p[18][23] , \p[18][22] , \p[18][21] ,
         \p[18][20] , \p[18][19] , \p[18][18] , \p[17][63] , \p[17][47] ,
         \p[17][46] , \p[17][45] , \p[17][44] , \p[17][43] , \p[17][42] ,
         \p[17][41] , \p[17][40] , \p[17][39] , \p[17][38] , \p[17][37] ,
         \p[17][36] , \p[17][35] , \p[17][34] , \p[17][33] , \p[17][32] ,
         \p[17][31] , \p[17][30] , \p[17][29] , \p[17][28] , \p[17][27] ,
         \p[17][26] , \p[17][25] , \p[17][24] , \p[17][23] , \p[17][22] ,
         \p[17][21] , \p[17][20] , \p[17][19] , \p[17][18] , \p[17][17] ,
         \p[16][63] , \p[16][46] , \p[16][45] , \p[16][44] , \p[16][43] ,
         \p[16][42] , \p[16][41] , \p[16][40] , \p[16][39] , \p[16][38] ,
         \p[16][37] , \p[16][36] , \p[16][35] , \p[16][34] , \p[16][33] ,
         \p[16][32] , \p[16][31] , \p[16][30] , \p[16][29] , \p[16][28] ,
         \p[16][27] , \p[16][26] , \p[16][25] , \p[16][24] , \p[16][23] ,
         \p[16][22] , \p[16][21] , \p[16][20] , \p[16][19] , \p[16][18] ,
         \p[16][17] , \p[16][16] , \p[15][63] , \p[15][45] , \p[15][44] ,
         \p[15][43] , \p[15][42] , \p[15][41] , \p[15][40] , \p[15][39] ,
         \p[15][38] , \p[15][37] , \p[15][36] , \p[15][35] , \p[15][34] ,
         \p[15][33] , \p[15][32] , \p[15][31] , \p[15][30] , \p[15][29] ,
         \p[15][28] , \p[15][27] , \p[15][26] , \p[15][25] , \p[15][24] ,
         \p[15][23] , \p[15][22] , \p[15][21] , \p[15][20] , \p[15][19] ,
         \p[15][18] , \p[15][17] , \p[15][16] , \p[15][15] , \p[14][63] ,
         \p[14][44] , \p[14][43] , \p[14][42] , \p[14][41] , \p[14][40] ,
         \p[14][39] , \p[14][38] , \p[14][37] , \p[14][36] , \p[14][35] ,
         \p[14][34] , \p[14][33] , \p[14][32] , \p[14][31] , \p[14][30] ,
         \p[14][29] , \p[14][28] , \p[14][27] , \p[14][26] , \p[14][25] ,
         \p[14][24] , \p[14][23] , \p[14][22] , \p[14][21] , \p[14][20] ,
         \p[14][19] , \p[14][18] , \p[14][17] , \p[14][16] , \p[14][15] ,
         \p[14][14] , \p[13][63] , \p[13][43] , \p[13][42] , \p[13][41] ,
         \p[13][40] , \p[13][39] , \p[13][38] , \p[13][37] , \p[13][36] ,
         \p[13][35] , \p[13][34] , \p[13][33] , \p[13][32] , \p[13][31] ,
         \p[13][30] , \p[13][29] , \p[13][28] , \p[13][27] , \p[13][26] ,
         \p[13][25] , \p[13][24] , \p[13][23] , \p[13][22] , \p[13][21] ,
         \p[13][20] , \p[13][19] , \p[13][18] , \p[13][17] , \p[13][16] ,
         \p[13][15] , \p[13][14] , \p[13][13] , \p[12][63] , \p[12][42] ,
         \p[12][41] , \p[12][40] , \p[12][39] , \p[12][38] , \p[12][37] ,
         \p[12][36] , \p[12][35] , \p[12][34] , \p[12][33] , \p[12][32] ,
         \p[12][31] , \p[12][30] , \p[12][29] , \p[12][28] , \p[12][27] ,
         \p[12][26] , \p[12][25] , \p[12][24] , \p[12][23] , \p[12][22] ,
         \p[12][21] , \p[12][20] , \p[12][19] , \p[12][18] , \p[12][17] ,
         \p[12][16] , \p[12][15] , \p[12][14] , \p[12][13] , \p[12][12] ,
         \p[11][63] , \p[11][41] , \p[11][40] , \p[11][39] , \p[11][38] ,
         \p[11][37] , \p[11][36] , \p[11][35] , \p[11][34] , \p[11][33] ,
         \p[11][32] , \p[11][31] , \p[11][30] , \p[11][29] , \p[11][28] ,
         \p[11][27] , \p[11][26] , \p[11][25] , \p[11][24] , \p[11][23] ,
         \p[11][22] , \p[11][21] , \p[11][20] , \p[11][19] , \p[11][18] ,
         \p[11][17] , \p[11][16] , \p[11][15] , \p[11][14] , \p[11][13] ,
         \p[11][12] , \p[11][11] , \p[10][63] , \p[10][40] , \p[10][39] ,
         \p[10][38] , \p[10][37] , \p[10][36] , \p[10][35] , \p[10][34] ,
         \p[10][33] , \p[10][32] , \p[10][31] , \p[10][30] , \p[10][29] ,
         \p[10][28] , \p[10][27] , \p[10][26] , \p[10][25] , \p[10][24] ,
         \p[10][23] , \p[10][22] , \p[10][21] , \p[10][20] , \p[10][19] ,
         \p[10][18] , \p[10][17] , \p[10][16] , \p[10][15] , \p[10][14] ,
         \p[10][13] , \p[10][12] , \p[10][11] , \p[10][10] , \p[9][63] ,
         \p[9][39] , \p[9][38] , \p[9][37] , \p[9][36] , \p[9][35] ,
         \p[9][34] , \p[9][33] , \p[9][32] , \p[9][31] , \p[9][30] ,
         \p[9][29] , \p[9][28] , \p[9][27] , \p[9][26] , \p[9][25] ,
         \p[9][24] , \p[9][23] , \p[9][22] , \p[9][21] , \p[9][20] ,
         \p[9][19] , \p[9][18] , \p[9][17] , \p[9][16] , \p[9][15] ,
         \p[9][14] , \p[9][13] , \p[9][12] , \p[9][11] , \p[9][10] , \p[9][9] ,
         \p[8][63] , \p[8][38] , \p[8][37] , \p[8][36] , \p[8][35] ,
         \p[8][34] , \p[8][33] , \p[8][32] , \p[8][31] , \p[8][30] ,
         \p[8][29] , \p[8][28] , \p[8][27] , \p[8][26] , \p[8][25] ,
         \p[8][24] , \p[8][23] , \p[8][22] , \p[8][21] , \p[8][20] ,
         \p[8][19] , \p[8][18] , \p[8][17] , \p[8][16] , \p[8][15] ,
         \p[8][14] , \p[8][13] , \p[8][12] , \p[8][11] , \p[8][10] , \p[8][9] ,
         \p[8][8] , \g[41][63] , \g[41][62] , \g[41][61] , \g[41][60] ,
         \g[41][59] , \g[41][58] , \g[41][57] , \g[41][56] , \g[41][55] ,
         \g[41][54] , \g[41][53] , \g[41][52] , \g[41][51] , \g[41][50] ,
         \g[41][49] , \g[41][48] , \g[41][47] , \g[41][46] , \g[41][45] ,
         \g[41][44] , \g[41][43] , \g[41][42] , \g[41][41] , \g[41][40] ,
         \g[41][39] , \g[41][38] , \g[41][37] , \g[41][36] , \g[41][35] ,
         \g[41][34] , \g[41][33] , \g[41][32] , \g[41][31] , \g[41][30] ,
         \g[41][29] , \g[41][28] , \g[41][27] , \g[41][26] , \g[41][25] ,
         \g[41][24] , \g[41][23] , \g[41][22] , \g[41][21] , \g[41][20] ,
         \g[41][19] , \g[41][18] , \g[41][17] , \g[41][16] , \g[41][15] ,
         \g[41][14] , \g[41][13] , \g[41][12] , \g[41][11] , \g[41][10] ,
         \g[41][9] , \g[41][8] , \g[41][7] , \g[41][6] , \g[41][5] ,
         \g[41][4] , \g[41][3] , \g[41][2] , \g[41][1] , \g[40][63] ,
         \g[40][62] , \g[40][61] , \g[40][60] , \g[40][59] , \g[40][58] ,
         \g[40][57] , \g[40][56] , \g[40][55] , \g[40][54] , \g[40][53] ,
         \g[40][52] , \g[40][51] , \g[40][50] , \g[40][49] , \g[40][48] ,
         \g[40][47] , \g[40][46] , \g[40][45] , \g[40][44] , \g[40][43] ,
         \g[40][42] , \g[40][41] , \g[40][40] , \g[40][39] , \g[40][38] ,
         \g[40][37] , \g[40][36] , \g[40][35] , \g[40][34] , \g[40][33] ,
         \g[40][32] , \g[40][31] , \g[40][30] , \g[40][29] , \g[40][28] ,
         \g[40][27] , \g[40][26] , \g[40][25] , \g[40][24] , \g[40][23] ,
         \g[40][22] , \g[40][21] , \g[40][20] , \g[40][19] , \g[40][18] ,
         \g[40][17] , \g[40][16] , \g[40][15] , \g[40][14] , \g[40][13] ,
         \g[40][12] , \g[40][11] , \g[40][10] , \g[40][9] , \g[40][8] ,
         \g[40][7] , \g[40][6] , \g[40][5] , \g[40][4] , \g[40][3] ,
         \g[40][2] , \g[40][1] , \g[39][63] , \g[39][62] , \g[39][61] ,
         \g[39][60] , \g[39][59] , \g[39][58] , \g[39][57] , \g[39][56] ,
         \g[39][55] , \g[39][54] , \g[39][53] , \g[39][52] , \g[39][51] ,
         \g[39][50] , \g[39][49] , \g[39][48] , \g[39][47] , \g[39][46] ,
         \g[39][45] , \g[39][44] , \g[39][43] , \g[39][42] , \g[39][41] ,
         \g[39][40] , \g[39][39] , \g[39][38] , \g[39][37] , \g[39][36] ,
         \g[39][35] , \g[39][34] , \g[39][33] , \g[39][32] , \g[39][31] ,
         \g[39][30] , \g[39][29] , \g[39][28] , \g[39][27] , \g[39][26] ,
         \g[39][25] , \g[39][24] , \g[39][23] , \g[39][22] , \g[39][21] ,
         \g[39][20] , \g[39][19] , \g[39][18] , \g[39][17] , \g[39][16] ,
         \g[39][15] , \g[39][14] , \g[39][13] , \g[39][12] , \g[39][11] ,
         \g[39][10] , \g[39][9] , \g[39][8] , \g[39][7] , \g[39][6] ,
         \g[39][5] , \g[39][4] , \g[39][3] , \g[39][2] , \g[39][1] ,
         \g[38][63] , \g[38][62] , \g[38][61] , \g[38][60] , \g[38][59] ,
         \g[38][58] , \g[38][57] , \g[38][56] , \g[38][55] , \g[38][54] ,
         \g[38][53] , \g[38][52] , \g[38][51] , \g[38][50] , \g[38][49] ,
         \g[38][48] , \g[38][47] , \g[38][46] , \g[38][45] , \g[38][44] ,
         \g[38][43] , \g[38][42] , \g[38][41] , \g[38][40] , \g[38][39] ,
         \g[38][38] , \g[38][37] , \g[38][36] , \g[38][35] , \g[38][34] ,
         \g[38][33] , \g[38][32] , \g[38][31] , \g[38][30] , \g[38][29] ,
         \g[38][28] , \g[38][27] , \g[38][26] , \g[38][25] , \g[38][24] ,
         \g[38][23] , \g[38][22] , \g[38][21] , \g[38][20] , \g[38][19] ,
         \g[38][18] , \g[38][17] , \g[38][16] , \g[38][15] , \g[38][14] ,
         \g[38][13] , \g[38][12] , \g[38][11] , \g[38][10] , \g[38][9] ,
         \g[38][8] , \g[38][7] , \g[38][6] , \g[38][5] , \g[38][4] ,
         \g[38][3] , \g[38][2] , \g[38][1] , \g[37][63] , \g[37][62] ,
         \g[37][61] , \g[37][60] , \g[37][59] , \g[37][58] , \g[37][57] ,
         \g[37][56] , \g[37][55] , \g[37][54] , \g[37][53] , \g[37][52] ,
         \g[37][51] , \g[37][50] , \g[37][49] , \g[37][48] , \g[37][47] ,
         \g[37][46] , \g[37][45] , \g[37][44] , \g[37][43] , \g[37][42] ,
         \g[37][41] , \g[37][40] , \g[37][39] , \g[37][38] , \g[37][37] ,
         \g[37][36] , \g[37][35] , \g[37][34] , \g[37][33] , \g[37][32] ,
         \g[37][31] , \g[37][30] , \g[37][29] , \g[37][28] , \g[37][27] ,
         \g[37][26] , \g[37][25] , \g[37][24] , \g[37][23] , \g[37][22] ,
         \g[37][21] , \g[37][20] , \g[37][19] , \g[37][18] , \g[37][17] ,
         \g[37][16] , \g[37][15] , \g[37][14] , \g[37][13] , \g[37][12] ,
         \g[37][11] , \g[37][10] , \g[37][9] , \g[37][8] , \g[37][7] ,
         \g[37][6] , \g[37][5] , \g[37][4] , \g[37][3] , \g[37][2] ,
         \g[37][1] , \g[36][63] , \g[36][62] , \g[36][61] , \g[36][60] ,
         \g[36][59] , \g[36][58] , \g[36][57] , \g[36][56] , \g[36][55] ,
         \g[36][54] , \g[36][53] , \g[36][52] , \g[36][51] , \g[36][50] ,
         \g[36][49] , \g[36][48] , \g[36][47] , \g[36][46] , \g[36][45] ,
         \g[36][44] , \g[36][43] , \g[36][42] , \g[36][41] , \g[36][40] ,
         \g[36][39] , \g[36][38] , \g[36][37] , \g[36][36] , \g[36][35] ,
         \g[36][34] , \g[36][33] , \g[36][32] , \g[36][31] , \g[36][30] ,
         \g[36][29] , \g[36][28] , \g[36][27] , \g[36][26] , \g[36][25] ,
         \g[36][24] , \g[36][23] , \g[36][22] , \g[36][21] , \g[36][20] ,
         \g[36][19] , \g[36][18] , \g[36][17] , \g[36][16] , \g[36][15] ,
         \g[36][14] , \g[36][13] , \g[36][12] , \g[36][11] , \g[36][10] ,
         \g[36][9] , \g[36][8] , \g[36][7] , \g[36][6] , \g[36][5] ,
         \g[36][4] , \g[36][3] , \g[36][2] , \g[36][1] , \g[35][63] ,
         \g[35][62] , \g[35][61] , \g[35][60] , \g[35][59] , \g[35][58] ,
         \g[35][57] , \g[35][56] , \g[35][55] , \g[35][54] , \g[35][53] ,
         \g[35][52] , \g[35][51] , \g[35][50] , \g[35][49] , \g[35][48] ,
         \g[35][47] , \g[35][46] , \g[35][45] , \g[35][44] , \g[35][43] ,
         \g[35][42] , \g[35][41] , \g[35][40] , \g[35][39] , \g[35][38] ,
         \g[35][37] , \g[35][36] , \g[35][35] , \g[35][34] , \g[35][33] ,
         \g[35][32] , \g[35][31] , \g[35][30] , \g[35][29] , \g[35][28] ,
         \g[35][27] , \g[35][26] , \g[35][25] , \g[35][24] , \g[35][23] ,
         \g[35][22] , \g[35][21] , \g[35][20] , \g[35][19] , \g[35][18] ,
         \g[35][17] , \g[35][16] , \g[35][15] , \g[35][14] , \g[35][13] ,
         \g[35][12] , \g[35][11] , \g[35][10] , \g[35][9] , \g[35][8] ,
         \g[35][7] , \g[35][6] , \g[35][5] , \g[35][4] , \g[35][3] ,
         \g[35][2] , \g[35][1] , \g[34][63] , \g[34][62] , \g[34][61] ,
         \g[34][60] , \g[34][59] , \g[34][58] , \g[34][57] , \g[34][56] ,
         \g[34][55] , \g[34][54] , \g[34][53] , \g[34][52] , \g[34][51] ,
         \g[34][50] , \g[34][49] , \g[34][48] , \g[34][47] , \g[34][46] ,
         \g[34][45] , \g[34][44] , \g[34][43] , \g[34][42] , \g[34][41] ,
         \g[34][40] , \g[34][39] , \g[34][38] , \g[34][37] , \g[34][36] ,
         \g[34][35] , \g[34][34] , \g[34][33] , \g[34][32] , \g[34][31] ,
         \g[34][30] , \g[34][29] , \g[34][28] , \g[34][27] , \g[34][26] ,
         \g[34][25] , \g[34][24] , \g[34][23] , \g[34][22] , \g[34][21] ,
         \g[34][20] , \g[34][19] , \g[34][18] , \g[34][17] , \g[34][16] ,
         \g[34][15] , \g[34][14] , \g[34][13] , \g[34][12] , \g[34][11] ,
         \g[34][10] , \g[34][9] , \g[34][8] , \g[34][7] , \g[34][6] ,
         \g[34][5] , \g[34][4] , \g[34][3] , \g[34][2] , \g[34][1] ,
         \g[33][63] , \g[33][62] , \g[33][61] , \g[33][60] , \g[33][59] ,
         \g[33][58] , \g[33][57] , \g[33][56] , \g[33][55] , \g[33][54] ,
         \g[33][53] , \g[33][52] , \g[33][51] , \g[33][50] , \g[33][49] ,
         \g[33][48] , \g[33][47] , \g[33][46] , \g[33][45] , \g[33][44] ,
         \g[33][43] , \g[33][42] , \g[33][41] , \g[33][40] , \g[33][39] ,
         \g[33][38] , \g[33][37] , \g[33][36] , \g[33][35] , \g[33][34] ,
         \g[33][33] , \g[33][32] , \g[33][31] , \g[33][30] , \g[33][29] ,
         \g[33][28] , \g[33][27] , \g[33][26] , \g[33][25] , \g[33][24] ,
         \g[33][23] , \g[33][22] , \g[33][21] , \g[33][20] , \g[33][19] ,
         \g[33][18] , \g[33][17] , \g[33][16] , \g[33][15] , \g[33][14] ,
         \g[33][13] , \g[33][12] , \g[33][11] , \g[33][10] , \g[33][9] ,
         \g[33][8] , \g[33][7] , \g[33][6] , \g[33][5] , \g[33][4] ,
         \g[33][3] , \g[33][2] , \g[33][1] , \g[32][63] , \g[32][62] ,
         \g[32][61] , \g[32][60] , \g[32][59] , \g[32][58] , \g[32][57] ,
         \g[32][56] , \g[32][55] , \g[32][54] , \g[32][53] , \g[32][52] ,
         \g[32][51] , \g[32][50] , \g[32][49] , \g[32][48] , \g[32][47] ,
         \g[32][46] , \g[32][45] , \g[32][44] , \g[32][43] , \g[32][42] ,
         \g[32][41] , \g[32][40] , \g[32][39] , \g[32][38] , \g[32][37] ,
         \g[32][36] , \g[32][35] , \g[32][34] , \g[32][33] , \g[32][32] ,
         \g[32][31] , \g[32][30] , \g[32][29] , \g[32][28] , \g[32][27] ,
         \g[32][26] , \g[32][25] , \g[32][24] , \g[32][23] , \g[32][22] ,
         \g[32][21] , \g[32][20] , \g[32][19] , \g[32][18] , \g[32][17] ,
         \g[32][16] , \g[32][15] , \g[32][14] , \g[32][13] , \g[32][12] ,
         \g[32][11] , \g[32][10] , \g[32][9] , \g[32][8] , \g[32][7] ,
         \g[32][6] , \g[32][5] , \g[32][4] , \g[32][3] , \g[32][2] ,
         \g[32][1] , \g[31][63] , \g[31][62] , \g[31][61] , \g[31][60] ,
         \g[31][59] , \g[31][58] , \g[31][57] , \g[31][56] , \g[31][55] ,
         \g[31][54] , \g[31][53] , \g[31][52] , \g[31][51] , \g[31][50] ,
         \g[31][49] , \g[31][48] , \g[31][47] , \g[31][46] , \g[31][45] ,
         \g[31][44] , \g[31][43] , \g[31][42] , \g[31][41] , \g[31][40] ,
         \g[31][39] , \g[31][38] , \g[31][37] , \g[31][36] , \g[31][35] ,
         \g[31][34] , \g[31][33] , \g[31][32] , \g[31][31] , \g[31][30] ,
         \g[31][29] , \g[31][28] , \g[31][27] , \g[31][26] , \g[31][25] ,
         \g[31][24] , \g[31][23] , \g[31][22] , \g[31][21] , \g[31][20] ,
         \g[31][19] , \g[31][18] , \g[31][17] , \g[31][16] , \g[31][15] ,
         \g[31][14] , \g[31][13] , \g[31][12] , \g[31][11] , \g[31][10] ,
         \g[31][9] , \g[31][8] , \g[31][7] , \g[31][6] , \g[31][5] ,
         \g[31][4] , \g[31][3] , \g[31][2] , \g[31][1] , \g[30][63] ,
         \g[30][62] , \g[30][61] , \g[30][60] , \g[30][59] , \g[30][58] ,
         \g[30][57] , \g[30][56] , \g[30][55] , \g[30][54] , \g[30][53] ,
         \g[30][52] , \g[30][51] , \g[30][50] , \g[30][49] , \g[30][48] ,
         \g[30][47] , \g[30][46] , \g[30][45] , \g[30][44] , \g[30][43] ,
         \g[30][42] , \g[30][41] , \g[30][40] , \g[30][39] , \g[30][38] ,
         \g[30][37] , \g[30][36] , \g[30][35] , \g[30][34] , \g[30][33] ,
         \g[30][32] , \g[30][31] , \g[30][30] , \g[30][29] , \g[30][28] ,
         \g[30][27] , \g[30][26] , \g[30][25] , \g[30][24] , \g[30][23] ,
         \g[30][22] , \g[30][21] , \g[30][20] , \g[30][19] , \g[30][18] ,
         \g[30][17] , \g[30][16] , \g[30][15] , \g[30][14] , \g[30][13] ,
         \g[30][12] , \g[30][11] , \g[30][10] , \g[30][9] , \g[30][8] ,
         \g[30][7] , \g[30][6] , \g[30][5] , \g[30][4] , \g[30][3] ,
         \g[30][2] , \g[30][1] , \g[29][63] , \g[29][62] , \g[29][61] ,
         \g[29][60] , \g[29][59] , \g[29][58] , \g[29][57] , \g[29][56] ,
         \g[29][55] , \g[29][54] , \g[29][53] , \g[29][52] , \g[29][51] ,
         \g[29][50] , \g[29][49] , \g[29][48] , \g[29][47] , \g[29][46] ,
         \g[29][45] , \g[29][44] , \g[29][43] , \g[29][42] , \g[29][41] ,
         \g[29][40] , \g[29][39] , \g[29][38] , \g[29][37] , \g[29][36] ,
         \g[29][35] , \g[29][34] , \g[29][33] , \g[29][32] , \g[29][31] ,
         \g[29][30] , \g[29][29] , \g[29][28] , \g[29][27] , \g[29][26] ,
         \g[29][25] , \g[29][24] , \g[29][23] , \g[29][22] , \g[29][21] ,
         \g[29][20] , \g[29][19] , \g[29][18] , \g[29][17] , \g[29][16] ,
         \g[29][15] , \g[29][14] , \g[29][13] , \g[29][12] , \g[29][11] ,
         \g[29][10] , \g[29][9] , \g[29][8] , \g[29][7] , \g[29][6] ,
         \g[29][5] , \g[29][4] , \g[29][3] , \g[29][2] , \g[29][1] ,
         \g[28][63] , \g[28][62] , \g[28][61] , \g[28][60] , \g[28][59] ,
         \g[28][58] , \g[28][57] , \g[28][56] , \g[28][55] , \g[28][54] ,
         \g[28][53] , \g[28][52] , \g[28][51] , \g[28][50] , \g[28][49] ,
         \g[28][48] , \g[28][47] , \g[28][46] , \g[28][45] , \g[28][44] ,
         \g[28][43] , \g[28][42] , \g[28][41] , \g[28][40] , \g[28][39] ,
         \g[28][38] , \g[28][37] , \g[28][36] , \g[28][35] , \g[28][34] ,
         \g[28][33] , \g[28][32] , \g[28][31] , \g[28][30] , \g[28][29] ,
         \g[28][28] , \g[28][27] , \g[28][26] , \g[28][25] , \g[28][24] ,
         \g[28][23] , \g[28][22] , \g[28][21] , \g[28][20] , \g[28][19] ,
         \g[28][18] , \g[28][17] , \g[28][16] , \g[28][15] , \g[28][14] ,
         \g[28][13] , \g[28][12] , \g[28][11] , \g[28][10] , \g[28][9] ,
         \g[28][8] , \g[28][7] , \g[28][6] , \g[28][5] , \g[28][4] ,
         \g[28][3] , \g[28][2] , \g[28][1] , \g[27][63] , \g[27][62] ,
         \g[27][61] , \g[27][60] , \g[27][59] , \g[27][58] , \g[27][57] ,
         \g[27][56] , \g[27][55] , \g[27][54] , \g[27][53] , \g[27][52] ,
         \g[27][51] , \g[27][50] , \g[27][49] , \g[27][48] , \g[27][47] ,
         \g[27][46] , \g[27][45] , \g[27][44] , \g[27][43] , \g[27][42] ,
         \g[27][41] , \g[27][40] , \g[27][39] , \g[27][38] , \g[27][37] ,
         \g[27][36] , \g[27][35] , \g[27][34] , \g[27][33] , \g[27][32] ,
         \g[27][31] , \g[27][30] , \g[27][29] , \g[27][28] , \g[27][27] ,
         \g[27][26] , \g[27][25] , \g[27][24] , \g[27][23] , \g[27][22] ,
         \g[27][21] , \g[27][20] , \g[27][19] , \g[27][18] , \g[27][17] ,
         \g[27][16] , \g[27][15] , \g[27][14] , \g[27][13] , \g[27][12] ,
         \g[27][11] , \g[27][10] , \g[27][9] , \g[27][8] , \g[27][7] ,
         \g[27][6] , \g[27][5] , \g[27][4] , \g[27][3] , \g[27][2] ,
         \g[27][1] , \g[26][63] , \g[26][62] , \g[26][61] , \g[26][60] ,
         \g[26][59] , \g[26][58] , \g[26][57] , \g[26][56] , \g[26][55] ,
         \g[26][54] , \g[26][53] , \g[26][52] , \g[26][51] , \g[26][50] ,
         \g[26][49] , \g[26][48] , \g[26][47] , \g[26][46] , \g[26][45] ,
         \g[26][44] , \g[26][43] , \g[26][42] , \g[26][41] , \g[26][40] ,
         \g[26][39] , \g[26][38] , \g[26][37] , \g[26][36] , \g[26][35] ,
         \g[26][34] , \g[26][33] , \g[26][32] , \g[26][31] , \g[26][30] ,
         \g[26][29] , \g[26][28] , \g[26][27] , \g[26][26] , \g[26][25] ,
         \g[26][24] , \g[26][23] , \g[26][22] , \g[26][21] , \g[26][20] ,
         \g[26][19] , \g[26][18] , \g[26][17] , \g[26][16] , \g[26][15] ,
         \g[26][14] , \g[26][13] , \g[26][12] , \g[26][11] , \g[26][10] ,
         \g[26][9] , \g[26][8] , \g[26][7] , \g[26][6] , \g[26][5] ,
         \g[26][4] , \g[26][3] , \g[26][2] , \g[26][1] , \g[25][63] ,
         \g[25][62] , \g[25][61] , \g[25][60] , \g[25][59] , \g[25][58] ,
         \g[25][57] , \g[25][56] , \g[25][55] , \g[25][54] , \g[25][53] ,
         \g[25][52] , \g[25][51] , \g[25][50] , \g[25][49] , \g[25][48] ,
         \g[25][47] , \g[25][46] , \g[25][45] , \g[25][44] , \g[25][43] ,
         \g[25][42] , \g[25][41] , \g[25][40] , \g[25][39] , \g[25][38] ,
         \g[25][37] , \g[25][36] , \g[25][35] , \g[25][34] , \g[25][33] ,
         \g[25][32] , \g[25][31] , \g[25][30] , \g[25][29] , \g[25][28] ,
         \g[25][27] , \g[25][26] , \g[25][25] , \g[25][24] , \g[25][23] ,
         \g[25][22] , \g[25][21] , \g[25][20] , \g[25][19] , \g[25][18] ,
         \g[25][17] , \g[25][16] , \g[25][15] , \g[25][14] , \g[25][13] ,
         \g[25][12] , \g[25][11] , \g[25][10] , \g[25][9] , \g[25][8] ,
         \g[25][7] , \g[25][6] , \g[25][5] , \g[25][4] , \g[25][3] ,
         \g[25][2] , \g[25][1] , \g[24][63] , \g[24][62] , \g[24][61] ,
         \g[24][60] , \g[24][59] , \g[24][58] , \g[24][57] , \g[24][56] ,
         \g[24][55] , \g[24][54] , \g[24][53] , \g[24][52] , \g[24][51] ,
         \g[24][50] , \g[24][49] , \g[24][48] , \g[24][47] , \g[24][46] ,
         \g[24][45] , \g[24][44] , \g[24][43] , \g[24][42] , \g[24][41] ,
         \g[24][40] , \g[24][39] , \g[24][38] , \g[24][37] , \g[24][36] ,
         \g[24][35] , \g[24][34] , \g[24][33] , \g[24][32] , \g[24][31] ,
         \g[24][30] , \g[24][29] , \g[24][28] , \g[24][27] , \g[24][26] ,
         \g[24][25] , \g[24][24] , \g[24][23] , \g[24][22] , \g[24][21] ,
         \g[24][20] , \g[24][19] , \g[24][18] , \g[24][17] , \g[24][16] ,
         \g[24][15] , \g[24][14] , \g[24][13] , \g[24][12] , \g[24][11] ,
         \g[24][10] , \g[24][9] , \g[24][8] , \g[24][7] , \g[24][6] ,
         \g[24][5] , \g[24][4] , \g[24][3] , \g[24][2] , \g[24][1] ,
         \g[23][63] , \g[23][62] , \g[23][61] , \g[23][60] , \g[23][59] ,
         \g[23][58] , \g[23][57] , \g[23][56] , \g[23][55] , \g[23][54] ,
         \g[23][53] , \g[23][52] , \g[23][51] , \g[23][50] , \g[23][49] ,
         \g[23][48] , \g[23][47] , \g[23][46] , \g[23][45] , \g[23][44] ,
         \g[23][43] , \g[23][42] , \g[23][41] , \g[23][40] , \g[23][39] ,
         \g[23][38] , \g[23][37] , \g[23][36] , \g[23][35] , \g[23][34] ,
         \g[23][33] , \g[23][32] , \g[23][31] , \g[23][30] , \g[23][29] ,
         \g[23][28] , \g[23][27] , \g[23][26] , \g[23][25] , \g[23][24] ,
         \g[23][23] , \g[23][22] , \g[23][21] , \g[23][20] , \g[23][19] ,
         \g[23][18] , \g[23][17] , \g[23][16] , \g[23][15] , \g[23][14] ,
         \g[23][13] , \g[23][12] , \g[23][11] , \g[23][10] , \g[23][9] ,
         \g[23][8] , \g[23][7] , \g[23][6] , \g[23][5] , \g[23][4] ,
         \g[23][3] , \g[23][2] , \g[23][1] , \g[22][63] , \g[22][62] ,
         \g[22][61] , \g[22][60] , \g[22][59] , \g[22][58] , \g[22][57] ,
         \g[22][56] , \g[22][55] , \g[22][54] , \g[22][53] , \g[22][52] ,
         \g[22][51] , \g[22][50] , \g[22][49] , \g[22][48] , \g[22][47] ,
         \g[22][46] , \g[22][45] , \g[22][44] , \g[22][43] , \g[22][42] ,
         \g[22][41] , \g[22][40] , \g[22][39] , \g[22][38] , \g[22][37] ,
         \g[22][36] , \g[22][35] , \g[22][34] , \g[22][33] , \g[22][32] ,
         \g[22][31] , \g[22][30] , \g[22][29] , \g[22][28] , \g[22][27] ,
         \g[22][26] , \g[22][25] , \g[22][24] , \g[22][23] , \g[22][22] ,
         \g[22][21] , \g[22][20] , \g[22][19] , \g[22][18] , \g[22][17] ,
         \g[22][16] , \g[22][15] , \g[22][14] , \g[22][13] , \g[22][12] ,
         \g[22][11] , \g[22][10] , \g[22][9] , \g[22][8] , \g[22][7] ,
         \g[22][6] , \g[22][5] , \g[22][4] , \g[22][3] , \g[22][2] ,
         \g[22][1] , \g[21][63] , \g[21][62] , \g[21][61] , \g[21][60] ,
         \g[21][59] , \g[21][58] , \g[21][57] , \g[21][56] , \g[21][55] ,
         \g[21][54] , \g[21][53] , \g[21][52] , \g[21][51] , \g[21][50] ,
         \g[21][49] , \g[21][48] , \g[21][47] , \g[21][46] , \g[21][45] ,
         \g[21][44] , \g[21][43] , \g[21][42] , \g[21][41] , \g[21][40] ,
         \g[21][39] , \g[21][38] , \g[21][37] , \g[21][36] , \g[21][35] ,
         \g[21][34] , \g[21][33] , \g[21][32] , \g[21][31] , \g[21][30] ,
         \g[21][29] , \g[21][28] , \g[21][27] , \g[21][26] , \g[21][25] ,
         \g[21][24] , \g[21][23] , \g[21][22] , \g[21][21] , \g[21][20] ,
         \g[21][19] , \g[21][18] , \g[21][17] , \g[21][16] , \g[21][15] ,
         \g[21][14] , \g[21][13] , \g[21][12] , \g[21][11] , \g[21][10] ,
         \g[21][9] , \g[21][8] , \g[21][7] , \g[21][6] , \g[21][5] ,
         \g[21][4] , \g[21][3] , \g[21][2] , \g[21][1] , \g[20][63] ,
         \g[20][62] , \g[20][61] , \g[20][60] , \g[20][59] , \g[20][58] ,
         \g[20][57] , \g[20][56] , \g[20][55] , \g[20][54] , \g[20][53] ,
         \g[20][52] , \g[20][51] , \g[20][50] , \g[20][49] , \g[20][48] ,
         \g[20][47] , \g[20][46] , \g[20][45] , \g[20][44] , \g[20][43] ,
         \g[20][42] , \g[20][41] , \g[20][40] , \g[20][39] , \g[20][38] ,
         \g[20][37] , \g[20][36] , \g[20][35] , \g[20][34] , \g[20][33] ,
         \g[20][32] , \g[20][31] , \g[20][30] , \g[20][29] , \g[20][28] ,
         \g[20][27] , \g[20][26] , \g[20][25] , \g[20][24] , \g[20][23] ,
         \g[20][22] , \g[20][21] , \g[20][20] , \g[20][19] , \g[20][18] ,
         \g[20][17] , \g[20][16] , \g[20][15] , \g[20][14] , \g[20][13] ,
         \g[20][12] , \g[20][11] , \g[20][10] , \g[20][9] , \g[20][8] ,
         \g[20][7] , \g[20][6] , \g[20][5] , \g[20][4] , \g[20][3] ,
         \g[20][2] , \g[20][1] , \g[20][0] , \g[19][63] , \g[19][62] ,
         \g[19][61] , \g[19][60] , \g[19][59] , \g[19][58] , \g[19][57] ,
         \g[19][56] , \g[19][55] , \g[19][54] , \g[19][53] , \g[19][52] ,
         \g[19][51] , \g[19][50] , \g[19][49] , \g[19][48] , \g[19][47] ,
         \g[19][46] , \g[19][45] , \g[19][44] , \g[19][43] , \g[19][42] ,
         \g[19][41] , \g[19][40] , \g[19][39] , \g[19][38] , \g[19][37] ,
         \g[19][36] , \g[19][35] , \g[19][34] , \g[19][33] , \g[19][32] ,
         \g[19][31] , \g[19][30] , \g[19][29] , \g[19][28] , \g[19][27] ,
         \g[19][26] , \g[19][25] , \g[19][24] , \g[19][23] , \g[19][22] ,
         \g[19][21] , \g[19][20] , \g[19][19] , \g[19][18] , \g[19][17] ,
         \g[19][16] , \g[19][15] , \g[19][14] , \g[19][13] , \g[19][12] ,
         \g[19][11] , \g[19][10] , \g[19][9] , \g[19][8] , \g[19][7] ,
         \g[19][6] , \g[19][5] , \g[19][4] , \g[19][3] , \g[19][2] ,
         \g[19][1] , \g[19][0] , \g[18][63] , \g[18][62] , \g[18][61] ,
         \g[18][60] , \g[18][59] , \g[18][58] , \g[18][57] , \g[18][56] ,
         \g[18][55] , \g[18][54] , \g[18][53] , \g[18][52] , \g[18][51] ,
         \g[18][50] , \g[18][49] , \g[18][48] , \g[18][47] , \g[18][46] ,
         \g[18][45] , \g[18][44] , \g[18][43] , \g[18][42] , \g[18][41] ,
         \g[18][40] , \g[18][39] , \g[18][38] , \g[18][37] , \g[18][36] ,
         \g[18][35] , \g[18][34] , \g[18][33] , \g[18][32] , \g[18][31] ,
         \g[18][30] , \g[18][29] , \g[18][28] , \g[18][27] , \g[18][26] ,
         \g[18][25] , \g[18][24] , \g[18][23] , \g[18][22] , \g[18][21] ,
         \g[18][20] , \g[18][19] , \g[18][18] , \g[18][17] , \g[18][16] ,
         \g[18][15] , \g[18][14] , \g[18][13] , \g[18][12] , \g[18][11] ,
         \g[18][10] , \g[18][9] , \g[18][8] , \g[18][7] , \g[18][6] ,
         \g[18][5] , \g[18][4] , \g[18][3] , \g[18][2] , \g[18][1] ,
         \g[18][0] , \g[17][63] , \g[17][62] , \g[17][61] , \g[17][60] ,
         \g[17][59] , \g[17][58] , \g[17][57] , \g[17][56] , \g[17][55] ,
         \g[17][54] , \g[17][53] , \g[17][52] , \g[17][51] , \g[17][50] ,
         \g[17][49] , \g[17][48] , \g[17][47] , \g[17][46] , \g[17][45] ,
         \g[17][44] , \g[17][43] , \g[17][42] , \g[17][41] , \g[17][40] ,
         \g[17][39] , \g[17][38] , \g[17][37] , \g[17][36] , \g[17][35] ,
         \g[17][34] , \g[17][33] , \g[17][32] , \g[17][31] , \g[17][30] ,
         \g[17][29] , \g[17][28] , \g[17][27] , \g[17][26] , \g[17][25] ,
         \g[17][24] , \g[17][23] , \g[17][22] , \g[17][21] , \g[17][20] ,
         \g[17][19] , \g[17][18] , \g[17][17] , \g[17][16] , \g[17][15] ,
         \g[17][14] , \g[17][13] , \g[17][12] , \g[17][11] , \g[17][10] ,
         \g[17][9] , \g[17][8] , \g[17][7] , \g[17][6] , \g[17][5] ,
         \g[17][4] , \g[17][3] , \g[17][2] , \g[17][1] , \g[17][0] ,
         \g[16][63] , \g[16][62] , \g[16][61] , \g[16][60] , \g[16][59] ,
         \g[16][58] , \g[16][57] , \g[16][56] , \g[16][55] , \g[16][54] ,
         \g[16][53] , \g[16][52] , \g[16][51] , \g[16][50] , \g[16][49] ,
         \g[16][48] , \g[16][47] , \g[16][46] , \g[16][45] , \g[16][44] ,
         \g[16][43] , \g[16][42] , \g[16][41] , \g[16][40] , \g[16][39] ,
         \g[16][38] , \g[16][37] , \g[16][36] , \g[16][35] , \g[16][34] ,
         \g[16][33] , \g[16][32] , \g[16][31] , \g[16][30] , \g[16][29] ,
         \g[16][28] , \g[16][27] , \g[16][26] , \g[16][25] , \g[16][24] ,
         \g[16][23] , \g[16][22] , \g[16][21] , \g[16][20] , \g[16][19] ,
         \g[16][18] , \g[16][17] , \g[16][16] , \g[16][15] , \g[16][14] ,
         \g[16][13] , \g[16][12] , \g[16][11] , \g[16][10] , \g[16][9] ,
         \g[16][8] , \g[16][7] , \g[16][6] , \g[16][5] , \g[16][4] ,
         \g[16][3] , \g[16][2] , \g[16][1] , \g[16][0] , \g[15][63] ,
         \g[15][62] , \g[15][61] , \g[15][60] , \g[15][59] , \g[15][58] ,
         \g[15][57] , \g[15][56] , \g[15][55] , \g[15][54] , \g[15][53] ,
         \g[15][52] , \g[15][51] , \g[15][50] , \g[15][49] , \g[15][48] ,
         \g[15][47] , \g[15][46] , \g[15][45] , \g[15][44] , \g[15][43] ,
         \g[15][42] , \g[15][41] , \g[15][40] , \g[15][39] , \g[15][38] ,
         \g[15][37] , \g[15][36] , \g[15][35] , \g[15][34] , \g[15][33] ,
         \g[15][32] , \g[15][31] , \g[15][30] , \g[15][29] , \g[15][28] ,
         \g[15][27] , \g[15][26] , \g[15][25] , \g[15][24] , \g[15][23] ,
         \g[15][22] , \g[15][21] , \g[15][20] , \g[15][19] , \g[15][18] ,
         \g[15][17] , \g[15][16] , \g[15][15] , \g[15][14] , \g[15][13] ,
         \g[15][12] , \g[15][11] , \g[15][10] , \g[15][9] , \g[15][8] ,
         \g[15][7] , \g[15][6] , \g[15][5] , \g[15][4] , \g[15][3] ,
         \g[15][2] , \g[15][1] , \g[15][0] , \g[14][63] , \g[14][62] ,
         \g[14][61] , \g[14][60] , \g[14][59] , \g[14][58] , \g[14][57] ,
         \g[14][56] , \g[14][55] , \g[14][54] , \g[14][53] , \g[14][52] ,
         \g[14][51] , \g[14][50] , \g[14][49] , \g[14][48] , \g[14][47] ,
         \g[14][46] , \g[14][45] , \g[14][44] , \g[14][43] , \g[14][42] ,
         \g[14][41] , \g[14][40] , \g[14][39] , \g[14][38] , \g[14][37] ,
         \g[14][36] , \g[14][35] , \g[14][34] , \g[14][33] , \g[14][32] ,
         \g[14][31] , \g[14][30] , \g[14][29] , \g[14][28] , \g[14][27] ,
         \g[14][26] , \g[14][25] , \g[14][24] , \g[14][23] , \g[14][22] ,
         \g[14][21] , \g[14][20] , \g[14][19] , \g[14][18] , \g[14][17] ,
         \g[14][16] , \g[14][15] , \g[14][14] , \g[14][13] , \g[14][12] ,
         \g[14][11] , \g[14][10] , \g[14][9] , \g[14][8] , \g[14][7] ,
         \g[14][6] , \g[14][5] , \g[14][4] , \g[14][3] , \g[14][2] ,
         \g[14][1] , \g[14][0] , \g[13][63] , \g[13][62] , \g[13][61] ,
         \g[13][60] , \g[13][59] , \g[13][58] , \g[13][57] , \g[13][56] ,
         \g[13][55] , \g[13][54] , \g[13][53] , \g[13][52] , \g[13][51] ,
         \g[13][50] , \g[13][49] , \g[13][48] , \g[13][47] , \g[13][46] ,
         \g[13][45] , \g[13][44] , \g[13][43] , \g[13][42] , \g[13][41] ,
         \g[13][40] , \g[13][39] , \g[13][38] , \g[13][37] , \g[13][36] ,
         \g[13][35] , \g[13][34] , \g[13][33] , \g[13][32] , \g[13][31] ,
         \g[13][30] , \g[13][29] , \g[13][28] , \g[13][27] , \g[13][26] ,
         \g[13][25] , \g[13][24] , \g[13][23] , \g[13][22] , \g[13][21] ,
         \g[13][20] , \g[13][19] , \g[13][18] , \g[13][17] , \g[13][16] ,
         \g[13][15] , \g[13][14] , \g[13][13] , \g[13][12] , \g[13][11] ,
         \g[13][10] , \g[13][9] , \g[13][8] , \g[13][7] , \g[13][6] ,
         \g[13][5] , \g[13][4] , \g[13][3] , \g[13][2] , \g[13][1] ,
         \g[13][0] , \g[12][63] , \g[12][62] , \g[12][61] , \g[12][60] ,
         \g[12][59] , \g[12][58] , \g[12][57] , \g[12][56] , \g[12][55] ,
         \g[12][54] , \g[12][53] , \g[12][52] , \g[12][51] , \g[12][50] ,
         \g[12][49] , \g[12][48] , \g[12][47] , \g[12][46] , \g[12][45] ,
         \g[12][44] , \g[12][43] , \g[12][42] , \g[12][41] , \g[12][40] ,
         \g[12][39] , \g[12][38] , \g[12][37] , \g[12][36] , \g[12][35] ,
         \g[12][34] , \g[12][33] , \g[12][32] , \g[12][31] , \g[12][30] ,
         \g[12][29] , \g[12][28] , \g[12][27] , \g[12][26] , \g[12][25] ,
         \g[12][24] , \g[12][23] , \g[12][22] , \g[12][21] , \g[12][20] ,
         \g[12][19] , \g[12][18] , \g[12][17] , \g[12][16] , \g[12][15] ,
         \g[12][14] , \g[12][13] , \g[12][12] , \g[12][11] , \g[12][10] ,
         \g[12][9] , \g[12][8] , \g[12][7] , \g[12][6] , \g[12][5] ,
         \g[12][4] , \g[12][3] , \g[12][2] , \g[12][1] , \g[12][0] ,
         \g[11][63] , \g[11][62] , \g[11][61] , \g[11][60] , \g[11][59] ,
         \g[11][58] , \g[11][57] , \g[11][56] , \g[11][55] , \g[11][54] ,
         \g[11][53] , \g[11][52] , \g[11][51] , \g[11][50] , \g[11][49] ,
         \g[11][48] , \g[11][47] , \g[11][46] , \g[11][45] , \g[11][44] ,
         \g[11][43] , \g[11][42] , \g[11][41] , \g[11][40] , \g[11][39] ,
         \g[11][38] , \g[11][37] , \g[11][36] , \g[11][35] , \g[11][34] ,
         \g[11][33] , \g[11][32] , \g[11][31] , \g[11][30] , \g[11][29] ,
         \g[11][28] , \g[11][27] , \g[11][26] , \g[11][25] , \g[11][24] ,
         \g[11][23] , \g[11][22] , \g[11][21] , \g[11][20] , \g[11][19] ,
         \g[11][18] , \g[11][17] , \g[11][16] , \g[11][15] , \g[11][14] ,
         \g[11][13] , \g[11][12] , \g[11][11] , \g[11][10] , \g[11][9] ,
         \g[11][8] , \g[11][7] , \g[11][6] , \g[11][5] , \g[11][4] ,
         \g[11][3] , \g[11][2] , \g[11][1] , \g[11][0] , \g[10][63] ,
         \g[10][62] , \g[10][61] , \g[10][60] , \g[10][59] , \g[10][58] ,
         \g[10][57] , \g[10][56] , \g[10][55] , \g[10][54] , \g[10][53] ,
         \g[10][52] , \g[10][51] , \g[10][50] , \g[10][49] , \g[10][48] ,
         \g[10][47] , \g[10][46] , \g[10][45] , \g[10][44] , \g[10][43] ,
         \g[10][42] , \g[10][41] , \g[10][40] , \g[10][39] , \g[10][38] ,
         \g[10][37] , \g[10][36] , \g[10][35] , \g[10][34] , \g[10][33] ,
         \g[10][32] , \g[10][31] , \g[10][30] , \g[10][29] , \g[10][28] ,
         \g[10][27] , \g[10][26] , \g[10][25] , \g[10][24] , \g[10][23] ,
         \g[10][22] , \g[10][21] , \g[10][20] , \g[10][19] , \g[10][18] ,
         \g[10][17] , \g[10][16] , \g[10][15] , \g[10][14] , \g[10][13] ,
         \g[10][12] , \g[10][11] , \g[10][10] , \g[10][9] , \g[10][8] ,
         \g[10][7] , \g[10][6] , \g[10][5] , \g[10][4] , \g[10][3] ,
         \g[10][2] , \g[10][1] , \g[10][0] , \g[9][63] , \g[9][62] ,
         \g[9][61] , \g[9][60] , \g[9][59] , \g[9][58] , \g[9][57] ,
         \g[9][56] , \g[9][55] , \g[9][54] , \g[9][53] , \g[9][52] ,
         \g[9][51] , \g[9][50] , \g[9][49] , \g[9][48] , \g[9][47] ,
         \g[9][46] , \g[9][45] , \g[9][44] , \g[9][43] , \g[9][42] ,
         \g[9][41] , \g[9][40] , \g[9][39] , \g[9][38] , \g[9][37] ,
         \g[9][36] , \g[9][35] , \g[9][34] , \g[9][33] , \g[9][32] ,
         \g[9][31] , \g[9][30] , \g[9][29] , \g[9][28] , \g[9][27] ,
         \g[9][26] , \g[9][25] , \g[9][24] , \g[9][23] , \g[9][22] ,
         \g[9][21] , \g[9][20] , \g[9][19] , \g[9][18] , \g[9][17] ,
         \g[9][16] , \g[9][15] , \g[9][14] , \g[9][13] , \g[9][12] ,
         \g[9][11] , \g[9][10] , \g[9][9] , \g[9][8] , \g[9][7] , \g[9][6] ,
         \g[9][5] , \g[9][4] , \g[9][3] , \g[9][2] , \g[9][1] , \g[9][0] ,
         \g[8][63] , \g[8][62] , \g[8][61] , \g[8][60] , \g[8][59] ,
         \g[8][58] , \g[8][57] , \g[8][56] , \g[8][55] , \g[8][54] ,
         \g[8][53] , \g[8][52] , \g[8][51] , \g[8][50] , \g[8][49] ,
         \g[8][48] , \g[8][47] , \g[8][46] , \g[8][45] , \g[8][44] ,
         \g[8][43] , \g[8][42] , \g[8][41] , \g[8][40] , \g[8][39] ,
         \g[8][38] , \g[8][37] , \g[8][36] , \g[8][35] , \g[8][34] ,
         \g[8][33] , \g[8][32] , \g[8][31] , \g[8][30] , \g[8][29] ,
         \g[8][28] , \g[8][27] , \g[8][26] , \g[8][25] , \g[8][24] ,
         \g[8][23] , \g[8][22] , \g[8][21] , \g[8][20] , \g[8][19] ,
         \g[8][18] , \g[8][17] , \g[8][16] , \g[8][15] , \g[8][14] ,
         \g[8][13] , \g[8][12] , \g[8][11] , \g[8][10] , \g[8][9] , \g[8][8] ,
         \g[8][7] , \g[8][6] , \g[8][5] , \g[8][4] , \g[8][3] , \g[8][2] ,
         \g[8][1] , \g[8][0] , \g[7][63] , \g[7][62] , \g[7][61] , \g[7][60] ,
         \g[7][59] , \g[7][58] , \g[7][57] , \g[7][56] , \g[7][55] ,
         \g[7][54] , \g[7][53] , \g[7][52] , \g[7][51] , \g[7][50] ,
         \g[7][49] , \g[7][48] , \g[7][47] , \g[7][46] , \g[7][45] ,
         \g[7][44] , \g[7][43] , \g[7][42] , \g[7][41] , \g[7][40] ,
         \g[7][39] , \g[7][38] , \g[7][37] , \g[7][36] , \g[7][35] ,
         \g[7][34] , \g[7][33] , \g[7][32] , \g[7][31] , \g[7][30] ,
         \g[7][29] , \g[7][28] , \g[7][27] , \g[7][26] , \g[7][25] ,
         \g[7][24] , \g[7][23] , \g[7][22] , \g[7][21] , \g[7][20] ,
         \g[7][19] , \g[7][18] , \g[7][17] , \g[7][16] , \g[7][15] ,
         \g[7][14] , \g[7][13] , \g[7][12] , \g[7][11] , \g[7][10] , \g[7][9] ,
         \g[7][8] , \g[7][7] , \g[7][6] , \g[7][5] , \g[7][4] , \g[7][3] ,
         \g[7][2] , \g[7][1] , \g[7][0] , \g[6][63] , \g[6][62] , \g[6][61] ,
         \g[6][60] , \g[6][59] , \g[6][58] , \g[6][57] , \g[6][56] ,
         \g[6][55] , \g[6][54] , \g[6][53] , \g[6][52] , \g[6][51] ,
         \g[6][50] , \g[6][49] , \g[6][48] , \g[6][47] , \g[6][46] ,
         \g[6][45] , \g[6][44] , \g[6][43] , \g[6][42] , \g[6][41] ,
         \g[6][40] , \g[6][39] , \g[6][38] , \g[6][37] , \g[6][36] ,
         \g[6][35] , \g[6][34] , \g[6][33] , \g[6][32] , \g[6][31] ,
         \g[6][30] , \g[6][29] , \g[6][28] , \g[6][27] , \g[6][26] ,
         \g[6][25] , \g[6][24] , \g[6][23] , \g[6][22] , \g[6][21] ,
         \g[6][20] , \g[6][19] , \g[6][18] , \g[6][17] , \g[6][16] ,
         \g[6][15] , \g[6][14] , \g[6][13] , \g[6][12] , \g[6][11] ,
         \g[6][10] , \g[6][9] , \g[6][8] , \g[6][7] , \g[6][6] , \g[6][5] ,
         \g[6][4] , \g[6][3] , \g[6][2] , \g[6][1] , \g[6][0] , \g[5][63] ,
         \g[5][62] , \g[5][61] , \g[5][60] , \g[5][59] , \g[5][58] ,
         \g[5][57] , \g[5][56] , \g[5][55] , \g[5][54] , \g[5][53] ,
         \g[5][52] , \g[5][51] , \g[5][50] , \g[5][49] , \g[5][48] ,
         \g[5][47] , \g[5][46] , \g[5][45] , \g[5][44] , \g[5][43] ,
         \g[5][42] , \g[5][41] , \g[5][40] , \g[5][39] , \g[5][38] ,
         \g[5][37] , \g[5][36] , \g[5][35] , \g[5][34] , \g[5][33] ,
         \g[5][32] , \g[5][31] , \g[5][30] , \g[5][29] , \g[5][28] ,
         \g[5][27] , \g[5][26] , \g[5][25] , \g[5][24] , \g[5][23] ,
         \g[5][22] , \g[5][21] , \g[5][20] , \g[5][19] , \g[5][18] ,
         \g[5][17] , \g[5][16] , \g[5][15] , \g[5][14] , \g[5][13] ,
         \g[5][12] , \g[5][11] , \g[5][10] , \g[5][9] , \g[5][8] , \g[5][7] ,
         \g[5][6] , \g[5][5] , \g[5][4] , \g[5][3] , \g[5][2] , \g[5][1] ,
         \g[5][0] , \g[4][63] , \g[4][62] , \g[4][61] , \g[4][60] , \g[4][59] ,
         \g[4][58] , \g[4][57] , \g[4][56] , \g[4][55] , \g[4][54] ,
         \g[4][53] , \g[4][52] , \g[4][51] , \g[4][50] , \g[4][49] ,
         \g[4][48] , \g[4][47] , \g[4][46] , \g[4][45] , \g[4][44] ,
         \g[4][43] , \g[4][42] , \g[4][41] , \g[4][40] , \g[4][39] ,
         \g[4][38] , \g[4][37] , \g[4][36] , \g[4][35] , \g[4][34] ,
         \g[4][33] , \g[4][32] , \g[4][31] , \g[4][30] , \g[4][29] ,
         \g[4][28] , \g[4][27] , \g[4][26] , \g[4][25] , \g[4][24] ,
         \g[4][23] , \g[4][22] , \g[4][21] , \g[4][20] , \g[4][19] ,
         \g[4][18] , \g[4][17] , \g[4][16] , \g[4][15] , \g[4][14] ,
         \g[4][13] , \g[4][12] , \g[4][11] , \g[4][10] , \g[4][9] , \g[4][8] ,
         \g[4][7] , \g[4][6] , \g[4][5] , \g[4][4] , \g[4][3] , \g[4][2] ,
         \g[4][1] , \g[4][0] , \g[3][63] , \g[3][62] , \g[3][61] , \g[3][60] ,
         \g[3][59] , \g[3][58] , \g[3][57] , \g[3][56] , \g[3][55] ,
         \g[3][54] , \g[3][53] , \g[3][52] , \g[3][51] , \g[3][50] ,
         \g[3][49] , \g[3][48] , \g[3][47] , \g[3][46] , \g[3][45] ,
         \g[3][44] , \g[3][43] , \g[3][42] , \g[3][41] , \g[3][40] ,
         \g[3][39] , \g[3][38] , \g[3][37] , \g[3][36] , \g[3][35] ,
         \g[3][34] , \g[3][33] , \g[3][32] , \g[3][31] , \g[3][30] ,
         \g[3][29] , \g[3][28] , \g[3][27] , \g[3][26] , \g[3][25] ,
         \g[3][24] , \g[3][23] , \g[3][22] , \g[3][21] , \g[3][20] ,
         \g[3][19] , \g[3][18] , \g[3][17] , \g[3][16] , \g[3][15] ,
         \g[3][14] , \g[3][13] , \g[3][12] , \g[3][11] , \g[3][10] , \g[3][9] ,
         \g[3][8] , \g[3][7] , \g[3][6] , \g[3][5] , \g[3][4] , \g[3][3] ,
         \g[3][2] , \g[3][1] , \g[3][0] , \g[2][63] , \g[2][62] , \g[2][61] ,
         \g[2][60] , \g[2][59] , \g[2][58] , \g[2][57] , \g[2][56] ,
         \g[2][55] , \g[2][54] , \g[2][53] , \g[2][52] , \g[2][51] ,
         \g[2][50] , \g[2][49] , \g[2][48] , \g[2][47] , \g[2][46] ,
         \g[2][45] , \g[2][44] , \g[2][43] , \g[2][42] , \g[2][41] ,
         \g[2][40] , \g[2][39] , \g[2][38] , \g[2][37] , \g[2][36] ,
         \g[2][35] , \g[2][34] , \g[2][33] , \g[2][32] , \g[2][31] ,
         \g[2][30] , \g[2][29] , \g[2][28] , \g[2][27] , \g[2][26] ,
         \g[2][25] , \g[2][24] , \g[2][23] , \g[2][22] , \g[2][21] ,
         \g[2][20] , \g[2][19] , \g[2][18] , \g[2][17] , \g[2][16] ,
         \g[2][15] , \g[2][14] , \g[2][13] , \g[2][12] , \g[2][11] ,
         \g[2][10] , \g[2][9] , \g[2][8] , \g[2][7] , \g[2][6] , \g[2][5] ,
         \g[2][4] , \g[2][3] , \g[2][2] , \g[2][1] , \g[2][0] , \g[1][63] ,
         \g[1][62] , \g[1][61] , \g[1][60] , \g[1][59] , \g[1][58] ,
         \g[1][57] , \g[1][56] , \g[1][55] , \g[1][54] , \g[1][53] ,
         \g[1][52] , \g[1][51] , \g[1][50] , \g[1][49] , \g[1][48] ,
         \g[1][47] , \g[1][46] , \g[1][45] , \g[1][44] , \g[1][43] ,
         \g[1][42] , \g[1][41] , \g[1][40] , \g[1][39] , \g[1][38] ,
         \g[1][37] , \g[1][36] , \g[1][35] , \g[1][34] , \g[1][33] ,
         \g[1][32] , \g[1][31] , \g[1][30] , \g[1][29] , \g[1][28] ,
         \g[1][27] , \g[1][26] , \g[1][25] , \g[1][24] , \g[1][23] ,
         \g[1][22] , \g[1][21] , \g[1][20] , \g[1][19] , \g[1][18] ,
         \g[1][17] , \g[1][16] , \g[1][15] , \g[1][14] , \g[1][13] ,
         \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] ,
         \g[1][6] , \g[1][5] , \g[1][4] , \g[1][3] , \g[1][2] , \g[1][1] ,
         \g[1][0] , \g[0][63] , \g[0][62] , \g[0][61] , \g[0][60] , \g[0][59] ,
         \g[0][58] , \g[0][57] , \g[0][56] , \g[0][55] , \g[0][54] ,
         \g[0][53] , \g[0][52] , \g[0][51] , \g[0][50] , \g[0][49] ,
         \g[0][48] , \g[0][47] , \g[0][46] , \g[0][45] , \g[0][44] ,
         \g[0][43] , \g[0][42] , \g[0][41] , \g[0][40] , \g[0][39] ,
         \g[0][38] , \g[0][37] , \g[0][36] , \g[0][35] , \g[0][34] ,
         \g[0][33] , \g[0][32] , \g[0][31] , \g[0][30] , \g[0][29] ,
         \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] , \g[0][24] ,
         \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , \g[0][19] ,
         \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] ,
         \g[0][13] , \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] ,
         \g[0][7] , \g[0][6] , \g[0][5] , \g[0][4] , \g[0][3] , \g[0][2] ,
         \g[0][1] , \g[0][0] , \g2[27][63] , \g2[27][62] , \g2[27][61] ,
         \g2[27][60] , \g2[27][59] , \g2[27][58] , \g2[27][57] , \g2[27][56] ,
         \g2[27][55] , \g2[27][54] , \g2[27][53] , \g2[27][52] , \g2[27][51] ,
         \g2[27][50] , \g2[27][49] , \g2[27][48] , \g2[27][47] , \g2[27][46] ,
         \g2[27][45] , \g2[27][44] , \g2[27][43] , \g2[27][42] , \g2[27][41] ,
         \g2[27][40] , \g2[27][39] , \g2[27][38] , \g2[27][37] , \g2[27][36] ,
         \g2[27][35] , \g2[27][34] , \g2[27][33] , \g2[27][32] , \g2[27][31] ,
         \g2[27][30] , \g2[27][29] , \g2[27][28] , \g2[27][27] , \g2[27][26] ,
         \g2[27][25] , \g2[27][24] , \g2[27][23] , \g2[27][22] , \g2[27][21] ,
         \g2[27][20] , \g2[27][19] , \g2[27][18] , \g2[27][17] , \g2[27][16] ,
         \g2[27][15] , \g2[27][14] , \g2[27][13] , \g2[27][12] , \g2[27][11] ,
         \g2[27][10] , \g2[27][9] , \g2[27][8] , \g2[27][7] , \g2[27][6] ,
         \g2[27][5] , \g2[27][4] , \g2[27][3] , \g2[27][2] , \g2[27][1] ,
         \g2[26][63] , \g2[26][62] , \g2[26][61] , \g2[26][60] , \g2[26][59] ,
         \g2[26][58] , \g2[26][57] , \g2[26][56] , \g2[26][55] , \g2[26][54] ,
         \g2[26][53] , \g2[26][52] , \g2[26][51] , \g2[26][50] , \g2[26][49] ,
         \g2[26][48] , \g2[26][47] , \g2[26][46] , \g2[26][45] , \g2[26][44] ,
         \g2[26][43] , \g2[26][42] , \g2[26][41] , \g2[26][40] , \g2[26][39] ,
         \g2[26][38] , \g2[26][37] , \g2[26][36] , \g2[26][35] , \g2[26][34] ,
         \g2[26][33] , \g2[26][32] , \g2[26][31] , \g2[26][30] , \g2[26][29] ,
         \g2[26][28] , \g2[26][27] , \g2[26][26] , \g2[26][25] , \g2[26][24] ,
         \g2[26][23] , \g2[26][22] , \g2[26][21] , \g2[26][20] , \g2[26][19] ,
         \g2[26][18] , \g2[26][17] , \g2[26][16] , \g2[26][15] , \g2[26][14] ,
         \g2[26][13] , \g2[26][12] , \g2[26][11] , \g2[26][10] , \g2[26][9] ,
         \g2[26][8] , \g2[26][7] , \g2[26][6] , \g2[26][5] , \g2[26][4] ,
         \g2[26][3] , \g2[26][2] , \g2[26][1] , \g2[25][63] , \g2[25][62] ,
         \g2[25][61] , \g2[25][60] , \g2[25][59] , \g2[25][58] , \g2[25][57] ,
         \g2[25][56] , \g2[25][55] , \g2[25][54] , \g2[25][53] , \g2[25][52] ,
         \g2[25][51] , \g2[25][50] , \g2[25][49] , \g2[25][48] , \g2[25][47] ,
         \g2[25][46] , \g2[25][45] , \g2[25][44] , \g2[25][43] , \g2[25][42] ,
         \g2[25][41] , \g2[25][40] , \g2[25][39] , \g2[25][38] , \g2[25][37] ,
         \g2[25][36] , \g2[25][35] , \g2[25][34] , \g2[25][33] , \g2[25][32] ,
         \g2[25][31] , \g2[25][30] , \g2[25][29] , \g2[25][28] , \g2[25][27] ,
         \g2[25][26] , \g2[25][25] , \g2[25][24] , \g2[25][23] , \g2[25][22] ,
         \g2[25][21] , \g2[25][20] , \g2[25][19] , \g2[25][18] , \g2[25][17] ,
         \g2[25][16] , \g2[25][15] , \g2[25][14] , \g2[25][13] , \g2[25][12] ,
         \g2[25][11] , \g2[25][10] , \g2[25][9] , \g2[25][8] , \g2[25][7] ,
         \g2[25][6] , \g2[25][5] , \g2[25][4] , \g2[25][3] , \g2[25][2] ,
         \g2[25][1] , \g2[24][63] , \g2[24][62] , \g2[24][61] , \g2[24][60] ,
         \g2[24][59] , \g2[24][58] , \g2[24][57] , \g2[24][56] , \g2[24][55] ,
         \g2[24][54] , \g2[24][53] , \g2[24][52] , \g2[24][51] , \g2[24][50] ,
         \g2[24][49] , \g2[24][48] , \g2[24][47] , \g2[24][46] , \g2[24][45] ,
         \g2[24][44] , \g2[24][43] , \g2[24][42] , \g2[24][41] , \g2[24][40] ,
         \g2[24][39] , \g2[24][38] , \g2[24][37] , \g2[24][36] , \g2[24][35] ,
         \g2[24][34] , \g2[24][33] , \g2[24][32] , \g2[24][31] , \g2[24][30] ,
         \g2[24][29] , \g2[24][28] , \g2[24][27] , \g2[24][26] , \g2[24][25] ,
         \g2[24][24] , \g2[24][23] , \g2[24][22] , \g2[24][21] , \g2[24][20] ,
         \g2[24][19] , \g2[24][18] , \g2[24][17] , \g2[24][16] , \g2[24][15] ,
         \g2[24][14] , \g2[24][13] , \g2[24][12] , \g2[24][11] , \g2[24][10] ,
         \g2[24][9] , \g2[24][8] , \g2[24][7] , \g2[24][6] , \g2[24][5] ,
         \g2[24][4] , \g2[24][3] , \g2[24][2] , \g2[24][1] , \g2[23][63] ,
         \g2[23][62] , \g2[23][61] , \g2[23][60] , \g2[23][59] , \g2[23][58] ,
         \g2[23][57] , \g2[23][56] , \g2[23][55] , \g2[23][54] , \g2[23][53] ,
         \g2[23][52] , \g2[23][51] , \g2[23][50] , \g2[23][49] , \g2[23][48] ,
         \g2[23][47] , \g2[23][46] , \g2[23][45] , \g2[23][44] , \g2[23][43] ,
         \g2[23][42] , \g2[23][41] , \g2[23][40] , \g2[23][39] , \g2[23][38] ,
         \g2[23][37] , \g2[23][36] , \g2[23][35] , \g2[23][34] , \g2[23][33] ,
         \g2[23][32] , \g2[23][31] , \g2[23][30] , \g2[23][29] , \g2[23][28] ,
         \g2[23][27] , \g2[23][26] , \g2[23][25] , \g2[23][24] , \g2[23][23] ,
         \g2[23][22] , \g2[23][21] , \g2[23][20] , \g2[23][19] , \g2[23][18] ,
         \g2[23][17] , \g2[23][16] , \g2[23][15] , \g2[23][14] , \g2[23][13] ,
         \g2[23][12] , \g2[23][11] , \g2[23][10] , \g2[23][9] , \g2[23][8] ,
         \g2[23][7] , \g2[23][6] , \g2[23][5] , \g2[23][4] , \g2[23][3] ,
         \g2[23][2] , \g2[23][1] , \g2[22][63] , \g2[22][62] , \g2[22][61] ,
         \g2[22][60] , \g2[22][59] , \g2[22][58] , \g2[22][57] , \g2[22][56] ,
         \g2[22][55] , \g2[22][54] , \g2[22][53] , \g2[22][52] , \g2[22][51] ,
         \g2[22][50] , \g2[22][49] , \g2[22][48] , \g2[22][47] , \g2[22][46] ,
         \g2[22][45] , \g2[22][44] , \g2[22][43] , \g2[22][42] , \g2[22][41] ,
         \g2[22][40] , \g2[22][39] , \g2[22][38] , \g2[22][37] , \g2[22][36] ,
         \g2[22][35] , \g2[22][34] , \g2[22][33] , \g2[22][32] , \g2[22][31] ,
         \g2[22][30] , \g2[22][29] , \g2[22][28] , \g2[22][27] , \g2[22][26] ,
         \g2[22][25] , \g2[22][24] , \g2[22][23] , \g2[22][22] , \g2[22][21] ,
         \g2[22][20] , \g2[22][19] , \g2[22][18] , \g2[22][17] , \g2[22][16] ,
         \g2[22][15] , \g2[22][14] , \g2[22][13] , \g2[22][12] , \g2[22][11] ,
         \g2[22][10] , \g2[22][9] , \g2[22][8] , \g2[22][7] , \g2[22][6] ,
         \g2[22][5] , \g2[22][4] , \g2[22][3] , \g2[22][2] , \g2[22][1] ,
         \g2[21][63] , \g2[21][62] , \g2[21][61] , \g2[21][60] , \g2[21][59] ,
         \g2[21][58] , \g2[21][57] , \g2[21][56] , \g2[21][55] , \g2[21][54] ,
         \g2[21][53] , \g2[21][52] , \g2[21][51] , \g2[21][50] , \g2[21][49] ,
         \g2[21][48] , \g2[21][47] , \g2[21][46] , \g2[21][45] , \g2[21][44] ,
         \g2[21][43] , \g2[21][42] , \g2[21][41] , \g2[21][40] , \g2[21][39] ,
         \g2[21][38] , \g2[21][37] , \g2[21][36] , \g2[21][35] , \g2[21][34] ,
         \g2[21][33] , \g2[21][32] , \g2[21][31] , \g2[21][30] , \g2[21][29] ,
         \g2[21][28] , \g2[21][27] , \g2[21][26] , \g2[21][25] , \g2[21][24] ,
         \g2[21][23] , \g2[21][22] , \g2[21][21] , \g2[21][20] , \g2[21][19] ,
         \g2[21][18] , \g2[21][17] , \g2[21][16] , \g2[21][15] , \g2[21][14] ,
         \g2[21][13] , \g2[21][12] , \g2[21][11] , \g2[21][10] , \g2[21][9] ,
         \g2[21][8] , \g2[21][7] , \g2[21][6] , \g2[21][5] , \g2[21][4] ,
         \g2[21][3] , \g2[21][2] , \g2[21][1] , \g2[20][63] , \g2[20][62] ,
         \g2[20][61] , \g2[20][60] , \g2[20][59] , \g2[20][58] , \g2[20][57] ,
         \g2[20][56] , \g2[20][55] , \g2[20][54] , \g2[20][53] , \g2[20][52] ,
         \g2[20][51] , \g2[20][50] , \g2[20][49] , \g2[20][48] , \g2[20][47] ,
         \g2[20][46] , \g2[20][45] , \g2[20][44] , \g2[20][43] , \g2[20][42] ,
         \g2[20][41] , \g2[20][40] , \g2[20][39] , \g2[20][38] , \g2[20][37] ,
         \g2[20][36] , \g2[20][35] , \g2[20][34] , \g2[20][33] , \g2[20][32] ,
         \g2[20][31] , \g2[20][30] , \g2[20][29] , \g2[20][28] , \g2[20][27] ,
         \g2[20][26] , \g2[20][25] , \g2[20][24] , \g2[20][23] , \g2[20][22] ,
         \g2[20][21] , \g2[20][20] , \g2[20][19] , \g2[20][18] , \g2[20][17] ,
         \g2[20][16] , \g2[20][15] , \g2[20][14] , \g2[20][13] , \g2[20][12] ,
         \g2[20][11] , \g2[20][10] , \g2[20][9] , \g2[20][8] , \g2[20][7] ,
         \g2[20][6] , \g2[20][5] , \g2[20][4] , \g2[20][3] , \g2[20][2] ,
         \g2[20][1] , \g2[19][63] , \g2[19][62] , \g2[19][61] , \g2[19][60] ,
         \g2[19][59] , \g2[19][58] , \g2[19][57] , \g2[19][56] , \g2[19][55] ,
         \g2[19][54] , \g2[19][53] , \g2[19][52] , \g2[19][51] , \g2[19][50] ,
         \g2[19][49] , \g2[19][48] , \g2[19][47] , \g2[19][46] , \g2[19][45] ,
         \g2[19][44] , \g2[19][43] , \g2[19][42] , \g2[19][41] , \g2[19][40] ,
         \g2[19][39] , \g2[19][38] , \g2[19][37] , \g2[19][36] , \g2[19][35] ,
         \g2[19][34] , \g2[19][33] , \g2[19][32] , \g2[19][31] , \g2[19][30] ,
         \g2[19][29] , \g2[19][28] , \g2[19][27] , \g2[19][26] , \g2[19][25] ,
         \g2[19][24] , \g2[19][23] , \g2[19][22] , \g2[19][21] , \g2[19][20] ,
         \g2[19][19] , \g2[19][18] , \g2[19][17] , \g2[19][16] , \g2[19][15] ,
         \g2[19][14] , \g2[19][13] , \g2[19][12] , \g2[19][11] , \g2[19][10] ,
         \g2[19][9] , \g2[19][8] , \g2[19][7] , \g2[19][6] , \g2[19][5] ,
         \g2[19][4] , \g2[19][3] , \g2[19][2] , \g2[19][1] , \g2[18][63] ,
         \g2[18][62] , \g2[18][61] , \g2[18][60] , \g2[18][59] , \g2[18][58] ,
         \g2[18][57] , \g2[18][56] , \g2[18][55] , \g2[18][54] , \g2[18][53] ,
         \g2[18][52] , \g2[18][51] , \g2[18][50] , \g2[18][49] , \g2[18][48] ,
         \g2[18][47] , \g2[18][46] , \g2[18][45] , \g2[18][44] , \g2[18][43] ,
         \g2[18][42] , \g2[18][41] , \g2[18][40] , \g2[18][39] , \g2[18][38] ,
         \g2[18][37] , \g2[18][36] , \g2[18][35] , \g2[18][34] , \g2[18][33] ,
         \g2[18][32] , \g2[18][31] , \g2[18][30] , \g2[18][29] , \g2[18][28] ,
         \g2[18][27] , \g2[18][26] , \g2[18][25] , \g2[18][24] , \g2[18][23] ,
         \g2[18][22] , \g2[18][21] , \g2[18][20] , \g2[18][19] , \g2[18][18] ,
         \g2[18][17] , \g2[18][16] , \g2[18][15] , \g2[18][14] , \g2[18][13] ,
         \g2[18][12] , \g2[18][11] , \g2[18][10] , \g2[18][9] , \g2[18][8] ,
         \g2[18][7] , \g2[18][6] , \g2[18][5] , \g2[18][4] , \g2[18][3] ,
         \g2[18][2] , \g2[18][1] , \g2[17][63] , \g2[17][62] , \g2[17][61] ,
         \g2[17][60] , \g2[17][59] , \g2[17][58] , \g2[17][57] , \g2[17][56] ,
         \g2[17][55] , \g2[17][54] , \g2[17][53] , \g2[17][52] , \g2[17][51] ,
         \g2[17][50] , \g2[17][49] , \g2[17][48] , \g2[17][47] , \g2[17][46] ,
         \g2[17][45] , \g2[17][44] , \g2[17][43] , \g2[17][42] , \g2[17][41] ,
         \g2[17][40] , \g2[17][39] , \g2[17][38] , \g2[17][37] , \g2[17][36] ,
         \g2[17][35] , \g2[17][34] , \g2[17][33] , \g2[17][32] , \g2[17][31] ,
         \g2[17][30] , \g2[17][29] , \g2[17][28] , \g2[17][27] , \g2[17][26] ,
         \g2[17][25] , \g2[17][24] , \g2[17][23] , \g2[17][22] , \g2[17][21] ,
         \g2[17][20] , \g2[17][19] , \g2[17][18] , \g2[17][17] , \g2[17][16] ,
         \g2[17][15] , \g2[17][14] , \g2[17][13] , \g2[17][12] , \g2[17][11] ,
         \g2[17][10] , \g2[17][9] , \g2[17][8] , \g2[17][7] , \g2[17][6] ,
         \g2[17][5] , \g2[17][4] , \g2[17][3] , \g2[17][2] , \g2[17][1] ,
         \g2[16][63] , \g2[16][62] , \g2[16][61] , \g2[16][60] , \g2[16][59] ,
         \g2[16][58] , \g2[16][57] , \g2[16][56] , \g2[16][55] , \g2[16][54] ,
         \g2[16][53] , \g2[16][52] , \g2[16][51] , \g2[16][50] , \g2[16][49] ,
         \g2[16][48] , \g2[16][47] , \g2[16][46] , \g2[16][45] , \g2[16][44] ,
         \g2[16][43] , \g2[16][42] , \g2[16][41] , \g2[16][40] , \g2[16][39] ,
         \g2[16][38] , \g2[16][37] , \g2[16][36] , \g2[16][35] , \g2[16][34] ,
         \g2[16][33] , \g2[16][32] , \g2[16][31] , \g2[16][30] , \g2[16][29] ,
         \g2[16][28] , \g2[16][27] , \g2[16][26] , \g2[16][25] , \g2[16][24] ,
         \g2[16][23] , \g2[16][22] , \g2[16][21] , \g2[16][20] , \g2[16][19] ,
         \g2[16][18] , \g2[16][17] , \g2[16][16] , \g2[16][15] , \g2[16][14] ,
         \g2[16][13] , \g2[16][12] , \g2[16][11] , \g2[16][10] , \g2[16][9] ,
         \g2[16][8] , \g2[16][7] , \g2[16][6] , \g2[16][5] , \g2[16][4] ,
         \g2[16][3] , \g2[16][2] , \g2[16][1] , \g2[15][63] , \g2[15][62] ,
         \g2[15][61] , \g2[15][60] , \g2[15][59] , \g2[15][58] , \g2[15][57] ,
         \g2[15][56] , \g2[15][55] , \g2[15][54] , \g2[15][53] , \g2[15][52] ,
         \g2[15][51] , \g2[15][50] , \g2[15][49] , \g2[15][48] , \g2[15][47] ,
         \g2[15][46] , \g2[15][45] , \g2[15][44] , \g2[15][43] , \g2[15][42] ,
         \g2[15][41] , \g2[15][40] , \g2[15][39] , \g2[15][38] , \g2[15][37] ,
         \g2[15][36] , \g2[15][35] , \g2[15][34] , \g2[15][33] , \g2[15][32] ,
         \g2[15][31] , \g2[15][30] , \g2[15][29] , \g2[15][28] , \g2[15][27] ,
         \g2[15][26] , \g2[15][25] , \g2[15][24] , \g2[15][23] , \g2[15][22] ,
         \g2[15][21] , \g2[15][20] , \g2[15][19] , \g2[15][18] , \g2[15][17] ,
         \g2[15][16] , \g2[15][15] , \g2[15][14] , \g2[15][13] , \g2[15][12] ,
         \g2[15][11] , \g2[15][10] , \g2[15][9] , \g2[15][8] , \g2[15][7] ,
         \g2[15][6] , \g2[15][5] , \g2[15][4] , \g2[15][3] , \g2[15][2] ,
         \g2[15][1] , \g2[14][63] , \g2[14][62] , \g2[14][61] , \g2[14][60] ,
         \g2[14][59] , \g2[14][58] , \g2[14][57] , \g2[14][56] , \g2[14][55] ,
         \g2[14][54] , \g2[14][53] , \g2[14][52] , \g2[14][51] , \g2[14][50] ,
         \g2[14][49] , \g2[14][48] , \g2[14][47] , \g2[14][46] , \g2[14][45] ,
         \g2[14][44] , \g2[14][43] , \g2[14][42] , \g2[14][41] , \g2[14][40] ,
         \g2[14][39] , \g2[14][38] , \g2[14][37] , \g2[14][36] , \g2[14][35] ,
         \g2[14][34] , \g2[14][33] , \g2[14][32] , \g2[14][31] , \g2[14][30] ,
         \g2[14][29] , \g2[14][28] , \g2[14][27] , \g2[14][26] , \g2[14][25] ,
         \g2[14][24] , \g2[14][23] , \g2[14][22] , \g2[14][21] , \g2[14][20] ,
         \g2[14][19] , \g2[14][18] , \g2[14][17] , \g2[14][16] , \g2[14][15] ,
         \g2[14][14] , \g2[14][13] , \g2[14][12] , \g2[14][11] , \g2[14][10] ,
         \g2[14][9] , \g2[14][8] , \g2[14][7] , \g2[14][6] , \g2[14][5] ,
         \g2[14][4] , \g2[14][3] , \g2[14][2] , \g2[14][1] , \g2[13][63] ,
         \g2[13][62] , \g2[13][61] , \g2[13][60] , \g2[13][59] , \g2[13][58] ,
         \g2[13][57] , \g2[13][56] , \g2[13][55] , \g2[13][54] , \g2[13][53] ,
         \g2[13][52] , \g2[13][51] , \g2[13][50] , \g2[13][49] , \g2[13][48] ,
         \g2[13][47] , \g2[13][46] , \g2[13][45] , \g2[13][44] , \g2[13][43] ,
         \g2[13][42] , \g2[13][41] , \g2[13][40] , \g2[13][39] , \g2[13][38] ,
         \g2[13][37] , \g2[13][36] , \g2[13][35] , \g2[13][34] , \g2[13][33] ,
         \g2[13][32] , \g2[13][31] , \g2[13][30] , \g2[13][29] , \g2[13][28] ,
         \g2[13][27] , \g2[13][26] , \g2[13][25] , \g2[13][24] , \g2[13][23] ,
         \g2[13][22] , \g2[13][21] , \g2[13][20] , \g2[13][19] , \g2[13][18] ,
         \g2[13][17] , \g2[13][16] , \g2[13][15] , \g2[13][14] , \g2[13][13] ,
         \g2[13][12] , \g2[13][11] , \g2[13][10] , \g2[13][9] , \g2[13][8] ,
         \g2[13][7] , \g2[13][6] , \g2[13][5] , \g2[13][4] , \g2[13][3] ,
         \g2[13][2] , \g2[13][1] , \g2[13][0] , \g2[12][63] , \g2[12][62] ,
         \g2[12][61] , \g2[12][60] , \g2[12][59] , \g2[12][58] , \g2[12][57] ,
         \g2[12][56] , \g2[12][55] , \g2[12][54] , \g2[12][53] , \g2[12][52] ,
         \g2[12][51] , \g2[12][50] , \g2[12][49] , \g2[12][48] , \g2[12][47] ,
         \g2[12][46] , \g2[12][45] , \g2[12][44] , \g2[12][43] , \g2[12][42] ,
         \g2[12][41] , \g2[12][40] , \g2[12][39] , \g2[12][38] , \g2[12][37] ,
         \g2[12][36] , \g2[12][35] , \g2[12][34] , \g2[12][33] , \g2[12][32] ,
         \g2[12][31] , \g2[12][30] , \g2[12][29] , \g2[12][28] , \g2[12][27] ,
         \g2[12][26] , \g2[12][25] , \g2[12][24] , \g2[12][23] , \g2[12][22] ,
         \g2[12][21] , \g2[12][20] , \g2[12][19] , \g2[12][18] , \g2[12][17] ,
         \g2[12][16] , \g2[12][15] , \g2[12][14] , \g2[12][13] , \g2[12][12] ,
         \g2[12][11] , \g2[12][10] , \g2[12][9] , \g2[12][8] , \g2[12][7] ,
         \g2[12][6] , \g2[12][5] , \g2[12][4] , \g2[12][3] , \g2[12][2] ,
         \g2[12][1] , \g2[12][0] , \g2[11][63] , \g2[11][62] , \g2[11][61] ,
         \g2[11][60] , \g2[11][59] , \g2[11][58] , \g2[11][57] , \g2[11][56] ,
         \g2[11][55] , \g2[11][54] , \g2[11][53] , \g2[11][52] , \g2[11][51] ,
         \g2[11][50] , \g2[11][49] , \g2[11][48] , \g2[11][47] , \g2[11][46] ,
         \g2[11][45] , \g2[11][44] , \g2[11][43] , \g2[11][42] , \g2[11][41] ,
         \g2[11][40] , \g2[11][39] , \g2[11][38] , \g2[11][37] , \g2[11][36] ,
         \g2[11][35] , \g2[11][34] , \g2[11][33] , \g2[11][32] , \g2[11][31] ,
         \g2[11][30] , \g2[11][29] , \g2[11][28] , \g2[11][27] , \g2[11][26] ,
         \g2[11][25] , \g2[11][24] , \g2[11][23] , \g2[11][22] , \g2[11][21] ,
         \g2[11][20] , \g2[11][19] , \g2[11][18] , \g2[11][17] , \g2[11][16] ,
         \g2[11][15] , \g2[11][14] , \g2[11][13] , \g2[11][12] , \g2[11][11] ,
         \g2[11][10] , \g2[11][9] , \g2[11][8] , \g2[11][7] , \g2[11][6] ,
         \g2[11][5] , \g2[11][4] , \g2[11][3] , \g2[11][2] , \g2[11][1] ,
         \g2[11][0] , \g2[10][63] , \g2[10][62] , \g2[10][61] , \g2[10][60] ,
         \g2[10][59] , \g2[10][58] , \g2[10][57] , \g2[10][56] , \g2[10][55] ,
         \g2[10][54] , \g2[10][53] , \g2[10][52] , \g2[10][51] , \g2[10][50] ,
         \g2[10][49] , \g2[10][48] , \g2[10][47] , \g2[10][46] , \g2[10][45] ,
         \g2[10][44] , \g2[10][43] , \g2[10][42] , \g2[10][41] , \g2[10][40] ,
         \g2[10][39] , \g2[10][38] , \g2[10][37] , \g2[10][36] , \g2[10][35] ,
         \g2[10][34] , \g2[10][33] , \g2[10][32] , \g2[10][31] , \g2[10][30] ,
         \g2[10][29] , \g2[10][28] , \g2[10][27] , \g2[10][26] , \g2[10][25] ,
         \g2[10][24] , \g2[10][23] , \g2[10][22] , \g2[10][21] , \g2[10][20] ,
         \g2[10][19] , \g2[10][18] , \g2[10][17] , \g2[10][16] , \g2[10][15] ,
         \g2[10][14] , \g2[10][13] , \g2[10][12] , \g2[10][11] , \g2[10][10] ,
         \g2[10][9] , \g2[10][8] , \g2[10][7] , \g2[10][6] , \g2[10][5] ,
         \g2[10][4] , \g2[10][3] , \g2[10][2] , \g2[10][1] , \g2[10][0] ,
         \g2[9][63] , \g2[9][62] , \g2[9][61] , \g2[9][60] , \g2[9][59] ,
         \g2[9][58] , \g2[9][57] , \g2[9][56] , \g2[9][55] , \g2[9][54] ,
         \g2[9][53] , \g2[9][52] , \g2[9][51] , \g2[9][50] , \g2[9][49] ,
         \g2[9][48] , \g2[9][47] , \g2[9][46] , \g2[9][45] , \g2[9][44] ,
         \g2[9][43] , \g2[9][42] , \g2[9][41] , \g2[9][40] , \g2[9][39] ,
         \g2[9][38] , \g2[9][37] , \g2[9][36] , \g2[9][35] , \g2[9][34] ,
         \g2[9][33] , \g2[9][32] , \g2[9][31] , \g2[9][30] , \g2[9][29] ,
         \g2[9][28] , \g2[9][27] , \g2[9][26] , \g2[9][25] , \g2[9][24] ,
         \g2[9][23] , \g2[9][22] , \g2[9][21] , \g2[9][20] , \g2[9][19] ,
         \g2[9][18] , \g2[9][17] , \g2[9][16] , \g2[9][15] , \g2[9][14] ,
         \g2[9][13] , \g2[9][12] , \g2[9][11] , \g2[9][10] , \g2[9][9] ,
         \g2[9][8] , \g2[9][7] , \g2[9][6] , \g2[9][5] , \g2[9][4] ,
         \g2[9][3] , \g2[9][2] , \g2[9][1] , \g2[9][0] , \g2[8][63] ,
         \g2[8][62] , \g2[8][61] , \g2[8][60] , \g2[8][59] , \g2[8][58] ,
         \g2[8][57] , \g2[8][56] , \g2[8][55] , \g2[8][54] , \g2[8][53] ,
         \g2[8][52] , \g2[8][51] , \g2[8][50] , \g2[8][49] , \g2[8][48] ,
         \g2[8][47] , \g2[8][46] , \g2[8][45] , \g2[8][44] , \g2[8][43] ,
         \g2[8][42] , \g2[8][41] , \g2[8][40] , \g2[8][39] , \g2[8][38] ,
         \g2[8][37] , \g2[8][36] , \g2[8][35] , \g2[8][34] , \g2[8][33] ,
         \g2[8][32] , \g2[8][31] , \g2[8][30] , \g2[8][29] , \g2[8][28] ,
         \g2[8][27] , \g2[8][26] , \g2[8][25] , \g2[8][24] , \g2[8][23] ,
         \g2[8][22] , \g2[8][21] , \g2[8][20] , \g2[8][19] , \g2[8][18] ,
         \g2[8][17] , \g2[8][16] , \g2[8][15] , \g2[8][14] , \g2[8][13] ,
         \g2[8][12] , \g2[8][11] , \g2[8][10] , \g2[8][9] , \g2[8][8] ,
         \g2[8][7] , \g2[8][6] , \g2[8][5] , \g2[8][4] , \g2[8][3] ,
         \g2[8][2] , \g2[8][1] , \g2[8][0] , \g2[7][63] , \g2[7][62] ,
         \g2[7][61] , \g2[7][60] , \g2[7][59] , \g2[7][58] , \g2[7][57] ,
         \g2[7][56] , \g2[7][55] , \g2[7][54] , \g2[7][53] , \g2[7][52] ,
         \g2[7][51] , \g2[7][50] , \g2[7][49] , \g2[7][48] , \g2[7][47] ,
         \g2[7][46] , \g2[7][45] , \g2[7][44] , \g2[7][43] , \g2[7][42] ,
         \g2[7][41] , \g2[7][40] , \g2[7][39] , \g2[7][38] , \g2[7][37] ,
         \g2[7][36] , \g2[7][35] , \g2[7][34] , \g2[7][33] , \g2[7][32] ,
         \g2[7][31] , \g2[7][30] , \g2[7][29] , \g2[7][28] , \g2[7][27] ,
         \g2[7][26] , \g2[7][25] , \g2[7][24] , \g2[7][23] , \g2[7][22] ,
         \g2[7][21] , \g2[7][20] , \g2[7][19] , \g2[7][18] , \g2[7][17] ,
         \g2[7][16] , \g2[7][15] , \g2[7][14] , \g2[7][13] , \g2[7][12] ,
         \g2[7][11] , \g2[7][10] , \g2[7][9] , \g2[7][8] , \g2[7][7] ,
         \g2[7][6] , \g2[7][5] , \g2[7][4] , \g2[7][3] , \g2[7][2] ,
         \g2[7][1] , \g2[7][0] , \g2[6][63] , \g2[6][62] , \g2[6][61] ,
         \g2[6][60] , \g2[6][59] , \g2[6][58] , \g2[6][57] , \g2[6][56] ,
         \g2[6][55] , \g2[6][54] , \g2[6][53] , \g2[6][52] , \g2[6][51] ,
         \g2[6][50] , \g2[6][49] , \g2[6][48] , \g2[6][47] , \g2[6][46] ,
         \g2[6][45] , \g2[6][44] , \g2[6][43] , \g2[6][42] , \g2[6][41] ,
         \g2[6][40] , \g2[6][39] , \g2[6][38] , \g2[6][37] , \g2[6][36] ,
         \g2[6][35] , \g2[6][34] , \g2[6][33] , \g2[6][32] , \g2[6][31] ,
         \g2[6][30] , \g2[6][29] , \g2[6][28] , \g2[6][27] , \g2[6][26] ,
         \g2[6][25] , \g2[6][24] , \g2[6][23] , \g2[6][22] , \g2[6][21] ,
         \g2[6][20] , \g2[6][19] , \g2[6][18] , \g2[6][17] , \g2[6][16] ,
         \g2[6][15] , \g2[6][14] , \g2[6][13] , \g2[6][12] , \g2[6][11] ,
         \g2[6][10] , \g2[6][9] , \g2[6][8] , \g2[6][7] , \g2[6][6] ,
         \g2[6][5] , \g2[6][4] , \g2[6][3] , \g2[6][2] , \g2[6][1] ,
         \g2[6][0] , \g2[5][63] , \g2[5][62] , \g2[5][61] , \g2[5][60] ,
         \g2[5][59] , \g2[5][58] , \g2[5][57] , \g2[5][56] , \g2[5][55] ,
         \g2[5][54] , \g2[5][53] , \g2[5][52] , \g2[5][51] , \g2[5][50] ,
         \g2[5][49] , \g2[5][48] , \g2[5][47] , \g2[5][46] , \g2[5][45] ,
         \g2[5][44] , \g2[5][43] , \g2[5][42] , \g2[5][41] , \g2[5][40] ,
         \g2[5][39] , \g2[5][38] , \g2[5][37] , \g2[5][36] , \g2[5][35] ,
         \g2[5][34] , \g2[5][33] , \g2[5][32] , \g2[5][31] , \g2[5][30] ,
         \g2[5][29] , \g2[5][28] , \g2[5][27] , \g2[5][26] , \g2[5][25] ,
         \g2[5][24] , \g2[5][23] , \g2[5][22] , \g2[5][21] , \g2[5][20] ,
         \g2[5][19] , \g2[5][18] , \g2[5][17] , \g2[5][16] , \g2[5][15] ,
         \g2[5][14] , \g2[5][13] , \g2[5][12] , \g2[5][11] , \g2[5][10] ,
         \g2[5][9] , \g2[5][8] , \g2[5][7] , \g2[5][6] , \g2[5][5] ,
         \g2[5][4] , \g2[5][3] , \g2[5][2] , \g2[5][1] , \g2[5][0] ,
         \g2[4][63] , \g2[4][62] , \g2[4][61] , \g2[4][60] , \g2[4][59] ,
         \g2[4][58] , \g2[4][57] , \g2[4][56] , \g2[4][55] , \g2[4][54] ,
         \g2[4][53] , \g2[4][52] , \g2[4][51] , \g2[4][50] , \g2[4][49] ,
         \g2[4][48] , \g2[4][47] , \g2[4][46] , \g2[4][45] , \g2[4][44] ,
         \g2[4][43] , \g2[4][42] , \g2[4][41] , \g2[4][40] , \g2[4][39] ,
         \g2[4][38] , \g2[4][37] , \g2[4][36] , \g2[4][35] , \g2[4][34] ,
         \g2[4][33] , \g2[4][32] , \g2[4][31] , \g2[4][30] , \g2[4][29] ,
         \g2[4][28] , \g2[4][27] , \g2[4][26] , \g2[4][25] , \g2[4][24] ,
         \g2[4][23] , \g2[4][22] , \g2[4][21] , \g2[4][20] , \g2[4][19] ,
         \g2[4][18] , \g2[4][17] , \g2[4][16] , \g2[4][15] , \g2[4][14] ,
         \g2[4][13] , \g2[4][12] , \g2[4][11] , \g2[4][10] , \g2[4][9] ,
         \g2[4][8] , \g2[4][7] , \g2[4][6] , \g2[4][5] , \g2[4][4] ,
         \g2[4][3] , \g2[4][2] , \g2[4][1] , \g2[4][0] , \g2[3][63] ,
         \g2[3][62] , \g2[3][61] , \g2[3][60] , \g2[3][59] , \g2[3][58] ,
         \g2[3][57] , \g2[3][56] , \g2[3][55] , \g2[3][54] , \g2[3][53] ,
         \g2[3][52] , \g2[3][51] , \g2[3][50] , \g2[3][49] , \g2[3][48] ,
         \g2[3][47] , \g2[3][46] , \g2[3][45] , \g2[3][44] , \g2[3][43] ,
         \g2[3][42] , \g2[3][41] , \g2[3][40] , \g2[3][39] , \g2[3][38] ,
         \g2[3][37] , \g2[3][36] , \g2[3][35] , \g2[3][34] , \g2[3][33] ,
         \g2[3][32] , \g2[3][31] , \g2[3][30] , \g2[3][29] , \g2[3][28] ,
         \g2[3][27] , \g2[3][26] , \g2[3][25] , \g2[3][24] , \g2[3][23] ,
         \g2[3][22] , \g2[3][21] , \g2[3][20] , \g2[3][19] , \g2[3][18] ,
         \g2[3][17] , \g2[3][16] , \g2[3][15] , \g2[3][14] , \g2[3][13] ,
         \g2[3][12] , \g2[3][11] , \g2[3][10] , \g2[3][9] , \g2[3][8] ,
         \g2[3][7] , \g2[3][6] , \g2[3][5] , \g2[3][4] , \g2[3][3] ,
         \g2[3][2] , \g2[3][1] , \g2[3][0] , \g2[2][63] , \g2[2][62] ,
         \g2[2][61] , \g2[2][60] , \g2[2][59] , \g2[2][58] , \g2[2][57] ,
         \g2[2][56] , \g2[2][55] , \g2[2][54] , \g2[2][53] , \g2[2][52] ,
         \g2[2][51] , \g2[2][50] , \g2[2][49] , \g2[2][48] , \g2[2][47] ,
         \g2[2][46] , \g2[2][45] , \g2[2][44] , \g2[2][43] , \g2[2][42] ,
         \g2[2][41] , \g2[2][40] , \g2[2][39] , \g2[2][38] , \g2[2][37] ,
         \g2[2][36] , \g2[2][35] , \g2[2][34] , \g2[2][33] , \g2[2][32] ,
         \g2[2][31] , \g2[2][30] , \g2[2][29] , \g2[2][28] , \g2[2][27] ,
         \g2[2][26] , \g2[2][25] , \g2[2][24] , \g2[2][23] , \g2[2][22] ,
         \g2[2][21] , \g2[2][20] , \g2[2][19] , \g2[2][18] , \g2[2][17] ,
         \g2[2][16] , \g2[2][15] , \g2[2][14] , \g2[2][13] , \g2[2][12] ,
         \g2[2][11] , \g2[2][10] , \g2[2][9] , \g2[2][8] , \g2[2][7] ,
         \g2[2][6] , \g2[2][5] , \g2[2][4] , \g2[2][3] , \g2[2][2] ,
         \g2[2][1] , \g2[2][0] , \g2[1][63] , \g2[1][62] , \g2[1][61] ,
         \g2[1][60] , \g2[1][59] , \g2[1][58] , \g2[1][57] , \g2[1][56] ,
         \g2[1][55] , \g2[1][54] , \g2[1][53] , \g2[1][52] , \g2[1][51] ,
         \g2[1][50] , \g2[1][49] , \g2[1][48] , \g2[1][47] , \g2[1][46] ,
         \g2[1][45] , \g2[1][44] , \g2[1][43] , \g2[1][42] , \g2[1][41] ,
         \g2[1][40] , \g2[1][39] , \g2[1][38] , \g2[1][37] , \g2[1][36] ,
         \g2[1][35] , \g2[1][34] , \g2[1][33] , \g2[1][32] , \g2[1][31] ,
         \g2[1][30] , \g2[1][29] , \g2[1][28] , \g2[1][27] , \g2[1][26] ,
         \g2[1][25] , \g2[1][24] , \g2[1][23] , \g2[1][22] , \g2[1][21] ,
         \g2[1][20] , \g2[1][19] , \g2[1][18] , \g2[1][17] , \g2[1][16] ,
         \g2[1][15] , \g2[1][14] , \g2[1][13] , \g2[1][12] , \g2[1][11] ,
         \g2[1][10] , \g2[1][9] , \g2[1][8] , \g2[1][7] , \g2[1][6] ,
         \g2[1][5] , \g2[1][4] , \g2[1][3] , \g2[1][2] , \g2[1][1] ,
         \g2[1][0] , \g2[0][63] , \g2[0][62] , \g2[0][61] , \g2[0][60] ,
         \g2[0][59] , \g2[0][58] , \g2[0][57] , \g2[0][56] , \g2[0][55] ,
         \g2[0][54] , \g2[0][53] , \g2[0][52] , \g2[0][51] , \g2[0][50] ,
         \g2[0][49] , \g2[0][48] , \g2[0][47] , \g2[0][46] , \g2[0][45] ,
         \g2[0][44] , \g2[0][43] , \g2[0][42] , \g2[0][41] , \g2[0][40] ,
         \g2[0][39] , \g2[0][38] , \g2[0][37] , \g2[0][36] , \g2[0][35] ,
         \g2[0][34] , \g2[0][33] , \g2[0][32] , \g2[0][31] , \g2[0][30] ,
         \g2[0][29] , \g2[0][28] , \g2[0][27] , \g2[0][26] , \g2[0][25] ,
         \g2[0][24] , \g2[0][23] , \g2[0][22] , \g2[0][21] , \g2[0][20] ,
         \g2[0][19] , \g2[0][18] , \g2[0][17] , \g2[0][16] , \g2[0][15] ,
         \g2[0][14] , \g2[0][13] , \g2[0][12] , \g2[0][11] , \g2[0][10] ,
         \g2[0][9] , \g2[0][8] , \g2[0][7] , \g2[0][6] , \g2[0][5] ,
         \g2[0][4] , \g2[0][3] , \g2[0][2] , \g2[0][1] , \g2[0][0] ,
         \g3[17][63] , \g3[17][62] , \g3[17][61] , \g3[17][60] , \g3[17][59] ,
         \g3[17][58] , \g3[17][57] , \g3[17][56] , \g3[17][55] , \g3[17][54] ,
         \g3[17][53] , \g3[17][52] , \g3[17][51] , \g3[17][50] , \g3[17][49] ,
         \g3[17][48] , \g3[17][47] , \g3[17][46] , \g3[17][45] , \g3[17][44] ,
         \g3[17][43] , \g3[17][42] , \g3[17][41] , \g3[17][40] , \g3[17][39] ,
         \g3[17][38] , \g3[17][37] , \g3[17][36] , \g3[17][35] , \g3[17][34] ,
         \g3[17][33] , \g3[17][32] , \g3[17][31] , \g3[17][30] , \g3[17][29] ,
         \g3[17][28] , \g3[17][27] , \g3[17][26] , \g3[17][25] , \g3[17][24] ,
         \g3[17][23] , \g3[17][22] , \g3[17][21] , \g3[17][20] , \g3[17][19] ,
         \g3[17][18] , \g3[17][17] , \g3[17][16] , \g3[17][15] , \g3[17][14] ,
         \g3[17][13] , \g3[17][12] , \g3[17][11] , \g3[17][10] , \g3[17][9] ,
         \g3[17][8] , \g3[17][7] , \g3[17][6] , \g3[17][5] , \g3[17][4] ,
         \g3[17][3] , \g3[17][2] , \g3[17][1] , \g3[16][63] , \g3[16][62] ,
         \g3[16][61] , \g3[16][60] , \g3[16][59] , \g3[16][58] , \g3[16][57] ,
         \g3[16][56] , \g3[16][55] , \g3[16][54] , \g3[16][53] , \g3[16][52] ,
         \g3[16][51] , \g3[16][50] , \g3[16][49] , \g3[16][48] , \g3[16][47] ,
         \g3[16][46] , \g3[16][45] , \g3[16][44] , \g3[16][43] , \g3[16][42] ,
         \g3[16][41] , \g3[16][40] , \g3[16][39] , \g3[16][38] , \g3[16][37] ,
         \g3[16][36] , \g3[16][35] , \g3[16][34] , \g3[16][33] , \g3[16][32] ,
         \g3[16][31] , \g3[16][30] , \g3[16][29] , \g3[16][28] , \g3[16][27] ,
         \g3[16][26] , \g3[16][25] , \g3[16][24] , \g3[16][23] , \g3[16][22] ,
         \g3[16][21] , \g3[16][20] , \g3[16][19] , \g3[16][18] , \g3[16][17] ,
         \g3[16][16] , \g3[16][15] , \g3[16][14] , \g3[16][13] , \g3[16][12] ,
         \g3[16][11] , \g3[16][10] , \g3[16][9] , \g3[16][8] , \g3[16][7] ,
         \g3[16][6] , \g3[16][5] , \g3[16][4] , \g3[16][3] , \g3[16][2] ,
         \g3[16][1] , \g3[15][63] , \g3[15][62] , \g3[15][61] , \g3[15][60] ,
         \g3[15][59] , \g3[15][58] , \g3[15][57] , \g3[15][56] , \g3[15][55] ,
         \g3[15][54] , \g3[15][53] , \g3[15][52] , \g3[15][51] , \g3[15][50] ,
         \g3[15][49] , \g3[15][48] , \g3[15][47] , \g3[15][46] , \g3[15][45] ,
         \g3[15][44] , \g3[15][43] , \g3[15][42] , \g3[15][41] , \g3[15][40] ,
         \g3[15][39] , \g3[15][38] , \g3[15][37] , \g3[15][36] , \g3[15][35] ,
         \g3[15][34] , \g3[15][33] , \g3[15][32] , \g3[15][31] , \g3[15][30] ,
         \g3[15][29] , \g3[15][28] , \g3[15][27] , \g3[15][26] , \g3[15][25] ,
         \g3[15][24] , \g3[15][23] , \g3[15][22] , \g3[15][21] , \g3[15][20] ,
         \g3[15][19] , \g3[15][18] , \g3[15][17] , \g3[15][16] , \g3[15][15] ,
         \g3[15][14] , \g3[15][13] , \g3[15][12] , \g3[15][11] , \g3[15][10] ,
         \g3[15][9] , \g3[15][8] , \g3[15][7] , \g3[15][6] , \g3[15][5] ,
         \g3[15][4] , \g3[15][3] , \g3[15][2] , \g3[15][1] , \g3[14][63] ,
         \g3[14][62] , \g3[14][61] , \g3[14][60] , \g3[14][59] , \g3[14][58] ,
         \g3[14][57] , \g3[14][56] , \g3[14][55] , \g3[14][54] , \g3[14][53] ,
         \g3[14][52] , \g3[14][51] , \g3[14][50] , \g3[14][49] , \g3[14][48] ,
         \g3[14][47] , \g3[14][46] , \g3[14][45] , \g3[14][44] , \g3[14][43] ,
         \g3[14][42] , \g3[14][41] , \g3[14][40] , \g3[14][39] , \g3[14][38] ,
         \g3[14][37] , \g3[14][36] , \g3[14][35] , \g3[14][34] , \g3[14][33] ,
         \g3[14][32] , \g3[14][31] , \g3[14][30] , \g3[14][29] , \g3[14][28] ,
         \g3[14][27] , \g3[14][26] , \g3[14][25] , \g3[14][24] , \g3[14][23] ,
         \g3[14][22] , \g3[14][21] , \g3[14][20] , \g3[14][19] , \g3[14][18] ,
         \g3[14][17] , \g3[14][16] , \g3[14][15] , \g3[14][14] , \g3[14][13] ,
         \g3[14][12] , \g3[14][11] , \g3[14][10] , \g3[14][9] , \g3[14][8] ,
         \g3[14][7] , \g3[14][6] , \g3[14][5] , \g3[14][4] , \g3[14][3] ,
         \g3[14][2] , \g3[14][1] , \g3[13][63] , \g3[13][62] , \g3[13][61] ,
         \g3[13][60] , \g3[13][59] , \g3[13][58] , \g3[13][57] , \g3[13][56] ,
         \g3[13][55] , \g3[13][54] , \g3[13][53] , \g3[13][52] , \g3[13][51] ,
         \g3[13][50] , \g3[13][49] , \g3[13][48] , \g3[13][47] , \g3[13][46] ,
         \g3[13][45] , \g3[13][44] , \g3[13][43] , \g3[13][42] , \g3[13][41] ,
         \g3[13][40] , \g3[13][39] , \g3[13][38] , \g3[13][37] , \g3[13][36] ,
         \g3[13][35] , \g3[13][34] , \g3[13][33] , \g3[13][32] , \g3[13][31] ,
         \g3[13][30] , \g3[13][29] , \g3[13][28] , \g3[13][27] , \g3[13][26] ,
         \g3[13][25] , \g3[13][24] , \g3[13][23] , \g3[13][22] , \g3[13][21] ,
         \g3[13][20] , \g3[13][19] , \g3[13][18] , \g3[13][17] , \g3[13][16] ,
         \g3[13][15] , \g3[13][14] , \g3[13][13] , \g3[13][12] , \g3[13][11] ,
         \g3[13][10] , \g3[13][9] , \g3[13][8] , \g3[13][7] , \g3[13][6] ,
         \g3[13][5] , \g3[13][4] , \g3[13][3] , \g3[13][2] , \g3[13][1] ,
         \g3[12][63] , \g3[12][62] , \g3[12][61] , \g3[12][60] , \g3[12][59] ,
         \g3[12][58] , \g3[12][57] , \g3[12][56] , \g3[12][55] , \g3[12][54] ,
         \g3[12][53] , \g3[12][52] , \g3[12][51] , \g3[12][50] , \g3[12][49] ,
         \g3[12][48] , \g3[12][47] , \g3[12][46] , \g3[12][45] , \g3[12][44] ,
         \g3[12][43] , \g3[12][42] , \g3[12][41] , \g3[12][40] , \g3[12][39] ,
         \g3[12][38] , \g3[12][37] , \g3[12][36] , \g3[12][35] , \g3[12][34] ,
         \g3[12][33] , \g3[12][32] , \g3[12][31] , \g3[12][30] , \g3[12][29] ,
         \g3[12][28] , \g3[12][27] , \g3[12][26] , \g3[12][25] , \g3[12][24] ,
         \g3[12][23] , \g3[12][22] , \g3[12][21] , \g3[12][20] , \g3[12][19] ,
         \g3[12][18] , \g3[12][17] , \g3[12][16] , \g3[12][15] , \g3[12][14] ,
         \g3[12][13] , \g3[12][12] , \g3[12][11] , \g3[12][10] , \g3[12][9] ,
         \g3[12][8] , \g3[12][7] , \g3[12][6] , \g3[12][5] , \g3[12][4] ,
         \g3[12][3] , \g3[12][2] , \g3[12][1] , \g3[11][63] , \g3[11][62] ,
         \g3[11][61] , \g3[11][60] , \g3[11][59] , \g3[11][58] , \g3[11][57] ,
         \g3[11][56] , \g3[11][55] , \g3[11][54] , \g3[11][53] , \g3[11][52] ,
         \g3[11][51] , \g3[11][50] , \g3[11][49] , \g3[11][48] , \g3[11][47] ,
         \g3[11][46] , \g3[11][45] , \g3[11][44] , \g3[11][43] , \g3[11][42] ,
         \g3[11][41] , \g3[11][40] , \g3[11][39] , \g3[11][38] , \g3[11][37] ,
         \g3[11][36] , \g3[11][35] , \g3[11][34] , \g3[11][33] , \g3[11][32] ,
         \g3[11][31] , \g3[11][30] , \g3[11][29] , \g3[11][28] , \g3[11][27] ,
         \g3[11][26] , \g3[11][25] , \g3[11][24] , \g3[11][23] , \g3[11][22] ,
         \g3[11][21] , \g3[11][20] , \g3[11][19] , \g3[11][18] , \g3[11][17] ,
         \g3[11][16] , \g3[11][15] , \g3[11][14] , \g3[11][13] , \g3[11][12] ,
         \g3[11][11] , \g3[11][10] , \g3[11][9] , \g3[11][8] , \g3[11][7] ,
         \g3[11][6] , \g3[11][5] , \g3[11][4] , \g3[11][3] , \g3[11][2] ,
         \g3[11][1] , \g3[10][63] , \g3[10][62] , \g3[10][61] , \g3[10][60] ,
         \g3[10][59] , \g3[10][58] , \g3[10][57] , \g3[10][56] , \g3[10][55] ,
         \g3[10][54] , \g3[10][53] , \g3[10][52] , \g3[10][51] , \g3[10][50] ,
         \g3[10][49] , \g3[10][48] , \g3[10][47] , \g3[10][46] , \g3[10][45] ,
         \g3[10][44] , \g3[10][43] , \g3[10][42] , \g3[10][41] , \g3[10][40] ,
         \g3[10][39] , \g3[10][38] , \g3[10][37] , \g3[10][36] , \g3[10][35] ,
         \g3[10][34] , \g3[10][33] , \g3[10][32] , \g3[10][31] , \g3[10][30] ,
         \g3[10][29] , \g3[10][28] , \g3[10][27] , \g3[10][26] , \g3[10][25] ,
         \g3[10][24] , \g3[10][23] , \g3[10][22] , \g3[10][21] , \g3[10][20] ,
         \g3[10][19] , \g3[10][18] , \g3[10][17] , \g3[10][16] , \g3[10][15] ,
         \g3[10][14] , \g3[10][13] , \g3[10][12] , \g3[10][11] , \g3[10][10] ,
         \g3[10][9] , \g3[10][8] , \g3[10][7] , \g3[10][6] , \g3[10][5] ,
         \g3[10][4] , \g3[10][3] , \g3[10][2] , \g3[10][1] , \g3[9][63] ,
         \g3[9][62] , \g3[9][61] , \g3[9][60] , \g3[9][59] , \g3[9][58] ,
         \g3[9][57] , \g3[9][56] , \g3[9][55] , \g3[9][54] , \g3[9][53] ,
         \g3[9][52] , \g3[9][51] , \g3[9][50] , \g3[9][49] , \g3[9][48] ,
         \g3[9][47] , \g3[9][46] , \g3[9][45] , \g3[9][44] , \g3[9][43] ,
         \g3[9][42] , \g3[9][41] , \g3[9][40] , \g3[9][39] , \g3[9][38] ,
         \g3[9][37] , \g3[9][36] , \g3[9][35] , \g3[9][34] , \g3[9][33] ,
         \g3[9][32] , \g3[9][31] , \g3[9][30] , \g3[9][29] , \g3[9][28] ,
         \g3[9][27] , \g3[9][26] , \g3[9][25] , \g3[9][24] , \g3[9][23] ,
         \g3[9][22] , \g3[9][21] , \g3[9][20] , \g3[9][19] , \g3[9][18] ,
         \g3[9][17] , \g3[9][16] , \g3[9][15] , \g3[9][14] , \g3[9][13] ,
         \g3[9][12] , \g3[9][11] , \g3[9][10] , \g3[9][9] , \g3[9][8] ,
         \g3[9][7] , \g3[9][6] , \g3[9][5] , \g3[9][4] , \g3[9][3] ,
         \g3[9][2] , \g3[9][1] , \g3[8][63] , \g3[8][62] , \g3[8][61] ,
         \g3[8][60] , \g3[8][59] , \g3[8][58] , \g3[8][57] , \g3[8][56] ,
         \g3[8][55] , \g3[8][54] , \g3[8][53] , \g3[8][52] , \g3[8][51] ,
         \g3[8][50] , \g3[8][49] , \g3[8][48] , \g3[8][47] , \g3[8][46] ,
         \g3[8][45] , \g3[8][44] , \g3[8][43] , \g3[8][42] , \g3[8][41] ,
         \g3[8][40] , \g3[8][39] , \g3[8][38] , \g3[8][37] , \g3[8][36] ,
         \g3[8][35] , \g3[8][34] , \g3[8][33] , \g3[8][32] , \g3[8][31] ,
         \g3[8][30] , \g3[8][29] , \g3[8][28] , \g3[8][27] , \g3[8][26] ,
         \g3[8][25] , \g3[8][24] , \g3[8][23] , \g3[8][22] , \g3[8][21] ,
         \g3[8][20] , \g3[8][19] , \g3[8][18] , \g3[8][17] , \g3[8][16] ,
         \g3[8][15] , \g3[8][14] , \g3[8][13] , \g3[8][12] , \g3[8][11] ,
         \g3[8][10] , \g3[8][9] , \g3[8][8] , \g3[8][7] , \g3[8][6] ,
         \g3[8][5] , \g3[8][4] , \g3[8][3] , \g3[8][2] , \g3[8][1] ,
         \g3[8][0] , \g3[7][63] , \g3[7][62] , \g3[7][61] , \g3[7][60] ,
         \g3[7][59] , \g3[7][58] , \g3[7][57] , \g3[7][56] , \g3[7][55] ,
         \g3[7][54] , \g3[7][53] , \g3[7][52] , \g3[7][51] , \g3[7][50] ,
         \g3[7][49] , \g3[7][48] , \g3[7][47] , \g3[7][46] , \g3[7][45] ,
         \g3[7][44] , \g3[7][43] , \g3[7][42] , \g3[7][41] , \g3[7][40] ,
         \g3[7][39] , \g3[7][38] , \g3[7][37] , \g3[7][36] , \g3[7][35] ,
         \g3[7][34] , \g3[7][33] , \g3[7][32] , \g3[7][31] , \g3[7][30] ,
         \g3[7][29] , \g3[7][28] , \g3[7][27] , \g3[7][26] , \g3[7][25] ,
         \g3[7][24] , \g3[7][23] , \g3[7][22] , \g3[7][21] , \g3[7][20] ,
         \g3[7][19] , \g3[7][18] , \g3[7][17] , \g3[7][16] , \g3[7][15] ,
         \g3[7][14] , \g3[7][13] , \g3[7][12] , \g3[7][11] , \g3[7][10] ,
         \g3[7][9] , \g3[7][8] , \g3[7][7] , \g3[7][6] , \g3[7][5] ,
         \g3[7][4] , \g3[7][3] , \g3[7][2] , \g3[7][1] , \g3[7][0] ,
         \g3[6][63] , \g3[6][62] , \g3[6][61] , \g3[6][60] , \g3[6][59] ,
         \g3[6][58] , \g3[6][57] , \g3[6][56] , \g3[6][55] , \g3[6][54] ,
         \g3[6][53] , \g3[6][52] , \g3[6][51] , \g3[6][50] , \g3[6][49] ,
         \g3[6][48] , \g3[6][47] , \g3[6][46] , \g3[6][45] , \g3[6][44] ,
         \g3[6][43] , \g3[6][42] , \g3[6][41] , \g3[6][40] , \g3[6][39] ,
         \g3[6][38] , \g3[6][37] , \g3[6][36] , \g3[6][35] , \g3[6][34] ,
         \g3[6][33] , \g3[6][32] , \g3[6][31] , \g3[6][30] , \g3[6][29] ,
         \g3[6][28] , \g3[6][27] , \g3[6][26] , \g3[6][25] , \g3[6][24] ,
         \g3[6][23] , \g3[6][22] , \g3[6][21] , \g3[6][20] , \g3[6][19] ,
         \g3[6][18] , \g3[6][17] , \g3[6][16] , \g3[6][15] , \g3[6][14] ,
         \g3[6][13] , \g3[6][12] , \g3[6][11] , \g3[6][10] , \g3[6][9] ,
         \g3[6][8] , \g3[6][7] , \g3[6][6] , \g3[6][5] , \g3[6][4] ,
         \g3[6][3] , \g3[6][2] , \g3[6][1] , \g3[6][0] , \g3[5][63] ,
         \g3[5][62] , \g3[5][61] , \g3[5][60] , \g3[5][59] , \g3[5][58] ,
         \g3[5][57] , \g3[5][56] , \g3[5][55] , \g3[5][54] , \g3[5][53] ,
         \g3[5][52] , \g3[5][51] , \g3[5][50] , \g3[5][49] , \g3[5][48] ,
         \g3[5][47] , \g3[5][46] , \g3[5][45] , \g3[5][44] , \g3[5][43] ,
         \g3[5][42] , \g3[5][41] , \g3[5][40] , \g3[5][39] , \g3[5][38] ,
         \g3[5][37] , \g3[5][36] , \g3[5][35] , \g3[5][34] , \g3[5][33] ,
         \g3[5][32] , \g3[5][31] , \g3[5][30] , \g3[5][29] , \g3[5][28] ,
         \g3[5][27] , \g3[5][26] , \g3[5][25] , \g3[5][24] , \g3[5][23] ,
         \g3[5][22] , \g3[5][21] , \g3[5][20] , \g3[5][19] , \g3[5][18] ,
         \g3[5][17] , \g3[5][16] , \g3[5][15] , \g3[5][14] , \g3[5][13] ,
         \g3[5][12] , \g3[5][11] , \g3[5][10] , \g3[5][9] , \g3[5][8] ,
         \g3[5][7] , \g3[5][6] , \g3[5][5] , \g3[5][4] , \g3[5][3] ,
         \g3[5][2] , \g3[5][1] , \g3[5][0] , \g3[4][63] , \g3[4][62] ,
         \g3[4][61] , \g3[4][60] , \g3[4][59] , \g3[4][58] , \g3[4][57] ,
         \g3[4][56] , \g3[4][55] , \g3[4][54] , \g3[4][53] , \g3[4][52] ,
         \g3[4][51] , \g3[4][50] , \g3[4][49] , \g3[4][48] , \g3[4][47] ,
         \g3[4][46] , \g3[4][45] , \g3[4][44] , \g3[4][43] , \g3[4][42] ,
         \g3[4][41] , \g3[4][40] , \g3[4][39] , \g3[4][38] , \g3[4][37] ,
         \g3[4][36] , \g3[4][35] , \g3[4][34] , \g3[4][33] , \g3[4][32] ,
         \g3[4][31] , \g3[4][30] , \g3[4][29] , \g3[4][28] , \g3[4][27] ,
         \g3[4][26] , \g3[4][25] , \g3[4][24] , \g3[4][23] , \g3[4][22] ,
         \g3[4][21] , \g3[4][20] , \g3[4][19] , \g3[4][18] , \g3[4][17] ,
         \g3[4][16] , \g3[4][15] , \g3[4][14] , \g3[4][13] , \g3[4][12] ,
         \g3[4][11] , \g3[4][10] , \g3[4][9] , \g3[4][8] , \g3[4][7] ,
         \g3[4][6] , \g3[4][5] , \g3[4][4] , \g3[4][3] , \g3[4][2] ,
         \g3[4][1] , \g3[4][0] , \g3[3][63] , \g3[3][62] , \g3[3][61] ,
         \g3[3][60] , \g3[3][59] , \g3[3][58] , \g3[3][57] , \g3[3][56] ,
         \g3[3][55] , \g3[3][54] , \g3[3][53] , \g3[3][52] , \g3[3][51] ,
         \g3[3][50] , \g3[3][49] , \g3[3][48] , \g3[3][47] , \g3[3][46] ,
         \g3[3][45] , \g3[3][44] , \g3[3][43] , \g3[3][42] , \g3[3][41] ,
         \g3[3][40] , \g3[3][39] , \g3[3][38] , \g3[3][37] , \g3[3][36] ,
         \g3[3][35] , \g3[3][34] , \g3[3][33] , \g3[3][32] , \g3[3][31] ,
         \g3[3][30] , \g3[3][29] , \g3[3][28] , \g3[3][27] , \g3[3][26] ,
         \g3[3][25] , \g3[3][24] , \g3[3][23] , \g3[3][22] , \g3[3][21] ,
         \g3[3][20] , \g3[3][19] , \g3[3][18] , \g3[3][17] , \g3[3][16] ,
         \g3[3][15] , \g3[3][14] , \g3[3][13] , \g3[3][12] , \g3[3][11] ,
         \g3[3][10] , \g3[3][9] , \g3[3][8] , \g3[3][7] , \g3[3][6] ,
         \g3[3][5] , \g3[3][4] , \g3[3][3] , \g3[3][2] , \g3[3][1] ,
         \g3[3][0] , \g3[2][63] , \g3[2][62] , \g3[2][61] , \g3[2][60] ,
         \g3[2][59] , \g3[2][58] , \g3[2][57] , \g3[2][56] , \g3[2][55] ,
         \g3[2][54] , \g3[2][53] , \g3[2][52] , \g3[2][51] , \g3[2][50] ,
         \g3[2][49] , \g3[2][48] , \g3[2][47] , \g3[2][46] , \g3[2][45] ,
         \g3[2][44] , \g3[2][43] , \g3[2][42] , \g3[2][41] , \g3[2][40] ,
         \g3[2][39] , \g3[2][38] , \g3[2][37] , \g3[2][36] , \g3[2][35] ,
         \g3[2][34] , \g3[2][33] , \g3[2][32] , \g3[2][31] , \g3[2][30] ,
         \g3[2][29] , \g3[2][28] , \g3[2][27] , \g3[2][26] , \g3[2][25] ,
         \g3[2][24] , \g3[2][23] , \g3[2][22] , \g3[2][21] , \g3[2][20] ,
         \g3[2][19] , \g3[2][18] , \g3[2][17] , \g3[2][16] , \g3[2][15] ,
         \g3[2][14] , \g3[2][13] , \g3[2][12] , \g3[2][11] , \g3[2][10] ,
         \g3[2][9] , \g3[2][8] , \g3[2][7] , \g3[2][6] , \g3[2][5] ,
         \g3[2][4] , \g3[2][3] , \g3[2][2] , \g3[2][1] , \g3[2][0] ,
         \g3[1][63] , \g3[1][62] , \g3[1][61] , \g3[1][60] , \g3[1][59] ,
         \g3[1][58] , \g3[1][57] , \g3[1][56] , \g3[1][55] , \g3[1][54] ,
         \g3[1][53] , \g3[1][52] , \g3[1][51] , \g3[1][50] , \g3[1][49] ,
         \g3[1][48] , \g3[1][47] , \g3[1][46] , \g3[1][45] , \g3[1][44] ,
         \g3[1][43] , \g3[1][42] , \g3[1][41] , \g3[1][40] , \g3[1][39] ,
         \g3[1][38] , \g3[1][37] , \g3[1][36] , \g3[1][35] , \g3[1][34] ,
         \g3[1][33] , \g3[1][32] , \g3[1][31] , \g3[1][30] , \g3[1][29] ,
         \g3[1][28] , \g3[1][27] , \g3[1][26] , \g3[1][25] , \g3[1][24] ,
         \g3[1][23] , \g3[1][22] , \g3[1][21] , \g3[1][20] , \g3[1][19] ,
         \g3[1][18] , \g3[1][17] , \g3[1][16] , \g3[1][15] , \g3[1][14] ,
         \g3[1][13] , \g3[1][12] , \g3[1][11] , \g3[1][10] , \g3[1][9] ,
         \g3[1][8] , \g3[1][7] , \g3[1][6] , \g3[1][5] , \g3[1][4] ,
         \g3[1][3] , \g3[1][2] , \g3[1][1] , \g3[1][0] , \g3[0][63] ,
         \g3[0][62] , \g3[0][61] , \g3[0][60] , \g3[0][59] , \g3[0][58] ,
         \g3[0][57] , \g3[0][56] , \g3[0][55] , \g3[0][54] , \g3[0][53] ,
         \g3[0][52] , \g3[0][51] , \g3[0][50] , \g3[0][49] , \g3[0][48] ,
         \g3[0][47] , \g3[0][46] , \g3[0][45] , \g3[0][44] , \g3[0][43] ,
         \g3[0][42] , \g3[0][41] , \g3[0][40] , \g3[0][39] , \g3[0][38] ,
         \g3[0][37] , \g3[0][36] , \g3[0][35] , \g3[0][34] , \g3[0][33] ,
         \g3[0][32] , \g3[0][31] , \g3[0][30] , \g3[0][29] , \g3[0][28] ,
         \g3[0][27] , \g3[0][26] , \g3[0][25] , \g3[0][24] , \g3[0][23] ,
         \g3[0][22] , \g3[0][21] , \g3[0][20] , \g3[0][19] , \g3[0][18] ,
         \g3[0][17] , \g3[0][16] , \g3[0][15] , \g3[0][14] , \g3[0][13] ,
         \g3[0][12] , \g3[0][11] , \g3[0][10] , \g3[0][9] , \g3[0][8] ,
         \g3[0][7] , \g3[0][6] , \g3[0][5] , \g3[0][4] , \g3[0][3] ,
         \g3[0][2] , \g3[0][1] , \g3[0][0] , \g4[11][63] , \g4[11][62] ,
         \g4[11][61] , \g4[11][60] , \g4[11][59] , \g4[11][58] , \g4[11][57] ,
         \g4[11][56] , \g4[11][55] , \g4[11][54] , \g4[11][53] , \g4[11][52] ,
         \g4[11][51] , \g4[11][50] , \g4[11][49] , \g4[11][48] , \g4[11][47] ,
         \g4[11][46] , \g4[11][45] , \g4[11][44] , \g4[11][43] , \g4[11][42] ,
         \g4[11][41] , \g4[11][40] , \g4[11][39] , \g4[11][38] , \g4[11][37] ,
         \g4[11][36] , \g4[11][35] , \g4[11][34] , \g4[11][33] , \g4[11][32] ,
         \g4[11][31] , \g4[11][30] , \g4[11][29] , \g4[11][28] , \g4[11][27] ,
         \g4[11][26] , \g4[11][25] , \g4[11][24] , \g4[11][23] , \g4[11][22] ,
         \g4[11][21] , \g4[11][20] , \g4[11][19] , \g4[11][18] , \g4[11][17] ,
         \g4[11][16] , \g4[11][15] , \g4[11][14] , \g4[11][13] , \g4[11][12] ,
         \g4[11][11] , \g4[11][10] , \g4[11][9] , \g4[11][8] , \g4[11][7] ,
         \g4[11][6] , \g4[11][5] , \g4[11][4] , \g4[11][3] , \g4[11][2] ,
         \g4[11][1] , \g4[10][63] , \g4[10][62] , \g4[10][61] , \g4[10][60] ,
         \g4[10][59] , \g4[10][58] , \g4[10][57] , \g4[10][56] , \g4[10][55] ,
         \g4[10][54] , \g4[10][53] , \g4[10][52] , \g4[10][51] , \g4[10][50] ,
         \g4[10][49] , \g4[10][48] , \g4[10][47] , \g4[10][46] , \g4[10][45] ,
         \g4[10][44] , \g4[10][43] , \g4[10][42] , \g4[10][41] , \g4[10][40] ,
         \g4[10][39] , \g4[10][38] , \g4[10][37] , \g4[10][36] , \g4[10][35] ,
         \g4[10][34] , \g4[10][33] , \g4[10][32] , \g4[10][31] , \g4[10][30] ,
         \g4[10][29] , \g4[10][28] , \g4[10][27] , \g4[10][26] , \g4[10][25] ,
         \g4[10][24] , \g4[10][23] , \g4[10][22] , \g4[10][21] , \g4[10][20] ,
         \g4[10][19] , \g4[10][18] , \g4[10][17] , \g4[10][16] , \g4[10][15] ,
         \g4[10][14] , \g4[10][13] , \g4[10][12] , \g4[10][11] , \g4[10][10] ,
         \g4[10][9] , \g4[10][8] , \g4[10][7] , \g4[10][6] , \g4[10][5] ,
         \g4[10][4] , \g4[10][3] , \g4[10][2] , \g4[10][1] , \g4[9][63] ,
         \g4[9][62] , \g4[9][61] , \g4[9][60] , \g4[9][59] , \g4[9][58] ,
         \g4[9][57] , \g4[9][56] , \g4[9][55] , \g4[9][54] , \g4[9][53] ,
         \g4[9][52] , \g4[9][51] , \g4[9][50] , \g4[9][49] , \g4[9][48] ,
         \g4[9][47] , \g4[9][46] , \g4[9][45] , \g4[9][44] , \g4[9][43] ,
         \g4[9][42] , \g4[9][41] , \g4[9][40] , \g4[9][39] , \g4[9][38] ,
         \g4[9][37] , \g4[9][36] , \g4[9][35] , \g4[9][34] , \g4[9][33] ,
         \g4[9][32] , \g4[9][31] , \g4[9][30] , \g4[9][29] , \g4[9][28] ,
         \g4[9][27] , \g4[9][26] , \g4[9][25] , \g4[9][24] , \g4[9][23] ,
         \g4[9][22] , \g4[9][21] , \g4[9][20] , \g4[9][19] , \g4[9][18] ,
         \g4[9][17] , \g4[9][16] , \g4[9][15] , \g4[9][14] , \g4[9][13] ,
         \g4[9][12] , \g4[9][11] , \g4[9][10] , \g4[9][9] , \g4[9][8] ,
         \g4[9][7] , \g4[9][6] , \g4[9][5] , \g4[9][4] , \g4[9][3] ,
         \g4[9][2] , \g4[9][1] , \g4[8][63] , \g4[8][62] , \g4[8][61] ,
         \g4[8][60] , \g4[8][59] , \g4[8][58] , \g4[8][57] , \g4[8][56] ,
         \g4[8][55] , \g4[8][54] , \g4[8][53] , \g4[8][52] , \g4[8][51] ,
         \g4[8][50] , \g4[8][49] , \g4[8][48] , \g4[8][47] , \g4[8][46] ,
         \g4[8][45] , \g4[8][44] , \g4[8][43] , \g4[8][42] , \g4[8][41] ,
         \g4[8][40] , \g4[8][39] , \g4[8][38] , \g4[8][37] , \g4[8][36] ,
         \g4[8][35] , \g4[8][34] , \g4[8][33] , \g4[8][32] , \g4[8][31] ,
         \g4[8][30] , \g4[8][29] , \g4[8][28] , \g4[8][27] , \g4[8][26] ,
         \g4[8][25] , \g4[8][24] , \g4[8][23] , \g4[8][22] , \g4[8][21] ,
         \g4[8][20] , \g4[8][19] , \g4[8][18] , \g4[8][17] , \g4[8][16] ,
         \g4[8][15] , \g4[8][14] , \g4[8][13] , \g4[8][12] , \g4[8][11] ,
         \g4[8][10] , \g4[8][9] , \g4[8][8] , \g4[8][7] , \g4[8][6] ,
         \g4[8][5] , \g4[8][4] , \g4[8][3] , \g4[8][2] , \g4[8][1] ,
         \g4[7][63] , \g4[7][62] , \g4[7][61] , \g4[7][60] , \g4[7][59] ,
         \g4[7][58] , \g4[7][57] , \g4[7][56] , \g4[7][55] , \g4[7][54] ,
         \g4[7][53] , \g4[7][52] , \g4[7][51] , \g4[7][50] , \g4[7][49] ,
         \g4[7][48] , \g4[7][47] , \g4[7][46] , \g4[7][45] , \g4[7][44] ,
         \g4[7][43] , \g4[7][42] , \g4[7][41] , \g4[7][40] , \g4[7][39] ,
         \g4[7][38] , \g4[7][37] , \g4[7][36] , \g4[7][35] , \g4[7][34] ,
         \g4[7][33] , \g4[7][32] , \g4[7][31] , \g4[7][30] , \g4[7][29] ,
         \g4[7][28] , \g4[7][27] , \g4[7][26] , \g4[7][25] , \g4[7][24] ,
         \g4[7][23] , \g4[7][22] , \g4[7][21] , \g4[7][20] , \g4[7][19] ,
         \g4[7][18] , \g4[7][17] , \g4[7][16] , \g4[7][15] , \g4[7][14] ,
         \g4[7][13] , \g4[7][12] , \g4[7][11] , \g4[7][10] , \g4[7][9] ,
         \g4[7][8] , \g4[7][7] , \g4[7][6] , \g4[7][5] , \g4[7][4] ,
         \g4[7][3] , \g4[7][2] , \g4[7][1] , \g4[6][63] , \g4[6][62] ,
         \g4[6][61] , \g4[6][60] , \g4[6][59] , \g4[6][58] , \g4[6][57] ,
         \g4[6][56] , \g4[6][55] , \g4[6][54] , \g4[6][53] , \g4[6][52] ,
         \g4[6][51] , \g4[6][50] , \g4[6][49] , \g4[6][48] , \g4[6][47] ,
         \g4[6][46] , \g4[6][45] , \g4[6][44] , \g4[6][43] , \g4[6][42] ,
         \g4[6][41] , \g4[6][40] , \g4[6][39] , \g4[6][38] , \g4[6][37] ,
         \g4[6][36] , \g4[6][35] , \g4[6][34] , \g4[6][33] , \g4[6][32] ,
         \g4[6][31] , \g4[6][30] , \g4[6][29] , \g4[6][28] , \g4[6][27] ,
         \g4[6][26] , \g4[6][25] , \g4[6][24] , \g4[6][23] , \g4[6][22] ,
         \g4[6][21] , \g4[6][20] , \g4[6][19] , \g4[6][18] , \g4[6][17] ,
         \g4[6][16] , \g4[6][15] , \g4[6][14] , \g4[6][13] , \g4[6][12] ,
         \g4[6][11] , \g4[6][10] , \g4[6][9] , \g4[6][8] , \g4[6][7] ,
         \g4[6][6] , \g4[6][5] , \g4[6][4] , \g4[6][3] , \g4[6][2] ,
         \g4[6][1] , \g4[5][63] , \g4[5][62] , \g4[5][61] , \g4[5][60] ,
         \g4[5][59] , \g4[5][58] , \g4[5][57] , \g4[5][56] , \g4[5][55] ,
         \g4[5][54] , \g4[5][53] , \g4[5][52] , \g4[5][51] , \g4[5][50] ,
         \g4[5][49] , \g4[5][48] , \g4[5][47] , \g4[5][46] , \g4[5][45] ,
         \g4[5][44] , \g4[5][43] , \g4[5][42] , \g4[5][41] , \g4[5][40] ,
         \g4[5][39] , \g4[5][38] , \g4[5][37] , \g4[5][36] , \g4[5][35] ,
         \g4[5][34] , \g4[5][33] , \g4[5][32] , \g4[5][31] , \g4[5][30] ,
         \g4[5][29] , \g4[5][28] , \g4[5][27] , \g4[5][26] , \g4[5][25] ,
         \g4[5][24] , \g4[5][23] , \g4[5][22] , \g4[5][21] , \g4[5][20] ,
         \g4[5][19] , \g4[5][18] , \g4[5][17] , \g4[5][16] , \g4[5][15] ,
         \g4[5][14] , \g4[5][13] , \g4[5][12] , \g4[5][11] , \g4[5][10] ,
         \g4[5][9] , \g4[5][8] , \g4[5][7] , \g4[5][6] , \g4[5][5] ,
         \g4[5][4] , \g4[5][3] , \g4[5][2] , \g4[5][1] , \g4[5][0] ,
         \g4[4][63] , \g4[4][62] , \g4[4][61] , \g4[4][60] , \g4[4][59] ,
         \g4[4][58] , \g4[4][57] , \g4[4][56] , \g4[4][55] , \g4[4][54] ,
         \g4[4][53] , \g4[4][52] , \g4[4][51] , \g4[4][50] , \g4[4][49] ,
         \g4[4][48] , \g4[4][47] , \g4[4][46] , \g4[4][45] , \g4[4][44] ,
         \g4[4][43] , \g4[4][42] , \g4[4][41] , \g4[4][40] , \g4[4][39] ,
         \g4[4][38] , \g4[4][37] , \g4[4][36] , \g4[4][35] , \g4[4][34] ,
         \g4[4][33] , \g4[4][32] , \g4[4][31] , \g4[4][30] , \g4[4][29] ,
         \g4[4][28] , \g4[4][27] , \g4[4][26] , \g4[4][25] , \g4[4][24] ,
         \g4[4][23] , \g4[4][22] , \g4[4][21] , \g4[4][20] , \g4[4][19] ,
         \g4[4][18] , \g4[4][17] , \g4[4][16] , \g4[4][15] , \g4[4][14] ,
         \g4[4][13] , \g4[4][12] , \g4[4][11] , \g4[4][10] , \g4[4][9] ,
         \g4[4][8] , \g4[4][7] , \g4[4][6] , \g4[4][5] , \g4[4][4] ,
         \g4[4][3] , \g4[4][2] , \g4[4][1] , \g4[4][0] , \g4[3][63] ,
         \g4[3][62] , \g4[3][61] , \g4[3][60] , \g4[3][59] , \g4[3][58] ,
         \g4[3][57] , \g4[3][56] , \g4[3][55] , \g4[3][54] , \g4[3][53] ,
         \g4[3][52] , \g4[3][51] , \g4[3][50] , \g4[3][49] , \g4[3][48] ,
         \g4[3][47] , \g4[3][46] , \g4[3][45] , \g4[3][44] , \g4[3][43] ,
         \g4[3][42] , \g4[3][41] , \g4[3][40] , \g4[3][39] , \g4[3][38] ,
         \g4[3][37] , \g4[3][36] , \g4[3][35] , \g4[3][34] , \g4[3][33] ,
         \g4[3][32] , \g4[3][31] , \g4[3][30] , \g4[3][29] , \g4[3][28] ,
         \g4[3][27] , \g4[3][26] , \g4[3][25] , \g4[3][24] , \g4[3][23] ,
         \g4[3][22] , \g4[3][21] , \g4[3][20] , \g4[3][19] , \g4[3][18] ,
         \g4[3][17] , \g4[3][16] , \g4[3][15] , \g4[3][14] , \g4[3][13] ,
         \g4[3][12] , \g4[3][11] , \g4[3][10] , \g4[3][9] , \g4[3][8] ,
         \g4[3][7] , \g4[3][6] , \g4[3][5] , \g4[3][4] , \g4[3][3] ,
         \g4[3][2] , \g4[3][1] , \g4[3][0] , \g4[2][63] , \g4[2][62] ,
         \g4[2][61] , \g4[2][60] , \g4[2][59] , \g4[2][58] , \g4[2][57] ,
         \g4[2][56] , \g4[2][55] , \g4[2][54] , \g4[2][53] , \g4[2][52] ,
         \g4[2][51] , \g4[2][50] , \g4[2][49] , \g4[2][48] , \g4[2][47] ,
         \g4[2][46] , \g4[2][45] , \g4[2][44] , \g4[2][43] , \g4[2][42] ,
         \g4[2][41] , \g4[2][40] , \g4[2][39] , \g4[2][38] , \g4[2][37] ,
         \g4[2][36] , \g4[2][35] , \g4[2][34] , \g4[2][33] , \g4[2][32] ,
         \g4[2][31] , \g4[2][30] , \g4[2][29] , \g4[2][28] , \g4[2][27] ,
         \g4[2][26] , \g4[2][25] , \g4[2][24] , \g4[2][23] , \g4[2][22] ,
         \g4[2][21] , \g4[2][20] , \g4[2][19] , \g4[2][18] , \g4[2][17] ,
         \g4[2][16] , \g4[2][15] , \g4[2][14] , \g4[2][13] , \g4[2][12] ,
         \g4[2][11] , \g4[2][10] , \g4[2][9] , \g4[2][8] , \g4[2][7] ,
         \g4[2][6] , \g4[2][5] , \g4[2][4] , \g4[2][3] , \g4[2][2] ,
         \g4[2][1] , \g4[2][0] , \g4[1][63] , \g4[1][62] , \g4[1][61] ,
         \g4[1][60] , \g4[1][59] , \g4[1][58] , \g4[1][57] , \g4[1][56] ,
         \g4[1][55] , \g4[1][54] , \g4[1][53] , \g4[1][52] , \g4[1][51] ,
         \g4[1][50] , \g4[1][49] , \g4[1][48] , \g4[1][47] , \g4[1][46] ,
         \g4[1][45] , \g4[1][44] , \g4[1][43] , \g4[1][42] , \g4[1][41] ,
         \g4[1][40] , \g4[1][39] , \g4[1][38] , \g4[1][37] , \g4[1][36] ,
         \g4[1][35] , \g4[1][34] , \g4[1][33] , \g4[1][32] , \g4[1][31] ,
         \g4[1][30] , \g4[1][29] , \g4[1][28] , \g4[1][27] , \g4[1][26] ,
         \g4[1][25] , \g4[1][24] , \g4[1][23] , \g4[1][22] , \g4[1][21] ,
         \g4[1][20] , \g4[1][19] , \g4[1][18] , \g4[1][17] , \g4[1][16] ,
         \g4[1][15] , \g4[1][14] , \g4[1][13] , \g4[1][12] , \g4[1][11] ,
         \g4[1][10] , \g4[1][9] , \g4[1][8] , \g4[1][7] , \g4[1][6] ,
         \g4[1][5] , \g4[1][4] , \g4[1][3] , \g4[1][2] , \g4[1][1] ,
         \g4[1][0] , \g4[0][63] , \g4[0][62] , \g4[0][61] , \g4[0][60] ,
         \g4[0][59] , \g4[0][58] , \g4[0][57] , \g4[0][56] , \g4[0][55] ,
         \g4[0][54] , \g4[0][53] , \g4[0][52] , \g4[0][51] , \g4[0][50] ,
         \g4[0][49] , \g4[0][48] , \g4[0][47] , \g4[0][46] , \g4[0][45] ,
         \g4[0][44] , \g4[0][43] , \g4[0][42] , \g4[0][41] , \g4[0][40] ,
         \g4[0][39] , \g4[0][38] , \g4[0][37] , \g4[0][36] , \g4[0][35] ,
         \g4[0][34] , \g4[0][33] , \g4[0][32] , \g4[0][31] , \g4[0][30] ,
         \g4[0][29] , \g4[0][28] , \g4[0][27] , \g4[0][26] , \g4[0][25] ,
         \g4[0][24] , \g4[0][23] , \g4[0][22] , \g4[0][21] , \g4[0][20] ,
         \g4[0][19] , \g4[0][18] , \g4[0][17] , \g4[0][16] , \g4[0][15] ,
         \g4[0][14] , \g4[0][13] , \g4[0][12] , \g4[0][11] , \g4[0][10] ,
         \g4[0][9] , \g4[0][8] , \g4[0][7] , \g4[0][6] , \g4[0][5] ,
         \g4[0][4] , \g4[0][3] , \g4[0][2] , \g4[0][1] , \g4[0][0] ,
         \g5[7][63] , \g5[7][62] , \g5[7][61] , \g5[7][60] , \g5[7][59] ,
         \g5[7][58] , \g5[7][57] , \g5[7][56] , \g5[7][55] , \g5[7][54] ,
         \g5[7][53] , \g5[7][52] , \g5[7][51] , \g5[7][50] , \g5[7][49] ,
         \g5[7][48] , \g5[7][47] , \g5[7][46] , \g5[7][45] , \g5[7][44] ,
         \g5[7][43] , \g5[7][42] , \g5[7][41] , \g5[7][40] , \g5[7][39] ,
         \g5[7][38] , \g5[7][37] , \g5[7][36] , \g5[7][35] , \g5[7][34] ,
         \g5[7][33] , \g5[7][32] , \g5[7][31] , \g5[7][30] , \g5[7][29] ,
         \g5[7][28] , \g5[7][27] , \g5[7][26] , \g5[7][25] , \g5[7][24] ,
         \g5[7][23] , \g5[7][22] , \g5[7][21] , \g5[7][20] , \g5[7][19] ,
         \g5[7][18] , \g5[7][17] , \g5[7][16] , \g5[7][15] , \g5[7][14] ,
         \g5[7][13] , \g5[7][12] , \g5[7][11] , \g5[7][10] , \g5[7][9] ,
         \g5[7][8] , \g5[7][7] , \g5[7][6] , \g5[7][5] , \g5[7][4] ,
         \g5[7][3] , \g5[7][2] , \g5[7][1] , \g5[6][63] , \g5[6][62] ,
         \g5[6][61] , \g5[6][60] , \g5[6][59] , \g5[6][58] , \g5[6][57] ,
         \g5[6][56] , \g5[6][55] , \g5[6][54] , \g5[6][53] , \g5[6][52] ,
         \g5[6][51] , \g5[6][50] , \g5[6][49] , \g5[6][48] , \g5[6][47] ,
         \g5[6][46] , \g5[6][45] , \g5[6][44] , \g5[6][43] , \g5[6][42] ,
         \g5[6][41] , \g5[6][40] , \g5[6][39] , \g5[6][38] , \g5[6][37] ,
         \g5[6][36] , \g5[6][35] , \g5[6][34] , \g5[6][33] , \g5[6][32] ,
         \g5[6][31] , \g5[6][30] , \g5[6][29] , \g5[6][28] , \g5[6][27] ,
         \g5[6][26] , \g5[6][25] , \g5[6][24] , \g5[6][23] , \g5[6][22] ,
         \g5[6][21] , \g5[6][20] , \g5[6][19] , \g5[6][18] , \g5[6][17] ,
         \g5[6][16] , \g5[6][15] , \g5[6][14] , \g5[6][13] , \g5[6][12] ,
         \g5[6][11] , \g5[6][10] , \g5[6][9] , \g5[6][8] , \g5[6][7] ,
         \g5[6][6] , \g5[6][5] , \g5[6][4] , \g5[6][3] , \g5[6][2] ,
         \g5[6][1] , \g5[5][63] , \g5[5][62] , \g5[5][61] , \g5[5][60] ,
         \g5[5][59] , \g5[5][58] , \g5[5][57] , \g5[5][56] , \g5[5][55] ,
         \g5[5][54] , \g5[5][53] , \g5[5][52] , \g5[5][51] , \g5[5][50] ,
         \g5[5][49] , \g5[5][48] , \g5[5][47] , \g5[5][46] , \g5[5][45] ,
         \g5[5][44] , \g5[5][43] , \g5[5][42] , \g5[5][41] , \g5[5][40] ,
         \g5[5][39] , \g5[5][38] , \g5[5][37] , \g5[5][36] , \g5[5][35] ,
         \g5[5][34] , \g5[5][33] , \g5[5][32] , \g5[5][31] , \g5[5][30] ,
         \g5[5][29] , \g5[5][28] , \g5[5][27] , \g5[5][26] , \g5[5][25] ,
         \g5[5][24] , \g5[5][23] , \g5[5][22] , \g5[5][21] , \g5[5][20] ,
         \g5[5][19] , \g5[5][18] , \g5[5][17] , \g5[5][16] , \g5[5][15] ,
         \g5[5][14] , \g5[5][13] , \g5[5][12] , \g5[5][11] , \g5[5][10] ,
         \g5[5][9] , \g5[5][8] , \g5[5][7] , \g5[5][6] , \g5[5][5] ,
         \g5[5][4] , \g5[5][3] , \g5[5][2] , \g5[5][1] , \g5[4][63] ,
         \g5[4][62] , \g5[4][61] , \g5[4][60] , \g5[4][59] , \g5[4][58] ,
         \g5[4][57] , \g5[4][56] , \g5[4][55] , \g5[4][54] , \g5[4][53] ,
         \g5[4][52] , \g5[4][51] , \g5[4][50] , \g5[4][49] , \g5[4][48] ,
         \g5[4][47] , \g5[4][46] , \g5[4][45] , \g5[4][44] , \g5[4][43] ,
         \g5[4][42] , \g5[4][41] , \g5[4][40] , \g5[4][39] , \g5[4][38] ,
         \g5[4][37] , \g5[4][36] , \g5[4][35] , \g5[4][34] , \g5[4][33] ,
         \g5[4][32] , \g5[4][31] , \g5[4][30] , \g5[4][29] , \g5[4][28] ,
         \g5[4][27] , \g5[4][26] , \g5[4][25] , \g5[4][24] , \g5[4][23] ,
         \g5[4][22] , \g5[4][21] , \g5[4][20] , \g5[4][19] , \g5[4][18] ,
         \g5[4][17] , \g5[4][16] , \g5[4][15] , \g5[4][14] , \g5[4][13] ,
         \g5[4][12] , \g5[4][11] , \g5[4][10] , \g5[4][9] , \g5[4][8] ,
         \g5[4][7] , \g5[4][6] , \g5[4][5] , \g5[4][4] , \g5[4][3] ,
         \g5[4][2] , \g5[4][1] , \g5[3][63] , \g5[3][62] , \g5[3][61] ,
         \g5[3][60] , \g5[3][59] , \g5[3][58] , \g5[3][57] , \g5[3][56] ,
         \g5[3][55] , \g5[3][54] , \g5[3][53] , \g5[3][52] , \g5[3][51] ,
         \g5[3][50] , \g5[3][49] , \g5[3][48] , \g5[3][47] , \g5[3][46] ,
         \g5[3][45] , \g5[3][44] , \g5[3][43] , \g5[3][42] , \g5[3][41] ,
         \g5[3][40] , \g5[3][39] , \g5[3][38] , \g5[3][37] , \g5[3][36] ,
         \g5[3][35] , \g5[3][34] , \g5[3][33] , \g5[3][32] , \g5[3][31] ,
         \g5[3][30] , \g5[3][29] , \g5[3][28] , \g5[3][27] , \g5[3][26] ,
         \g5[3][25] , \g5[3][24] , \g5[3][23] , \g5[3][22] , \g5[3][21] ,
         \g5[3][20] , \g5[3][19] , \g5[3][18] , \g5[3][17] , \g5[3][16] ,
         \g5[3][15] , \g5[3][14] , \g5[3][13] , \g5[3][12] , \g5[3][11] ,
         \g5[3][10] , \g5[3][9] , \g5[3][8] , \g5[3][7] , \g5[3][6] ,
         \g5[3][5] , \g5[3][4] , \g5[3][3] , \g5[3][2] , \g5[3][1] ,
         \g5[3][0] , \g5[2][63] , \g5[2][62] , \g5[2][61] , \g5[2][60] ,
         \g5[2][59] , \g5[2][58] , \g5[2][57] , \g5[2][56] , \g5[2][55] ,
         \g5[2][54] , \g5[2][53] , \g5[2][52] , \g5[2][51] , \g5[2][50] ,
         \g5[2][49] , \g5[2][48] , \g5[2][47] , \g5[2][46] , \g5[2][45] ,
         \g5[2][44] , \g5[2][43] , \g5[2][42] , \g5[2][41] , \g5[2][40] ,
         \g5[2][39] , \g5[2][38] , \g5[2][37] , \g5[2][36] , \g5[2][35] ,
         \g5[2][34] , \g5[2][33] , \g5[2][32] , \g5[2][31] , \g5[2][30] ,
         \g5[2][29] , \g5[2][28] , \g5[2][27] , \g5[2][26] , \g5[2][25] ,
         \g5[2][24] , \g5[2][23] , \g5[2][22] , \g5[2][21] , \g5[2][20] ,
         \g5[2][19] , \g5[2][18] , \g5[2][17] , \g5[2][16] , \g5[2][15] ,
         \g5[2][14] , \g5[2][13] , \g5[2][12] , \g5[2][11] , \g5[2][10] ,
         \g5[2][9] , \g5[2][8] , \g5[2][7] , \g5[2][6] , \g5[2][5] ,
         \g5[2][4] , \g5[2][3] , \g5[2][2] , \g5[2][1] , \g5[2][0] ,
         \g5[1][63] , \g5[1][62] , \g5[1][61] , \g5[1][60] , \g5[1][59] ,
         \g5[1][58] , \g5[1][57] , \g5[1][56] , \g5[1][55] , \g5[1][54] ,
         \g5[1][53] , \g5[1][52] , \g5[1][51] , \g5[1][50] , \g5[1][49] ,
         \g5[1][48] , \g5[1][47] , \g5[1][46] , \g5[1][45] , \g5[1][44] ,
         \g5[1][43] , \g5[1][42] , \g5[1][41] , \g5[1][40] , \g5[1][39] ,
         \g5[1][38] , \g5[1][37] , \g5[1][36] , \g5[1][35] , \g5[1][34] ,
         \g5[1][33] , \g5[1][32] , \g5[1][31] , \g5[1][30] , \g5[1][29] ,
         \g5[1][28] , \g5[1][27] , \g5[1][26] , \g5[1][25] , \g5[1][24] ,
         \g5[1][23] , \g5[1][22] , \g5[1][21] , \g5[1][20] , \g5[1][19] ,
         \g5[1][18] , \g5[1][17] , \g5[1][16] , \g5[1][15] , \g5[1][14] ,
         \g5[1][13] , \g5[1][12] , \g5[1][11] , \g5[1][10] , \g5[1][9] ,
         \g5[1][8] , \g5[1][7] , \g5[1][6] , \g5[1][5] , \g5[1][4] ,
         \g5[1][3] , \g5[1][2] , \g5[1][1] , \g5[1][0] , \g5[0][63] ,
         \g5[0][62] , \g5[0][61] , \g5[0][60] , \g5[0][59] , \g5[0][58] ,
         \g5[0][57] , \g5[0][56] , \g5[0][55] , \g5[0][54] , \g5[0][53] ,
         \g5[0][52] , \g5[0][51] , \g5[0][50] , \g5[0][49] , \g5[0][48] ,
         \g5[0][47] , \g5[0][46] , \g5[0][45] , \g5[0][44] , \g5[0][43] ,
         \g5[0][42] , \g5[0][41] , \g5[0][40] , \g5[0][39] , \g5[0][38] ,
         \g5[0][37] , \g5[0][36] , \g5[0][35] , \g5[0][34] , \g5[0][33] ,
         \g5[0][32] , \g5[0][31] , \g5[0][30] , \g5[0][29] , \g5[0][28] ,
         \g5[0][27] , \g5[0][26] , \g5[0][25] , \g5[0][24] , \g5[0][23] ,
         \g5[0][22] , \g5[0][21] , \g5[0][20] , \g5[0][19] , \g5[0][18] ,
         \g5[0][17] , \g5[0][16] , \g5[0][15] , \g5[0][14] , \g5[0][13] ,
         \g5[0][12] , \g5[0][11] , \g5[0][10] , \g5[0][9] , \g5[0][8] ,
         \g5[0][7] , \g5[0][6] , \g5[0][5] , \g5[0][4] , \g5[0][3] ,
         \g5[0][2] , \g5[0][1] , \g5[0][0] , \g6[5][63] , \g6[5][62] ,
         \g6[5][61] , \g6[5][60] , \g6[5][59] , \g6[5][58] , \g6[5][57] ,
         \g6[5][56] , \g6[5][55] , \g6[5][54] , \g6[5][53] , \g6[5][52] ,
         \g6[5][51] , \g6[5][50] , \g6[5][49] , \g6[5][48] , \g6[5][47] ,
         \g6[5][46] , \g6[5][45] , \g6[5][44] , \g6[5][43] , \g6[5][42] ,
         \g6[5][41] , \g6[5][40] , \g6[5][39] , \g6[5][38] , \g6[5][37] ,
         \g6[5][36] , \g6[5][35] , \g6[5][34] , \g6[5][33] , \g6[5][32] ,
         \g6[5][31] , \g6[5][30] , \g6[5][29] , \g6[5][28] , \g6[5][27] ,
         \g6[5][26] , \g6[5][25] , \g6[5][24] , \g6[5][23] , \g6[5][22] ,
         \g6[5][21] , \g6[5][20] , \g6[5][19] , \g6[5][18] , \g6[5][17] ,
         \g6[5][16] , \g6[5][15] , \g6[5][14] , \g6[5][13] , \g6[5][12] ,
         \g6[5][11] , \g6[5][10] , \g6[5][9] , \g6[5][8] , \g6[5][7] ,
         \g6[5][6] , \g6[5][5] , \g6[5][4] , \g6[5][3] , \g6[5][2] ,
         \g6[5][1] , \g6[4][63] , \g6[4][62] , \g6[4][61] , \g6[4][60] ,
         \g6[4][59] , \g6[4][58] , \g6[4][57] , \g6[4][56] , \g6[4][55] ,
         \g6[4][54] , \g6[4][53] , \g6[4][52] , \g6[4][51] , \g6[4][50] ,
         \g6[4][49] , \g6[4][48] , \g6[4][47] , \g6[4][46] , \g6[4][45] ,
         \g6[4][44] , \g6[4][43] , \g6[4][42] , \g6[4][41] , \g6[4][40] ,
         \g6[4][39] , \g6[4][38] , \g6[4][37] , \g6[4][36] , \g6[4][35] ,
         \g6[4][34] , \g6[4][33] , \g6[4][32] , \g6[4][31] , \g6[4][30] ,
         \g6[4][29] , \g6[4][28] , \g6[4][27] , \g6[4][26] , \g6[4][25] ,
         \g6[4][24] , \g6[4][23] , \g6[4][22] , \g6[4][21] , \g6[4][20] ,
         \g6[4][19] , \g6[4][18] , \g6[4][17] , \g6[4][16] , \g6[4][15] ,
         \g6[4][14] , \g6[4][13] , \g6[4][12] , \g6[4][11] , \g6[4][10] ,
         \g6[4][9] , \g6[4][8] , \g6[4][7] , \g6[4][6] , \g6[4][5] ,
         \g6[4][4] , \g6[4][3] , \g6[4][2] , \g6[4][1] , \g6[4][0] ,
         \g6[3][63] , \g6[3][62] , \g6[3][61] , \g6[3][60] , \g6[3][59] ,
         \g6[3][58] , \g6[3][57] , \g6[3][56] , \g6[3][55] , \g6[3][54] ,
         \g6[3][53] , \g6[3][52] , \g6[3][51] , \g6[3][50] , \g6[3][49] ,
         \g6[3][48] , \g6[3][47] , \g6[3][46] , \g6[3][45] , \g6[3][44] ,
         \g6[3][43] , \g6[3][42] , \g6[3][41] , \g6[3][40] , \g6[3][39] ,
         \g6[3][38] , \g6[3][37] , \g6[3][36] , \g6[3][35] , \g6[3][34] ,
         \g6[3][33] , \g6[3][32] , \g6[3][31] , \g6[3][30] , \g6[3][29] ,
         \g6[3][28] , \g6[3][27] , \g6[3][26] , \g6[3][25] , \g6[3][24] ,
         \g6[3][23] , \g6[3][22] , \g6[3][21] , \g6[3][20] , \g6[3][19] ,
         \g6[3][18] , \g6[3][17] , \g6[3][16] , \g6[3][15] , \g6[3][14] ,
         \g6[3][13] , \g6[3][12] , \g6[3][11] , \g6[3][10] , \g6[3][9] ,
         \g6[3][8] , \g6[3][7] , \g6[3][6] , \g6[3][5] , \g6[3][4] ,
         \g6[3][3] , \g6[3][2] , \g6[3][1] , \g6[2][63] , \g6[2][62] ,
         \g6[2][61] , \g6[2][60] , \g6[2][59] , \g6[2][58] , \g6[2][57] ,
         \g6[2][56] , \g6[2][55] , \g6[2][54] , \g6[2][53] , \g6[2][52] ,
         \g6[2][51] , \g6[2][50] , \g6[2][49] , \g6[2][48] , \g6[2][47] ,
         \g6[2][46] , \g6[2][45] , \g6[2][44] , \g6[2][43] , \g6[2][42] ,
         \g6[2][41] , \g6[2][40] , \g6[2][39] , \g6[2][38] , \g6[2][37] ,
         \g6[2][36] , \g6[2][35] , \g6[2][34] , \g6[2][33] , \g6[2][32] ,
         \g6[2][31] , \g6[2][30] , \g6[2][29] , \g6[2][28] , \g6[2][27] ,
         \g6[2][26] , \g6[2][25] , \g6[2][24] , \g6[2][23] , \g6[2][22] ,
         \g6[2][21] , \g6[2][20] , \g6[2][19] , \g6[2][18] , \g6[2][17] ,
         \g6[2][16] , \g6[2][15] , \g6[2][14] , \g6[2][13] , \g6[2][12] ,
         \g6[2][11] , \g6[2][10] , \g6[2][9] , \g6[2][8] , \g6[2][7] ,
         \g6[2][6] , \g6[2][5] , \g6[2][4] , \g6[2][3] , \g6[2][2] ,
         \g6[2][1] , \g6[2][0] , \g6[1][63] , \g6[1][62] , \g6[1][61] ,
         \g6[1][60] , \g6[1][59] , \g6[1][58] , \g6[1][57] , \g6[1][56] ,
         \g6[1][55] , \g6[1][54] , \g6[1][53] , \g6[1][52] , \g6[1][51] ,
         \g6[1][50] , \g6[1][49] , \g6[1][48] , \g6[1][47] , \g6[1][46] ,
         \g6[1][45] , \g6[1][44] , \g6[1][43] , \g6[1][42] , \g6[1][41] ,
         \g6[1][40] , \g6[1][39] , \g6[1][38] , \g6[1][37] , \g6[1][36] ,
         \g6[1][35] , \g6[1][34] , \g6[1][33] , \g6[1][32] , \g6[1][31] ,
         \g6[1][30] , \g6[1][29] , \g6[1][28] , \g6[1][27] , \g6[1][26] ,
         \g6[1][25] , \g6[1][24] , \g6[1][23] , \g6[1][22] , \g6[1][21] ,
         \g6[1][20] , \g6[1][19] , \g6[1][18] , \g6[1][17] , \g6[1][16] ,
         \g6[1][15] , \g6[1][14] , \g6[1][13] , \g6[1][12] , \g6[1][11] ,
         \g6[1][10] , \g6[1][9] , \g6[1][8] , \g6[1][7] , \g6[1][6] ,
         \g6[1][5] , \g6[1][4] , \g6[1][3] , \g6[1][2] , \g6[1][1] ,
         \g6[0][63] , \g6[0][62] , \g6[0][61] , \g6[0][60] , \g6[0][59] ,
         \g6[0][58] , \g6[0][57] , \g6[0][56] , \g6[0][55] , \g6[0][54] ,
         \g6[0][53] , \g6[0][52] , \g6[0][51] , \g6[0][50] , \g6[0][49] ,
         \g6[0][48] , \g6[0][47] , \g6[0][46] , \g6[0][45] , \g6[0][44] ,
         \g6[0][43] , \g6[0][42] , \g6[0][41] , \g6[0][40] , \g6[0][39] ,
         \g6[0][38] , \g6[0][37] , \g6[0][36] , \g6[0][35] , \g6[0][34] ,
         \g6[0][33] , \g6[0][32] , \g6[0][31] , \g6[0][30] , \g6[0][29] ,
         \g6[0][28] , \g6[0][27] , \g6[0][26] , \g6[0][25] , \g6[0][24] ,
         \g6[0][23] , \g6[0][22] , \g6[0][21] , \g6[0][20] , \g6[0][19] ,
         \g6[0][18] , \g6[0][17] , \g6[0][16] , \g6[0][15] , \g6[0][14] ,
         \g6[0][13] , \g6[0][12] , \g6[0][11] , \g6[0][10] , \g6[0][9] ,
         \g6[0][8] , \g6[0][7] , \g6[0][6] , \g6[0][5] , \g6[0][4] ,
         \g6[0][3] , \g6[0][2] , \g6[0][1] , \g6[0][0] , \g7[3][63] ,
         \g7[3][62] , \g7[3][61] , \g7[3][60] , \g7[3][59] , \g7[3][58] ,
         \g7[3][57] , \g7[3][56] , \g7[3][55] , \g7[3][54] , \g7[3][53] ,
         \g7[3][52] , \g7[3][51] , \g7[3][50] , \g7[3][49] , \g7[3][48] ,
         \g7[3][47] , \g7[3][46] , \g7[3][45] , \g7[3][44] , \g7[3][43] ,
         \g7[3][42] , \g7[3][41] , \g7[3][40] , \g7[3][39] , \g7[3][38] ,
         \g7[3][37] , \g7[3][36] , \g7[3][35] , \g7[3][34] , \g7[3][33] ,
         \g7[3][32] , \g7[3][31] , \g7[3][30] , \g7[3][29] , \g7[3][28] ,
         \g7[3][27] , \g7[3][26] , \g7[3][25] , \g7[3][24] , \g7[3][23] ,
         \g7[3][22] , \g7[3][21] , \g7[3][20] , \g7[3][19] , \g7[3][18] ,
         \g7[3][17] , \g7[3][16] , \g7[3][15] , \g7[3][14] , \g7[3][13] ,
         \g7[3][12] , \g7[3][11] , \g7[3][10] , \g7[3][9] , \g7[3][8] ,
         \g7[3][7] , \g7[3][6] , \g7[3][5] , \g7[3][4] , \g7[3][3] ,
         \g7[3][2] , \g7[3][1] , \g7[2][63] , \g7[2][62] , \g7[2][61] ,
         \g7[2][60] , \g7[2][59] , \g7[2][58] , \g7[2][57] , \g7[2][56] ,
         \g7[2][55] , \g7[2][54] , \g7[2][53] , \g7[2][52] , \g7[2][51] ,
         \g7[2][50] , \g7[2][49] , \g7[2][48] , \g7[2][47] , \g7[2][46] ,
         \g7[2][45] , \g7[2][44] , \g7[2][43] , \g7[2][42] , \g7[2][41] ,
         \g7[2][40] , \g7[2][39] , \g7[2][38] , \g7[2][37] , \g7[2][36] ,
         \g7[2][35] , \g7[2][34] , \g7[2][33] , \g7[2][32] , \g7[2][31] ,
         \g7[2][30] , \g7[2][29] , \g7[2][28] , \g7[2][27] , \g7[2][26] ,
         \g7[2][25] , \g7[2][24] , \g7[2][23] , \g7[2][22] , \g7[2][21] ,
         \g7[2][20] , \g7[2][19] , \g7[2][18] , \g7[2][17] , \g7[2][16] ,
         \g7[2][15] , \g7[2][14] , \g7[2][13] , \g7[2][12] , \g7[2][11] ,
         \g7[2][10] , \g7[2][9] , \g7[2][8] , \g7[2][7] , \g7[2][6] ,
         \g7[2][5] , \g7[2][4] , \g7[2][3] , \g7[2][2] , \g7[2][1] ,
         \g7[2][0] , \g7[1][63] , \g7[1][62] , \g7[1][61] , \g7[1][60] ,
         \g7[1][59] , \g7[1][58] , \g7[1][57] , \g7[1][56] , \g7[1][55] ,
         \g7[1][54] , \g7[1][53] , \g7[1][52] , \g7[1][51] , \g7[1][50] ,
         \g7[1][49] , \g7[1][48] , \g7[1][47] , \g7[1][46] , \g7[1][45] ,
         \g7[1][44] , \g7[1][43] , \g7[1][42] , \g7[1][41] , \g7[1][40] ,
         \g7[1][39] , \g7[1][38] , \g7[1][37] , \g7[1][36] , \g7[1][35] ,
         \g7[1][34] , \g7[1][33] , \g7[1][32] , \g7[1][31] , \g7[1][30] ,
         \g7[1][29] , \g7[1][28] , \g7[1][27] , \g7[1][26] , \g7[1][25] ,
         \g7[1][24] , \g7[1][23] , \g7[1][22] , \g7[1][21] , \g7[1][20] ,
         \g7[1][19] , \g7[1][18] , \g7[1][17] , \g7[1][16] , \g7[1][15] ,
         \g7[1][14] , \g7[1][13] , \g7[1][12] , \g7[1][11] , \g7[1][10] ,
         \g7[1][9] , \g7[1][8] , \g7[1][7] , \g7[1][6] , \g7[1][5] ,
         \g7[1][4] , \g7[1][3] , \g7[1][2] , \g7[1][1] , \g7[0][63] ,
         \g7[0][62] , \g7[0][61] , \g7[0][60] , \g7[0][59] , \g7[0][58] ,
         \g7[0][57] , \g7[0][56] , \g7[0][55] , \g7[0][54] , \g7[0][53] ,
         \g7[0][52] , \g7[0][51] , \g7[0][50] , \g7[0][49] , \g7[0][48] ,
         \g7[0][47] , \g7[0][46] , \g7[0][45] , \g7[0][44] , \g7[0][43] ,
         \g7[0][42] , \g7[0][41] , \g7[0][40] , \g7[0][39] , \g7[0][38] ,
         \g7[0][37] , \g7[0][36] , \g7[0][35] , \g7[0][34] , \g7[0][33] ,
         \g7[0][32] , \g7[0][31] , \g7[0][30] , \g7[0][29] , \g7[0][28] ,
         \g7[0][27] , \g7[0][26] , \g7[0][25] , \g7[0][24] , \g7[0][23] ,
         \g7[0][22] , \g7[0][21] , \g7[0][20] , \g7[0][19] , \g7[0][18] ,
         \g7[0][17] , \g7[0][16] , \g7[0][15] , \g7[0][14] , \g7[0][13] ,
         \g7[0][12] , \g7[0][11] , \g7[0][10] , \g7[0][9] , \g7[0][8] ,
         \g7[0][7] , \g7[0][6] , \g7[0][5] , \g7[0][4] , \g7[0][3] ,
         \g7[0][2] , \g7[0][1] , \g7[0][0] , \g8[1][63] , \g8[1][62] ,
         \g8[1][61] , \g8[1][60] , \g8[1][59] , \g8[1][58] , \g8[1][57] ,
         \g8[1][56] , \g8[1][55] , \g8[1][54] , \g8[1][53] , \g8[1][52] ,
         \g8[1][51] , \g8[1][50] , \g8[1][49] , \g8[1][48] , \g8[1][47] ,
         \g8[1][46] , \g8[1][45] , \g8[1][44] , \g8[1][43] , \g8[1][42] ,
         \g8[1][41] , \g8[1][40] , \g8[1][39] , \g8[1][38] , \g8[1][37] ,
         \g8[1][36] , \g8[1][35] , \g8[1][34] , \g8[1][33] , \g8[1][32] ,
         \g8[1][31] , \g8[1][30] , \g8[1][29] , \g8[1][28] , \g8[1][27] ,
         \g8[1][26] , \g8[1][25] , \g8[1][24] , \g8[1][23] , \g8[1][22] ,
         \g8[1][21] , \g8[1][20] , \g8[1][19] , \g8[1][18] , \g8[1][17] ,
         \g8[1][16] , \g8[1][15] , \g8[1][14] , \g8[1][13] , \g8[1][12] ,
         \g8[1][11] , \g8[1][10] , \g8[1][9] , \g8[1][8] , \g8[1][7] ,
         \g8[1][6] , \g8[1][5] , \g8[1][4] , \g8[1][3] , \g8[1][2] ,
         \g8[1][1] , \g8[0][63] , \g8[0][62] , \g8[0][61] , \g8[0][60] ,
         \g8[0][59] , \g8[0][58] , \g8[0][57] , \g8[0][56] , \g8[0][55] ,
         \g8[0][54] , \g8[0][53] , \g8[0][52] , \g8[0][51] , \g8[0][50] ,
         \g8[0][49] , \g8[0][48] , \g8[0][47] , \g8[0][46] , \g8[0][45] ,
         \g8[0][44] , \g8[0][43] , \g8[0][42] , \g8[0][41] , \g8[0][40] ,
         \g8[0][39] , \g8[0][38] , \g8[0][37] , \g8[0][36] , \g8[0][35] ,
         \g8[0][34] , \g8[0][33] , \g8[0][32] , \g8[0][31] , \g8[0][30] ,
         \g8[0][29] , \g8[0][28] , \g8[0][27] , \g8[0][26] , \g8[0][25] ,
         \g8[0][24] , \g8[0][23] , \g8[0][22] , \g8[0][21] , \g8[0][20] ,
         \g8[0][19] , \g8[0][18] , \g8[0][17] , \g8[0][16] , \g8[0][15] ,
         \g8[0][14] , \g8[0][13] , \g8[0][12] , \g8[0][11] , \g8[0][10] ,
         \g8[0][9] , \g8[0][8] , \g8[0][7] , \g8[0][6] , \g8[0][5] ,
         \g8[0][4] , \g8[0][3] , \g8[0][2] , \g8[0][1] , \g8[0][0] ,
         \g9[1][63] , \g9[1][62] , \g9[1][61] , \g9[1][60] , \g9[1][59] ,
         \g9[1][58] , \g9[1][57] , \g9[1][56] , \g9[1][55] , \g9[1][54] ,
         \g9[1][53] , \g9[1][52] , \g9[1][51] , \g9[1][50] , \g9[1][49] ,
         \g9[1][48] , \g9[1][47] , \g9[1][46] , \g9[1][45] , \g9[1][44] ,
         \g9[1][43] , \g9[1][42] , \g9[1][41] , \g9[1][40] , \g9[1][39] ,
         \g9[1][38] , \g9[1][37] , \g9[1][36] , \g9[1][35] , \g9[1][34] ,
         \g9[1][33] , \g9[1][32] , \g9[1][31] , \g9[1][30] , \g9[1][29] ,
         \g9[1][28] , \g9[1][27] , \g9[1][26] , \g9[1][25] , \g9[1][24] ,
         \g9[1][23] , \g9[1][22] , \g9[1][21] , \g9[1][20] , \g9[1][19] ,
         \g9[1][18] , \g9[1][17] , \g9[1][16] , \g9[1][15] , \g9[1][14] ,
         \g9[1][13] , \g9[1][12] , \g9[1][11] , \g9[1][10] , \g9[1][9] ,
         \g9[1][8] , \g9[1][7] , \g9[1][6] , \g9[1][5] , \g9[1][4] ,
         \g9[1][3] , \g9[1][2] , \g9[1][1] , \g9[0][63] , \g9[0][62] ,
         \g9[0][61] , \g9[0][60] , \g9[0][59] , \g9[0][58] , \g9[0][57] ,
         \g9[0][56] , \g9[0][55] , \g9[0][54] , \g9[0][53] , \g9[0][52] ,
         \g9[0][51] , \g9[0][50] , \g9[0][49] , \g9[0][48] , \g9[0][47] ,
         \g9[0][46] , \g9[0][45] , \g9[0][44] , \g9[0][43] , \g9[0][42] ,
         \g9[0][41] , \g9[0][40] , \g9[0][39] , \g9[0][38] , \g9[0][37] ,
         \g9[0][36] , \g9[0][35] , \g9[0][34] , \g9[0][33] , \g9[0][32] ,
         \g9[0][31] , \g9[0][30] , \g9[0][29] , \g9[0][28] , \g9[0][27] ,
         \g9[0][26] , \g9[0][25] , \g9[0][24] , \g9[0][23] , \g9[0][22] ,
         \g9[0][21] , \g9[0][20] , \g9[0][19] , \g9[0][18] , \g9[0][17] ,
         \g9[0][16] , \g9[0][15] , \g9[0][14] , \g9[0][13] , \g9[0][12] ,
         \g9[0][11] , \g9[0][10] , \g9[0][9] , \g9[0][8] , \g9[0][7] ,
         \g9[0][6] , \g9[0][5] , \g9[0][4] , \g9[0][3] , \g9[0][2] ,
         \g9[0][1] , \g9[0][0] , \g10[1][63] , \g10[1][62] , \g10[1][61] ,
         \g10[1][60] , \g10[1][59] , \g10[1][58] , \g10[1][57] , \g10[1][56] ,
         \g10[1][55] , \g10[1][54] , \g10[1][53] , \g10[1][52] , \g10[1][51] ,
         \g10[1][50] , \g10[1][49] , \g10[1][48] , \g10[1][47] , \g10[1][46] ,
         \g10[1][45] , \g10[1][44] , \g10[1][43] , \g10[1][42] , \g10[1][41] ,
         \g10[1][40] , \g10[1][39] , \g10[1][38] , \g10[1][37] , \g10[1][36] ,
         \g10[1][35] , \g10[1][34] , \g10[1][33] , \g10[1][32] , \g10[1][31] ,
         \g10[1][30] , \g10[1][29] , \g10[1][28] , \g10[1][27] , \g10[1][26] ,
         \g10[1][25] , \g10[1][24] , \g10[1][23] , \g10[1][22] , \g10[1][21] ,
         \g10[1][20] , \g10[1][19] , \g10[1][18] , \g10[1][17] , \g10[1][16] ,
         \g10[1][15] , \g10[1][14] , \g10[1][13] , \g10[1][12] , \g10[1][11] ,
         \g10[1][10] , \g10[1][9] , \g10[1][8] , \g10[1][7] , \g10[1][6] ,
         \g10[1][5] , \g10[1][4] , \g10[1][3] , \g10[1][2] , \g10[1][1] ,
         \g10[0][63] , \g10[0][62] , \g10[0][61] , \g10[0][60] , \g10[0][59] ,
         \g10[0][58] , \g10[0][57] , \g10[0][56] , \g10[0][55] , \g10[0][54] ,
         \g10[0][53] , \g10[0][52] , \g10[0][51] , \g10[0][50] , \g10[0][49] ,
         \g10[0][48] , \g10[0][47] , \g10[0][46] , \g10[0][45] , \g10[0][44] ,
         \g10[0][43] , \g10[0][42] , \g10[0][41] , \g10[0][40] , \g10[0][39] ,
         \g10[0][38] , \g10[0][37] , \g10[0][36] , \g10[0][35] , \g10[0][34] ,
         \g10[0][33] , \g10[0][32] , \g10[0][31] , \g10[0][30] , \g10[0][29] ,
         \g10[0][28] , \g10[0][27] , \g10[0][26] , \g10[0][25] , \g10[0][24] ,
         \g10[0][23] , \g10[0][22] , \g10[0][21] , \g10[0][20] , \g10[0][19] ,
         \g10[0][18] , \g10[0][17] , \g10[0][16] , \g10[0][15] , \g10[0][14] ,
         \g10[0][13] , \g10[0][12] , \g10[0][11] , \g10[0][10] , \g10[0][9] ,
         \g10[0][8] , \g10[0][7] , \g10[0][6] , \g10[0][5] , \g10[0][4] ,
         \g10[0][3] , \g10[0][2] , \g10[0][1] , \g10[0][0] , N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564;
  wire   [31:0] A_reg;
  wire   [31:0] B_reg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61;

  DFFX1 \A_reg_reg[31]  ( .D(N66), .CLK(clk), .Q(A_reg[31]) );
  DFFX1 \A_reg_reg[30]  ( .D(N65), .CLK(clk), .Q(A_reg[30]), .QN(n103) );
  DFFX1 \A_reg_reg[29]  ( .D(N64), .CLK(clk), .Q(A_reg[29]), .QN(n97) );
  DFFX1 \A_reg_reg[28]  ( .D(N63), .CLK(clk), .Q(A_reg[28]), .QN(n92) );
  DFFX1 \A_reg_reg[27]  ( .D(N62), .CLK(clk), .Q(A_reg[27]), .QN(n93) );
  DFFX1 \A_reg_reg[26]  ( .D(N61), .CLK(clk), .Q(A_reg[26]), .QN(n94) );
  DFFX1 \A_reg_reg[25]  ( .D(N60), .CLK(clk), .Q(A_reg[25]), .QN(n95) );
  DFFX1 \A_reg_reg[24]  ( .D(N59), .CLK(clk), .Q(A_reg[24]), .QN(n96) );
  DFFX1 \A_reg_reg[23]  ( .D(N58), .CLK(clk), .Q(A_reg[23]), .QN(n90) );
  DFFX1 \A_reg_reg[22]  ( .D(N57), .CLK(clk), .Q(A_reg[22]), .QN(n73) );
  DFFX1 \A_reg_reg[21]  ( .D(N56), .CLK(clk), .Q(A_reg[21]), .QN(n74) );
  DFFX1 \A_reg_reg[20]  ( .D(N55), .CLK(clk), .Q(A_reg[20]), .QN(n76) );
  DFFX1 \A_reg_reg[19]  ( .D(N54), .CLK(clk), .Q(A_reg[19]), .QN(n75) );
  DFFX1 \A_reg_reg[18]  ( .D(N53), .CLK(clk), .Q(A_reg[18]), .QN(n77) );
  DFFX1 \A_reg_reg[17]  ( .D(N52), .CLK(clk), .Q(A_reg[17]), .QN(n78) );
  DFFX1 \A_reg_reg[16]  ( .D(N51), .CLK(clk), .Q(A_reg[16]), .QN(n80) );
  DFFX1 \A_reg_reg[15]  ( .D(N50), .CLK(clk), .Q(A_reg[15]), .QN(n79) );
  DFFX1 \A_reg_reg[14]  ( .D(N49), .CLK(clk), .Q(A_reg[14]), .QN(n88) );
  DFFX1 \A_reg_reg[13]  ( .D(N48), .CLK(clk), .Q(A_reg[13]), .QN(n89) );
  DFFX1 \A_reg_reg[12]  ( .D(N47), .CLK(clk), .Q(A_reg[12]), .QN(n118) );
  DFFX1 \A_reg_reg[11]  ( .D(N46), .CLK(clk), .Q(A_reg[11]), .QN(n110) );
  DFFX1 \A_reg_reg[9]  ( .D(N44), .CLK(clk), .Q(A_reg[9]), .QN(n119) );
  DFFX1 \A_reg_reg[8]  ( .D(N43), .CLK(clk), .Q(A_reg[8]), .QN(n113) );
  DFFX1 \A_reg_reg[7]  ( .D(N42), .CLK(clk), .Q(A_reg[7]), .QN(n152) );
  DFFX1 \A_reg_reg[6]  ( .D(N41), .CLK(clk), .Q(A_reg[6]), .QN(n148) );
  DFFX1 \A_reg_reg[5]  ( .D(N40), .CLK(clk), .Q(A_reg[5]), .QN(n138) );
  DFFX1 \A_reg_reg[4]  ( .D(N39), .CLK(clk), .Q(A_reg[4]), .QN(n149) );
  DFFX1 \A_reg_reg[3]  ( .D(N38), .CLK(clk), .Q(A_reg[3]), .QN(n146) );
  DFFX1 \A_reg_reg[2]  ( .D(N37), .CLK(clk), .Q(A_reg[2]), .QN(n147) );
  DFFX1 \A_reg_reg[1]  ( .D(N36), .CLK(clk), .Q(A_reg[1]), .QN(n130) );
  DFFX1 \A_reg_reg[0]  ( .D(N35), .CLK(clk), .Q(A_reg[0]), .QN(n120) );
  DFFX1 \B_reg_reg[31]  ( .D(N98), .CLK(clk), .Q(B_reg[31]) );
  DFFX1 \B_reg_reg[30]  ( .D(N97), .CLK(clk), .Q(B_reg[30]), .QN(n104) );
  DFFX1 \B_reg_reg[29]  ( .D(N96), .CLK(clk), .Q(B_reg[29]), .QN(n98) );
  DFFX1 \B_reg_reg[28]  ( .D(N95), .CLK(clk), .Q(B_reg[28]), .QN(n91) );
  DFFX1 \B_reg_reg[27]  ( .D(N94), .CLK(clk), .Q(B_reg[27]), .QN(n99) );
  DFFX1 \B_reg_reg[26]  ( .D(N93), .CLK(clk), .Q(B_reg[26]), .QN(n101) );
  DFFX1 \B_reg_reg[25]  ( .D(N92), .CLK(clk), .Q(B_reg[25]), .QN(n102) );
  DFFX1 \B_reg_reg[24]  ( .D(N91), .CLK(clk), .Q(B_reg[24]), .QN(n100) );
  DFFX1 \B_reg_reg[23]  ( .D(N90), .CLK(clk), .Q(B_reg[23]), .QN(n122) );
  DFFX1 \B_reg_reg[22]  ( .D(N89), .CLK(clk), .Q(B_reg[22]), .QN(n83) );
  DFFX1 \B_reg_reg[21]  ( .D(N88), .CLK(clk), .Q(B_reg[21]), .QN(n84) );
  DFFX1 \B_reg_reg[20]  ( .D(N87), .CLK(clk), .Q(B_reg[20]), .QN(n85) );
  DFFX1 \B_reg_reg[19]  ( .D(N86), .CLK(clk), .Q(B_reg[19]), .QN(n81) );
  DFFX1 \B_reg_reg[18]  ( .D(N85), .CLK(clk), .Q(B_reg[18]), .QN(n86) );
  DFFX1 \B_reg_reg[17]  ( .D(N84), .CLK(clk), .Q(B_reg[17]), .QN(n87) );
  DFFX1 \B_reg_reg[16]  ( .D(N83), .CLK(clk), .Q(B_reg[16]), .QN(n82) );
  DFFX1 \B_reg_reg[15]  ( .D(N82), .CLK(clk), .Q(B_reg[15]), .QN(n107) );
  DFFX1 \B_reg_reg[14]  ( .D(N81), .CLK(clk), .Q(B_reg[14]), .QN(n108) );
  DFFX1 \B_reg_reg[13]  ( .D(N80), .CLK(clk), .Q(B_reg[13]), .QN(n116) );
  DFFX1 \B_reg_reg[12]  ( .D(N79), .CLK(clk), .Q(B_reg[12]), .QN(n111) );
  DFFX1 \B_reg_reg[11]  ( .D(N78), .CLK(clk), .QN(n129) );
  DFFX1 \B_reg_reg[10]  ( .D(N77), .CLK(clk), .Q(B_reg[10]), .QN(n139) );
  DFFX1 \B_reg_reg[9]  ( .D(N76), .CLK(clk), .Q(B_reg[9]), .QN(n123) );
  DFFX1 \B_reg_reg[8]  ( .D(N75), .CLK(clk), .Q(B_reg[8]), .QN(n126) );
  DFFX1 \B_reg_reg[7]  ( .D(N74), .CLK(clk), .Q(B_reg[7]), .QN(n125) );
  DFFX1 \B_reg_reg[6]  ( .D(N73), .CLK(clk), .Q(B_reg[6]), .QN(n133) );
  DFFX1 \B_reg_reg[5]  ( .D(N72), .CLK(clk), .Q(B_reg[5]), .QN(n115) );
  DFFX1 \out_reg[63]  ( .D(N258), .CLK(clk), .Q(out[63]) );
  DFFX1 \out_reg[62]  ( .D(N257), .CLK(clk), .Q(out[62]) );
  DFFX1 \out_reg[61]  ( .D(N256), .CLK(clk), .Q(out[61]) );
  DFFX1 \out_reg[60]  ( .D(N255), .CLK(clk), .Q(out[60]) );
  DFFX1 \out_reg[59]  ( .D(N254), .CLK(clk), .Q(out[59]) );
  DFFX1 \out_reg[58]  ( .D(N253), .CLK(clk), .Q(out[58]) );
  DFFX1 \out_reg[57]  ( .D(N252), .CLK(clk), .Q(out[57]) );
  DFFX1 \out_reg[56]  ( .D(N251), .CLK(clk), .Q(out[56]) );
  DFFX1 \out_reg[55]  ( .D(N250), .CLK(clk), .Q(out[55]) );
  DFFX1 \out_reg[54]  ( .D(N249), .CLK(clk), .Q(out[54]) );
  DFFX1 \out_reg[53]  ( .D(N248), .CLK(clk), .Q(out[53]) );
  DFFX1 \out_reg[52]  ( .D(N247), .CLK(clk), .Q(out[52]) );
  DFFX1 \out_reg[51]  ( .D(N246), .CLK(clk), .Q(out[51]) );
  DFFX1 \out_reg[50]  ( .D(N245), .CLK(clk), .Q(out[50]) );
  DFFX1 \out_reg[49]  ( .D(N244), .CLK(clk), .Q(out[49]) );
  DFFX1 \out_reg[48]  ( .D(N243), .CLK(clk), .Q(out[48]) );
  DFFX1 \out_reg[47]  ( .D(N242), .CLK(clk), .Q(out[47]) );
  DFFX1 \out_reg[46]  ( .D(N241), .CLK(clk), .Q(out[46]) );
  DFFX1 \out_reg[45]  ( .D(N240), .CLK(clk), .Q(out[45]) );
  DFFX1 \out_reg[44]  ( .D(N239), .CLK(clk), .Q(out[44]) );
  DFFX1 \out_reg[43]  ( .D(N238), .CLK(clk), .Q(out[43]) );
  DFFX1 \out_reg[42]  ( .D(N237), .CLK(clk), .Q(out[42]) );
  DFFX1 \out_reg[41]  ( .D(N236), .CLK(clk), .Q(out[41]) );
  DFFX1 \out_reg[40]  ( .D(N235), .CLK(clk), .Q(out[40]) );
  DFFX1 \out_reg[39]  ( .D(N234), .CLK(clk), .Q(out[39]) );
  DFFX1 \out_reg[38]  ( .D(N233), .CLK(clk), .Q(out[38]) );
  DFFX1 \out_reg[37]  ( .D(N232), .CLK(clk), .Q(out[37]) );
  DFFX1 \out_reg[36]  ( .D(N231), .CLK(clk), .Q(out[36]) );
  DFFX1 \out_reg[35]  ( .D(N230), .CLK(clk), .Q(out[35]) );
  DFFX1 \out_reg[34]  ( .D(N229), .CLK(clk), .Q(out[34]) );
  DFFX1 \out_reg[33]  ( .D(N228), .CLK(clk), .Q(out[33]) );
  DFFX1 \out_reg[32]  ( .D(N227), .CLK(clk), .Q(out[32]) );
  DFFX1 \out_reg[31]  ( .D(N226), .CLK(clk), .Q(out[31]) );
  DFFX1 \out_reg[30]  ( .D(N225), .CLK(clk), .Q(out[30]) );
  DFFX1 \out_reg[29]  ( .D(N224), .CLK(clk), .Q(out[29]) );
  DFFX1 \out_reg[28]  ( .D(N223), .CLK(clk), .Q(out[28]) );
  DFFX1 \out_reg[27]  ( .D(N222), .CLK(clk), .Q(out[27]) );
  DFFX1 \out_reg[26]  ( .D(N221), .CLK(clk), .Q(out[26]) );
  DFFX1 \out_reg[25]  ( .D(N220), .CLK(clk), .Q(out[25]) );
  DFFX1 \out_reg[24]  ( .D(N219), .CLK(clk), .Q(out[24]) );
  DFFX1 \out_reg[23]  ( .D(N218), .CLK(clk), .Q(out[23]) );
  DFFX1 \out_reg[22]  ( .D(N217), .CLK(clk), .Q(out[22]) );
  DFFX1 \out_reg[21]  ( .D(N216), .CLK(clk), .Q(out[21]) );
  DFFX1 \out_reg[20]  ( .D(N215), .CLK(clk), .Q(out[20]) );
  DFFX1 \out_reg[19]  ( .D(N214), .CLK(clk), .Q(out[19]) );
  DFFX1 \out_reg[18]  ( .D(N213), .CLK(clk), .Q(out[18]) );
  DFFX1 \out_reg[17]  ( .D(N212), .CLK(clk), .Q(out[17]) );
  DFFX1 \out_reg[16]  ( .D(N211), .CLK(clk), .Q(out[16]) );
  DFFX1 \out_reg[15]  ( .D(N210), .CLK(clk), .Q(out[15]) );
  DFFX1 \out_reg[14]  ( .D(N209), .CLK(clk), .Q(out[14]) );
  DFFX1 \out_reg[13]  ( .D(N208), .CLK(clk), .Q(out[13]) );
  DFFX1 \out_reg[12]  ( .D(N207), .CLK(clk), .Q(out[12]) );
  DFFX1 \out_reg[11]  ( .D(N206), .CLK(clk), .Q(out[11]) );
  DFFX1 \out_reg[10]  ( .D(N205), .CLK(clk), .Q(out[10]) );
  DFFX1 \out_reg[9]  ( .D(N204), .CLK(clk), .Q(out[9]) );
  DFFX1 \out_reg[8]  ( .D(N203), .CLK(clk), .Q(out[8]) );
  DFFX1 \out_reg[7]  ( .D(N202), .CLK(clk), .Q(out[7]) );
  DFFX1 \out_reg[6]  ( .D(N201), .CLK(clk), .Q(out[6]) );
  DFFX1 \out_reg[5]  ( .D(N200), .CLK(clk), .Q(out[5]) );
  DFFX1 \out_reg[4]  ( .D(N199), .CLK(clk), .Q(out[4]) );
  DFFX1 \out_reg[3]  ( .D(N198), .CLK(clk), .Q(out[3]) );
  DFFX1 \out_reg[2]  ( .D(N197), .CLK(clk), .Q(out[2]) );
  DFFX1 \out_reg[1]  ( .D(N196), .CLK(clk), .Q(out[1]) );
  DFFX1 \out_reg[0]  ( .D(N195), .CLK(clk), .Q(out[0]) );
  AND2X1 U1029 ( .IN1(B_reg[8]), .IN2(n545), .Q(\p[8][63] ) );
  AND2X1 U1030 ( .IN1(B_reg[7]), .IN2(n545), .Q(\p[7][63] ) );
  AND2X1 U1031 ( .IN1(B_reg[6]), .IN2(n545), .Q(\p[6][63] ) );
  AND2X1 U1032 ( .IN1(B_reg[5]), .IN2(n545), .Q(\p[5][63] ) );
  AND2X1 U1035 ( .IN1(n542), .IN2(n545), .Q(\p[32][63] ) );
  AND2X1 U1036 ( .IN1(n542), .IN2(A_reg[30]), .Q(\p[33][63] ) );
  AND2X1 U1037 ( .IN1(n542), .IN2(A_reg[29]), .Q(\p[34][63] ) );
  AND2X1 U1038 ( .IN1(n542), .IN2(A_reg[28]), .Q(\p[35][63] ) );
  AND2X1 U1039 ( .IN1(n542), .IN2(A_reg[27]), .Q(\p[36][63] ) );
  AND2X1 U1040 ( .IN1(n542), .IN2(A_reg[26]), .Q(\p[37][63] ) );
  AND2X1 U1041 ( .IN1(n542), .IN2(A_reg[25]), .Q(\p[38][63] ) );
  AND2X1 U1046 ( .IN1(n541), .IN2(A_reg[20]), .Q(\p[43][63] ) );
  AND2X1 U1047 ( .IN1(n541), .IN2(A_reg[19]), .Q(\p[44][63] ) );
  AND2X1 U1048 ( .IN1(n541), .IN2(A_reg[18]), .Q(\p[45][63] ) );
  AND2X1 U1049 ( .IN1(n541), .IN2(A_reg[17]), .Q(\p[46][63] ) );
  AND2X1 U1050 ( .IN1(n541), .IN2(A_reg[16]), .Q(\p[47][63] ) );
  AND2X1 U1051 ( .IN1(n541), .IN2(A_reg[15]), .Q(\p[48][63] ) );
  AND2X1 U1052 ( .IN1(n541), .IN2(A_reg[14]), .Q(\p[49][63] ) );
  AND2X1 U1053 ( .IN1(n541), .IN2(A_reg[13]), .Q(\p[50][63] ) );
  AND2X1 U1054 ( .IN1(n541), .IN2(A_reg[12]), .Q(\p[51][63] ) );
  AND2X1 U1056 ( .IN1(n540), .IN2(A_reg[10]), .Q(\p[53][63] ) );
  AND2X1 U1057 ( .IN1(n540), .IN2(A_reg[9]), .Q(\p[54][63] ) );
  AND2X1 U1058 ( .IN1(n540), .IN2(A_reg[8]), .Q(\p[55][63] ) );
  AND2X1 U1059 ( .IN1(n540), .IN2(A_reg[7]), .Q(\p[56][63] ) );
  AND2X1 U1066 ( .IN1(n540), .IN2(A_reg[0]), .Q(\p[63][63] ) );
  AND2X1 U1067 ( .IN1(B_reg[30]), .IN2(n544), .Q(\p[30][63] ) );
  AND2X1 U1069 ( .IN1(B_reg[29]), .IN2(n544), .Q(\p[29][63] ) );
  AND2X1 U1070 ( .IN1(B_reg[28]), .IN2(n544), .Q(\p[28][63] ) );
  AND2X1 U1071 ( .IN1(B_reg[27]), .IN2(n544), .Q(\p[27][63] ) );
  AND2X1 U1072 ( .IN1(B_reg[26]), .IN2(n544), .Q(\p[26][63] ) );
  AND2X1 U1073 ( .IN1(B_reg[25]), .IN2(n544), .Q(\p[25][63] ) );
  AND2X1 U1078 ( .IN1(B_reg[20]), .IN2(n544), .Q(\p[20][63] ) );
  AND2X1 U1080 ( .IN1(B_reg[19]), .IN2(n543), .Q(\p[19][63] ) );
  AND2X1 U1081 ( .IN1(B_reg[18]), .IN2(n543), .Q(\p[18][63] ) );
  AND2X1 U1082 ( .IN1(B_reg[17]), .IN2(n543), .Q(\p[17][63] ) );
  AND2X1 U1083 ( .IN1(B_reg[16]), .IN2(n543), .Q(\p[16][63] ) );
  AND2X1 U1084 ( .IN1(B_reg[15]), .IN2(n543), .Q(\p[15][63] ) );
  AND2X1 U1085 ( .IN1(B_reg[14]), .IN2(n543), .Q(\p[14][63] ) );
  AND2X1 U1086 ( .IN1(B_reg[13]), .IN2(n543), .Q(\p[13][63] ) );
  AND2X1 U1087 ( .IN1(B_reg[12]), .IN2(n543), .Q(\p[12][63] ) );
  AND2X1 U1088 ( .IN1(n66), .IN2(n543), .Q(\p[11][63] ) );
  AND2X1 U1091 ( .IN1(B[31]), .IN2(n159), .Q(N98) );
  AND2X1 U1092 ( .IN1(B[30]), .IN2(n159), .Q(N97) );
  AND2X1 U1093 ( .IN1(B[29]), .IN2(n159), .Q(N96) );
  AND2X1 U1094 ( .IN1(B[28]), .IN2(n159), .Q(N95) );
  AND2X1 U1095 ( .IN1(B[27]), .IN2(n159), .Q(N94) );
  AND2X1 U1096 ( .IN1(B[26]), .IN2(n159), .Q(N93) );
  AND2X1 U1097 ( .IN1(B[25]), .IN2(n159), .Q(N92) );
  AND2X1 U1098 ( .IN1(B[24]), .IN2(n159), .Q(N91) );
  AND2X1 U1099 ( .IN1(B[23]), .IN2(n159), .Q(N90) );
  AND2X1 U1100 ( .IN1(B[22]), .IN2(n159), .Q(N89) );
  AND2X1 U1101 ( .IN1(B[21]), .IN2(n159), .Q(N88) );
  AND2X1 U1102 ( .IN1(B[20]), .IN2(n159), .Q(N87) );
  AND2X1 U1103 ( .IN1(B[19]), .IN2(n160), .Q(N86) );
  AND2X1 U1104 ( .IN1(B[18]), .IN2(n160), .Q(N85) );
  AND2X1 U1105 ( .IN1(B[17]), .IN2(n160), .Q(N84) );
  AND2X1 U1106 ( .IN1(B[16]), .IN2(n160), .Q(N83) );
  AND2X1 U1107 ( .IN1(B[15]), .IN2(n160), .Q(N82) );
  AND2X1 U1108 ( .IN1(B[14]), .IN2(n160), .Q(N81) );
  AND2X1 U1109 ( .IN1(B[13]), .IN2(n160), .Q(N80) );
  AND2X1 U1110 ( .IN1(B[12]), .IN2(n160), .Q(N79) );
  AND2X1 U1111 ( .IN1(B[11]), .IN2(n160), .Q(N78) );
  AND2X1 U1112 ( .IN1(B[10]), .IN2(n160), .Q(N77) );
  AND2X1 U1113 ( .IN1(B[9]), .IN2(n160), .Q(N76) );
  AND2X1 U1114 ( .IN1(B[8]), .IN2(n160), .Q(N75) );
  AND2X1 U1115 ( .IN1(B[7]), .IN2(n161), .Q(N74) );
  AND2X1 U1116 ( .IN1(B[6]), .IN2(n161), .Q(N73) );
  AND2X1 U1117 ( .IN1(B[5]), .IN2(n161), .Q(N72) );
  AND2X1 U1118 ( .IN1(B[4]), .IN2(n161), .Q(N71) );
  AND2X1 U1119 ( .IN1(B[3]), .IN2(n161), .Q(N70) );
  AND2X1 U1120 ( .IN1(B[2]), .IN2(n161), .Q(N69) );
  AND2X1 U1121 ( .IN1(B[1]), .IN2(n161), .Q(N68) );
  AND2X1 U1122 ( .IN1(B[0]), .IN2(n161), .Q(N67) );
  AND2X1 U1123 ( .IN1(A[31]), .IN2(n161), .Q(N66) );
  AND2X1 U1124 ( .IN1(A[30]), .IN2(n161), .Q(N65) );
  AND2X1 U1125 ( .IN1(A[29]), .IN2(n161), .Q(N64) );
  AND2X1 U1126 ( .IN1(A[28]), .IN2(n161), .Q(N63) );
  AND2X1 U1127 ( .IN1(A[27]), .IN2(n162), .Q(N62) );
  AND2X1 U1128 ( .IN1(A[26]), .IN2(n162), .Q(N61) );
  AND2X1 U1129 ( .IN1(A[25]), .IN2(n162), .Q(N60) );
  AND2X1 U1130 ( .IN1(A[24]), .IN2(n162), .Q(N59) );
  AND2X1 U1131 ( .IN1(A[23]), .IN2(n162), .Q(N58) );
  AND2X1 U1132 ( .IN1(A[22]), .IN2(n162), .Q(N57) );
  AND2X1 U1133 ( .IN1(A[21]), .IN2(n162), .Q(N56) );
  AND2X1 U1134 ( .IN1(A[20]), .IN2(n162), .Q(N55) );
  AND2X1 U1135 ( .IN1(A[19]), .IN2(n162), .Q(N54) );
  AND2X1 U1136 ( .IN1(A[18]), .IN2(n162), .Q(N53) );
  AND2X1 U1137 ( .IN1(A[17]), .IN2(n162), .Q(N52) );
  AND2X1 U1138 ( .IN1(A[16]), .IN2(n162), .Q(N51) );
  AND2X1 U1139 ( .IN1(A[15]), .IN2(n163), .Q(N50) );
  AND2X1 U1140 ( .IN1(A[14]), .IN2(n163), .Q(N49) );
  AND2X1 U1141 ( .IN1(A[13]), .IN2(n163), .Q(N48) );
  AND2X1 U1142 ( .IN1(A[12]), .IN2(n163), .Q(N47) );
  AND2X1 U1143 ( .IN1(A[11]), .IN2(n163), .Q(N46) );
  AND2X1 U1144 ( .IN1(A[10]), .IN2(n163), .Q(N45) );
  AND2X1 U1145 ( .IN1(A[9]), .IN2(n163), .Q(N44) );
  AND2X1 U1146 ( .IN1(A[8]), .IN2(n163), .Q(N43) );
  AND2X1 U1147 ( .IN1(A[7]), .IN2(n163), .Q(N42) );
  AND2X1 U1148 ( .IN1(A[6]), .IN2(n163), .Q(N41) );
  AND2X1 U1149 ( .IN1(A[5]), .IN2(n163), .Q(N40) );
  AND2X1 U1150 ( .IN1(A[4]), .IN2(n163), .Q(N39) );
  AND2X1 U1151 ( .IN1(A[3]), .IN2(n164), .Q(N38) );
  AND2X1 U1152 ( .IN1(A[2]), .IN2(n164), .Q(N37) );
  AND2X1 U1153 ( .IN1(A[1]), .IN2(n164), .Q(N36) );
  AND2X1 U1154 ( .IN1(A[0]), .IN2(n164), .Q(N35) );
  AND2X1 U1155 ( .IN1(N194), .IN2(n164), .Q(N258) );
  AND2X1 U1156 ( .IN1(N193), .IN2(n164), .Q(N257) );
  AND2X1 U1157 ( .IN1(N192), .IN2(n164), .Q(N256) );
  AND2X1 U1158 ( .IN1(N191), .IN2(n164), .Q(N255) );
  AND2X1 U1159 ( .IN1(N190), .IN2(n164), .Q(N254) );
  AND2X1 U1160 ( .IN1(N189), .IN2(n164), .Q(N253) );
  AND2X1 U1161 ( .IN1(N188), .IN2(n164), .Q(N252) );
  AND2X1 U1162 ( .IN1(N187), .IN2(n164), .Q(N251) );
  AND2X1 U1163 ( .IN1(N186), .IN2(n165), .Q(N250) );
  AND2X1 U1164 ( .IN1(N185), .IN2(n165), .Q(N249) );
  AND2X1 U1165 ( .IN1(N184), .IN2(n165), .Q(N248) );
  AND2X1 U1166 ( .IN1(N183), .IN2(n165), .Q(N247) );
  AND2X1 U1167 ( .IN1(N182), .IN2(n165), .Q(N246) );
  AND2X1 U1168 ( .IN1(N181), .IN2(n165), .Q(N245) );
  AND2X1 U1169 ( .IN1(N180), .IN2(n165), .Q(N244) );
  AND2X1 U1170 ( .IN1(N179), .IN2(n165), .Q(N243) );
  AND2X1 U1171 ( .IN1(N178), .IN2(n165), .Q(N242) );
  AND2X1 U1172 ( .IN1(N177), .IN2(n165), .Q(N241) );
  AND2X1 U1173 ( .IN1(N176), .IN2(n165), .Q(N240) );
  AND2X1 U1174 ( .IN1(N175), .IN2(n165), .Q(N239) );
  AND2X1 U1175 ( .IN1(N174), .IN2(n166), .Q(N238) );
  AND2X1 U1176 ( .IN1(N173), .IN2(n166), .Q(N237) );
  AND2X1 U1177 ( .IN1(N172), .IN2(n166), .Q(N236) );
  AND2X1 U1178 ( .IN1(N171), .IN2(n166), .Q(N235) );
  AND2X1 U1179 ( .IN1(N170), .IN2(n166), .Q(N234) );
  AND2X1 U1180 ( .IN1(N169), .IN2(n166), .Q(N233) );
  AND2X1 U1181 ( .IN1(N168), .IN2(n166), .Q(N232) );
  AND2X1 U1182 ( .IN1(N167), .IN2(n166), .Q(N231) );
  AND2X1 U1183 ( .IN1(N166), .IN2(n166), .Q(N230) );
  AND2X1 U1184 ( .IN1(N165), .IN2(n166), .Q(N229) );
  AND2X1 U1185 ( .IN1(N164), .IN2(n166), .Q(N228) );
  AND2X1 U1186 ( .IN1(N163), .IN2(n166), .Q(N227) );
  AND2X1 U1187 ( .IN1(N162), .IN2(n167), .Q(N226) );
  AND2X1 U1188 ( .IN1(N161), .IN2(n167), .Q(N225) );
  AND2X1 U1189 ( .IN1(N160), .IN2(n167), .Q(N224) );
  AND2X1 U1190 ( .IN1(N159), .IN2(n167), .Q(N223) );
  AND2X1 U1191 ( .IN1(N158), .IN2(n167), .Q(N222) );
  AND2X1 U1192 ( .IN1(N157), .IN2(n167), .Q(N221) );
  AND2X1 U1193 ( .IN1(N156), .IN2(n167), .Q(N220) );
  AND2X1 U1194 ( .IN1(N155), .IN2(n167), .Q(N219) );
  AND2X1 U1195 ( .IN1(N154), .IN2(n167), .Q(N218) );
  AND2X1 U1196 ( .IN1(N153), .IN2(n167), .Q(N217) );
  AND2X1 U1197 ( .IN1(N152), .IN2(n167), .Q(N216) );
  AND2X1 U1198 ( .IN1(N151), .IN2(n167), .Q(N215) );
  AND2X1 U1199 ( .IN1(N150), .IN2(n168), .Q(N214) );
  AND2X1 U1200 ( .IN1(N149), .IN2(n168), .Q(N213) );
  AND2X1 U1201 ( .IN1(N148), .IN2(n168), .Q(N212) );
  AND2X1 U1202 ( .IN1(N147), .IN2(n168), .Q(N211) );
  AND2X1 U1203 ( .IN1(N146), .IN2(n168), .Q(N210) );
  AND2X1 U1204 ( .IN1(N145), .IN2(n168), .Q(N209) );
  AND2X1 U1205 ( .IN1(N144), .IN2(n168), .Q(N208) );
  AND2X1 U1206 ( .IN1(N143), .IN2(n168), .Q(N207) );
  AND2X1 U1207 ( .IN1(N142), .IN2(n168), .Q(N206) );
  AND2X1 U1208 ( .IN1(N141), .IN2(n168), .Q(N205) );
  AND2X1 U1209 ( .IN1(N140), .IN2(n168), .Q(N204) );
  AND2X1 U1210 ( .IN1(N139), .IN2(n168), .Q(N203) );
  AND2X1 U1211 ( .IN1(N138), .IN2(n169), .Q(N202) );
  AND2X1 U1212 ( .IN1(N137), .IN2(n169), .Q(N201) );
  AND2X1 U1213 ( .IN1(N136), .IN2(n169), .Q(N200) );
  AND2X1 U1214 ( .IN1(N135), .IN2(n169), .Q(N199) );
  AND2X1 U1215 ( .IN1(N134), .IN2(n169), .Q(N198) );
  AND2X1 U1216 ( .IN1(N133), .IN2(n169), .Q(N197) );
  AND2X1 U1217 ( .IN1(N132), .IN2(n169), .Q(N196) );
  AND2X1 U1218 ( .IN1(N131), .IN2(n169), .Q(N195) );
  FullAdder_0 \level1[0].x6  ( .a({n508, n508, n508, n507, n507, n507, n507, 
        n507, n507, n506, n506, n506, n506, n506, n506, n505, n505, n505, n505, 
        n505, n505, n504, n504, n504, n504, n504, n504, n503, n503, n503, n503, 
        n503, n503, \p[0][30] , \p[0][29] , \p[0][28] , \p[0][27] , \p[0][26] , 
        \p[0][25] , \p[0][24] , \p[0][23] , \p[0][22] , \p[0][21] , \p[0][20] , 
        \p[0][19] , \p[0][18] , \p[0][17] , \p[0][16] , \p[0][15] , \p[0][14] , 
        \p[0][13] , \p[0][12] , \p[0][11] , \p[0][10] , \p[0][9] , \p[0][8] , 
        \p[0][7] , \p[0][6] , \p[0][5] , \p[0][4] , \p[0][3] , \p[0][2] , 
        \p[0][1] , \p[0][0] }), .b({n513, n513, n513, n513, n512, n512, n512, 
        n512, n512, n512, n512, n511, n511, n511, n511, n511, n511, n511, n510, 
        n510, n510, n510, n510, n510, n510, n509, n509, n509, n509, n509, n509, 
        n509, \p[1][31] , \p[1][30] , \p[1][29] , \p[1][28] , \p[1][27] , 
        \p[1][26] , \p[1][25] , \p[1][24] , \p[1][23] , \p[1][22] , \p[1][21] , 
        \p[1][20] , \p[1][19] , \p[1][18] , \p[1][17] , \p[1][16] , \p[1][15] , 
        \p[1][14] , \p[1][13] , \p[1][12] , \p[1][11] , \p[1][10] , \p[1][9] , 
        \p[1][8] , \p[1][7] , \p[1][6] , \p[1][5] , \p[1][4] , \p[1][3] , 
        \p[1][2] , \p[1][1] , 1'b0}), .cin({n517, n517, n517, n517, n517, n517, 
        n517, n516, n516, n516, n516, n516, n516, n516, n516, n515, n515, n515, 
        n515, n515, n515, n515, n515, n514, n514, n514, n514, n514, n514, n514, 
        n514, \p[2][32] , \p[2][31] , \p[2][30] , \p[2][29] , \p[2][28] , 
        \p[2][27] , \p[2][26] , \p[2][25] , \p[2][24] , \p[2][23] , \p[2][22] , 
        \p[2][21] , \p[2][20] , \p[2][19] , \p[2][18] , \p[2][17] , \p[2][16] , 
        \p[2][15] , \p[2][14] , \p[2][13] , \p[2][12] , \p[2][11] , \p[2][10] , 
        \p[2][9] , \p[2][8] , \p[2][7] , \p[2][6] , \p[2][5] , \p[2][4] , 
        \p[2][3] , \p[2][2] , 1'b0, 1'b0}), .sum({\g[0][63] , \g[0][62] , 
        \g[0][61] , \g[0][60] , \g[0][59] , \g[0][58] , \g[0][57] , \g[0][56] , 
        \g[0][55] , \g[0][54] , \g[0][53] , \g[0][52] , \g[0][51] , \g[0][50] , 
        \g[0][49] , \g[0][48] , \g[0][47] , \g[0][46] , \g[0][45] , \g[0][44] , 
        \g[0][43] , \g[0][42] , \g[0][41] , \g[0][40] , \g[0][39] , \g[0][38] , 
        \g[0][37] , \g[0][36] , \g[0][35] , \g[0][34] , \g[0][33] , \g[0][32] , 
        \g[0][31] , \g[0][30] , \g[0][29] , \g[0][28] , \g[0][27] , \g[0][26] , 
        \g[0][25] , \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , 
        \g[0][19] , \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] , 
        \g[0][13] , \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] , 
        \g[0][7] , \g[0][6] , \g[0][5] , \g[0][4] , \g[0][3] , \g[0][2] , 
        \g[0][1] , \g[0][0] }), .cout({\g[21][63] , \g[21][62] , \g[21][61] , 
        \g[21][60] , \g[21][59] , \g[21][58] , \g[21][57] , \g[21][56] , 
        \g[21][55] , \g[21][54] , \g[21][53] , \g[21][52] , \g[21][51] , 
        \g[21][50] , \g[21][49] , \g[21][48] , \g[21][47] , \g[21][46] , 
        \g[21][45] , \g[21][44] , \g[21][43] , \g[21][42] , \g[21][41] , 
        \g[21][40] , \g[21][39] , \g[21][38] , \g[21][37] , \g[21][36] , 
        \g[21][35] , \g[21][34] , \g[21][33] , \g[21][32] , \g[21][31] , 
        \g[21][30] , \g[21][29] , \g[21][28] , \g[21][27] , \g[21][26] , 
        \g[21][25] , \g[21][24] , \g[21][23] , \g[21][22] , \g[21][21] , 
        \g[21][20] , \g[21][19] , \g[21][18] , \g[21][17] , \g[21][16] , 
        \g[21][15] , \g[21][14] , \g[21][13] , \g[21][12] , \g[21][11] , 
        \g[21][10] , \g[21][9] , \g[21][8] , \g[21][7] , \g[21][6] , 
        \g[21][5] , \g[21][4] , \g[21][3] , \g[21][2] , \g[21][1] , 
        SYNOPSYS_UNCONNECTED__0}) );
  FullAdder_61 \level1[1].x6  ( .a({n522, n522, n522, n522, n522, n522, n521, 
        n521, n521, n521, n521, n521, n520, n520, n520, n520, n520, n520, n519, 
        n519, n519, n519, n519, n519, n518, n518, n518, n518, n518, n518, 
        \p[3][33] , \p[3][32] , \p[3][31] , \p[3][30] , \p[3][29] , \p[3][28] , 
        \p[3][27] , \p[3][26] , \p[3][25] , \p[3][24] , \p[3][23] , \p[3][22] , 
        \p[3][21] , \p[3][20] , \p[3][19] , \p[3][18] , \p[3][17] , \p[3][16] , 
        \p[3][15] , \p[3][14] , \p[3][13] , \p[3][12] , \p[3][11] , \p[3][10] , 
        \p[3][9] , \p[3][8] , \p[3][7] , \p[3][6] , \p[3][5] , \p[3][4] , 
        \p[3][3] , 1'b0, 1'b0, 1'b0}), .b({n525, n525, n525, n525, n525, n525, 
        n525, n525, n525, n524, n524, n524, n524, n524, n524, n524, n524, n524, 
        n524, n523, n523, n523, n523, n523, n523, n523, n523, n523, n523, 
        \p[4][34] , \p[4][33] , \p[4][32] , \p[4][31] , \p[4][30] , \p[4][29] , 
        \p[4][28] , \p[4][27] , \p[4][26] , \p[4][25] , \p[4][24] , \p[4][23] , 
        \p[4][22] , \p[4][21] , \p[4][20] , \p[4][19] , \p[4][18] , \p[4][17] , 
        \p[4][16] , \p[4][15] , \p[4][14] , \p[4][13] , \p[4][12] , \p[4][11] , 
        \p[4][10] , \p[4][9] , \p[4][8] , \p[4][7] , \p[4][6] , \p[4][5] , 
        \p[4][4] , 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n530, n530, n530, n530, 
        n529, n529, n529, n529, n529, n529, n528, n528, n528, n528, n528, n528, 
        n527, n527, n527, n527, n527, n527, n526, n526, n526, n526, n526, n526, 
        \p[5][35] , \p[5][34] , \p[5][33] , \p[5][32] , \p[5][31] , \p[5][30] , 
        \p[5][29] , \p[5][28] , \p[5][27] , \p[5][26] , \p[5][25] , \p[5][24] , 
        \p[5][23] , \p[5][22] , \p[5][21] , \p[5][20] , \p[5][19] , \p[5][18] , 
        \p[5][17] , \p[5][16] , \p[5][15] , \p[5][14] , \p[5][13] , \p[5][12] , 
        \p[5][11] , \p[5][10] , \p[5][9] , \p[5][8] , \p[5][7] , \p[5][6] , 
        \p[5][5] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[1][63] , 
        \g[1][62] , \g[1][61] , \g[1][60] , \g[1][59] , \g[1][58] , \g[1][57] , 
        \g[1][56] , \g[1][55] , \g[1][54] , \g[1][53] , \g[1][52] , \g[1][51] , 
        \g[1][50] , \g[1][49] , \g[1][48] , \g[1][47] , \g[1][46] , \g[1][45] , 
        \g[1][44] , \g[1][43] , \g[1][42] , \g[1][41] , \g[1][40] , \g[1][39] , 
        \g[1][38] , \g[1][37] , \g[1][36] , \g[1][35] , \g[1][34] , \g[1][33] , 
        \g[1][32] , \g[1][31] , \g[1][30] , \g[1][29] , \g[1][28] , \g[1][27] , 
        \g[1][26] , \g[1][25] , \g[1][24] , \g[1][23] , \g[1][22] , \g[1][21] , 
        \g[1][20] , \g[1][19] , \g[1][18] , \g[1][17] , \g[1][16] , \g[1][15] , 
        \g[1][14] , \g[1][13] , \g[1][12] , \g[1][11] , \g[1][10] , \g[1][9] , 
        \g[1][8] , \g[1][7] , \g[1][6] , \g[1][5] , \g[1][4] , \g[1][3] , 
        \g[1][2] , \g[1][1] , \g[1][0] }), .cout({\g[22][63] , \g[22][62] , 
        \g[22][61] , \g[22][60] , \g[22][59] , \g[22][58] , \g[22][57] , 
        \g[22][56] , \g[22][55] , \g[22][54] , \g[22][53] , \g[22][52] , 
        \g[22][51] , \g[22][50] , \g[22][49] , \g[22][48] , \g[22][47] , 
        \g[22][46] , \g[22][45] , \g[22][44] , \g[22][43] , \g[22][42] , 
        \g[22][41] , \g[22][40] , \g[22][39] , \g[22][38] , \g[22][37] , 
        \g[22][36] , \g[22][35] , \g[22][34] , \g[22][33] , \g[22][32] , 
        \g[22][31] , \g[22][30] , \g[22][29] , \g[22][28] , \g[22][27] , 
        \g[22][26] , \g[22][25] , \g[22][24] , \g[22][23] , \g[22][22] , 
        \g[22][21] , \g[22][20] , \g[22][19] , \g[22][18] , \g[22][17] , 
        \g[22][16] , \g[22][15] , \g[22][14] , \g[22][13] , \g[22][12] , 
        \g[22][11] , \g[22][10] , \g[22][9] , \g[22][8] , \g[22][7] , 
        \g[22][6] , \g[22][5] , \g[22][4] , \g[22][3] , \g[22][2] , \g[22][1] , 
        SYNOPSYS_UNCONNECTED__1}) );
  FullAdder_60 \level1[2].x6  ( .a({n535, n535, n535, n534, n534, n534, n534, 
        n534, n534, n533, n533, n533, n533, n533, n533, n532, n532, n532, n532, 
        n532, n532, n531, n531, n531, n531, n531, n531, \p[6][36] , \p[6][35] , 
        \p[6][34] , \p[6][33] , \p[6][32] , \p[6][31] , \p[6][30] , \p[6][29] , 
        \p[6][28] , \p[6][27] , \p[6][26] , \p[6][25] , \p[6][24] , \p[6][23] , 
        \p[6][22] , \p[6][21] , \p[6][20] , \p[6][19] , \p[6][18] , \p[6][17] , 
        \p[6][16] , \p[6][15] , \p[6][14] , \p[6][13] , \p[6][12] , \p[6][11] , 
        \p[6][10] , \p[6][9] , \p[6][8] , \p[6][7] , \p[6][6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .b({n539, n539, n539, n539, n539, n538, n538, 
        n538, n538, n538, n538, n538, n537, n537, n537, n537, n537, n537, n537, 
        n536, n536, n536, n536, n536, n536, n536, \p[7][37] , \p[7][36] , 
        \p[7][35] , \p[7][34] , \p[7][33] , \p[7][32] , \p[7][31] , \p[7][30] , 
        \p[7][29] , \p[7][28] , \p[7][27] , \p[7][26] , \p[7][25] , \p[7][24] , 
        \p[7][23] , \p[7][22] , \p[7][21] , \p[7][20] , \p[7][19] , \p[7][18] , 
        \p[7][17] , \p[7][16] , \p[7][15] , \p[7][14] , \p[7][13] , \p[7][12] , 
        \p[7][11] , \p[7][10] , \p[7][9] , \p[7][8] , \p[7][7] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n375, n375, n375, n375, n375, 
        n375, n375, n374, n374, n374, n374, n374, n374, n373, n373, n373, n373, 
        n373, n373, n372, n372, n372, n372, n372, n372, \p[8][38] , \p[8][37] , 
        \p[8][36] , \p[8][35] , \p[8][34] , \p[8][33] , \p[8][32] , \p[8][31] , 
        \p[8][30] , \p[8][29] , \p[8][28] , \p[8][27] , \p[8][26] , \p[8][25] , 
        \p[8][24] , \p[8][23] , \p[8][22] , \p[8][21] , \p[8][20] , \p[8][19] , 
        \p[8][18] , \p[8][17] , \p[8][16] , \p[8][15] , \p[8][14] , \p[8][13] , 
        \p[8][12] , \p[8][11] , \p[8][10] , \p[8][9] , \p[8][8] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[2][63] , \g[2][62] , 
        \g[2][61] , \g[2][60] , \g[2][59] , \g[2][58] , \g[2][57] , \g[2][56] , 
        \g[2][55] , \g[2][54] , \g[2][53] , \g[2][52] , \g[2][51] , \g[2][50] , 
        \g[2][49] , \g[2][48] , \g[2][47] , \g[2][46] , \g[2][45] , \g[2][44] , 
        \g[2][43] , \g[2][42] , \g[2][41] , \g[2][40] , \g[2][39] , \g[2][38] , 
        \g[2][37] , \g[2][36] , \g[2][35] , \g[2][34] , \g[2][33] , \g[2][32] , 
        \g[2][31] , \g[2][30] , \g[2][29] , \g[2][28] , \g[2][27] , \g[2][26] , 
        \g[2][25] , \g[2][24] , \g[2][23] , \g[2][22] , \g[2][21] , \g[2][20] , 
        \g[2][19] , \g[2][18] , \g[2][17] , \g[2][16] , \g[2][15] , \g[2][14] , 
        \g[2][13] , \g[2][12] , \g[2][11] , \g[2][10] , \g[2][9] , \g[2][8] , 
        \g[2][7] , \g[2][6] , \g[2][5] , \g[2][4] , \g[2][3] , \g[2][2] , 
        \g[2][1] , \g[2][0] }), .cout({\g[23][63] , \g[23][62] , \g[23][61] , 
        \g[23][60] , \g[23][59] , \g[23][58] , \g[23][57] , \g[23][56] , 
        \g[23][55] , \g[23][54] , \g[23][53] , \g[23][52] , \g[23][51] , 
        \g[23][50] , \g[23][49] , \g[23][48] , \g[23][47] , \g[23][46] , 
        \g[23][45] , \g[23][44] , \g[23][43] , \g[23][42] , \g[23][41] , 
        \g[23][40] , \g[23][39] , \g[23][38] , \g[23][37] , \g[23][36] , 
        \g[23][35] , \g[23][34] , \g[23][33] , \g[23][32] , \g[23][31] , 
        \g[23][30] , \g[23][29] , \g[23][28] , \g[23][27] , \g[23][26] , 
        \g[23][25] , \g[23][24] , \g[23][23] , \g[23][22] , \g[23][21] , 
        \g[23][20] , \g[23][19] , \g[23][18] , \g[23][17] , \g[23][16] , 
        \g[23][15] , \g[23][14] , \g[23][13] , \g[23][12] , \g[23][11] , 
        \g[23][10] , \g[23][9] , \g[23][8] , \g[23][7] , \g[23][6] , 
        \g[23][5] , \g[23][4] , \g[23][3] , \g[23][2] , \g[23][1] , 
        SYNOPSYS_UNCONNECTED__2}) );
  FullAdder_59 \level1[3].x6  ( .a({n379, n379, n379, n379, n379, n379, n378, 
        n378, n378, n378, n378, n378, n377, n377, n377, n377, n377, n377, n376, 
        n376, n376, n376, n376, n376, \p[9][39] , \p[9][38] , \p[9][37] , 
        \p[9][36] , \p[9][35] , \p[9][34] , \p[9][33] , \p[9][32] , \p[9][31] , 
        \p[9][30] , \p[9][29] , \p[9][28] , \p[9][27] , \p[9][26] , \p[9][25] , 
        \p[9][24] , \p[9][23] , \p[9][22] , \p[9][21] , \p[9][20] , \p[9][19] , 
        \p[9][18] , \p[9][17] , \p[9][16] , \p[9][15] , \p[9][14] , \p[9][13] , 
        \p[9][12] , \p[9][11] , \p[9][10] , \p[9][9] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n383, n383, n382, n382, n382, n382, 
        n382, n382, n382, n381, n381, n381, n381, n381, n381, n381, n380, n380, 
        n380, n380, n380, n380, n380, \p[10][40] , \p[10][39] , \p[10][38] , 
        \p[10][37] , \p[10][36] , \p[10][35] , \p[10][34] , \p[10][33] , 
        \p[10][32] , \p[10][31] , \p[10][30] , \p[10][29] , \p[10][28] , 
        \p[10][27] , \p[10][26] , \p[10][25] , \p[10][24] , \p[10][23] , 
        \p[10][22] , \p[10][21] , \p[10][20] , \p[10][19] , \p[10][18] , 
        \p[10][17] , \p[10][16] , \p[10][15] , \p[10][14] , \p[10][13] , 
        \p[10][12] , \p[10][11] , \p[10][10] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n387, n387, n387, n387, n386, 
        n386, n386, n386, n386, n386, n385, n385, n385, n385, n385, n385, n384, 
        n384, n384, n384, n384, n384, \p[11][41] , \p[11][40] , \p[11][39] , 
        \p[11][38] , \p[11][37] , \p[11][36] , \p[11][35] , \p[11][34] , 
        \p[11][33] , \p[11][32] , \p[11][31] , \p[11][30] , \p[11][29] , 
        \p[11][28] , \p[11][27] , \p[11][26] , \p[11][25] , \p[11][24] , 
        \p[11][23] , \p[11][22] , \p[11][21] , \p[11][20] , \p[11][19] , 
        \p[11][18] , \p[11][17] , \p[11][16] , \p[11][15] , \p[11][14] , 
        \p[11][13] , \p[11][12] , \p[11][11] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[3][63] , \g[3][62] , 
        \g[3][61] , \g[3][60] , \g[3][59] , \g[3][58] , \g[3][57] , \g[3][56] , 
        \g[3][55] , \g[3][54] , \g[3][53] , \g[3][52] , \g[3][51] , \g[3][50] , 
        \g[3][49] , \g[3][48] , \g[3][47] , \g[3][46] , \g[3][45] , \g[3][44] , 
        \g[3][43] , \g[3][42] , \g[3][41] , \g[3][40] , \g[3][39] , \g[3][38] , 
        \g[3][37] , \g[3][36] , \g[3][35] , \g[3][34] , \g[3][33] , \g[3][32] , 
        \g[3][31] , \g[3][30] , \g[3][29] , \g[3][28] , \g[3][27] , \g[3][26] , 
        \g[3][25] , \g[3][24] , \g[3][23] , \g[3][22] , \g[3][21] , \g[3][20] , 
        \g[3][19] , \g[3][18] , \g[3][17] , \g[3][16] , \g[3][15] , \g[3][14] , 
        \g[3][13] , \g[3][12] , \g[3][11] , \g[3][10] , \g[3][9] , \g[3][8] , 
        \g[3][7] , \g[3][6] , \g[3][5] , \g[3][4] , \g[3][3] , \g[3][2] , 
        \g[3][1] , \g[3][0] }), .cout({\g[24][63] , \g[24][62] , \g[24][61] , 
        \g[24][60] , \g[24][59] , \g[24][58] , \g[24][57] , \g[24][56] , 
        \g[24][55] , \g[24][54] , \g[24][53] , \g[24][52] , \g[24][51] , 
        \g[24][50] , \g[24][49] , \g[24][48] , \g[24][47] , \g[24][46] , 
        \g[24][45] , \g[24][44] , \g[24][43] , \g[24][42] , \g[24][41] , 
        \g[24][40] , \g[24][39] , \g[24][38] , \g[24][37] , \g[24][36] , 
        \g[24][35] , \g[24][34] , \g[24][33] , \g[24][32] , \g[24][31] , 
        \g[24][30] , \g[24][29] , \g[24][28] , \g[24][27] , \g[24][26] , 
        \g[24][25] , \g[24][24] , \g[24][23] , \g[24][22] , \g[24][21] , 
        \g[24][20] , \g[24][19] , \g[24][18] , \g[24][17] , \g[24][16] , 
        \g[24][15] , \g[24][14] , \g[24][13] , \g[24][12] , \g[24][11] , 
        \g[24][10] , \g[24][9] , \g[24][8] , \g[24][7] , \g[24][6] , 
        \g[24][5] , \g[24][4] , \g[24][3] , \g[24][2] , \g[24][1] , 
        SYNOPSYS_UNCONNECTED__3}) );
  FullAdder_58 \level1[4].x6  ( .a({n391, n391, n391, n390, n390, n390, n390, 
        n390, n390, n389, n389, n389, n389, n389, n389, n388, n388, n388, n388, 
        n388, n388, \p[12][42] , \p[12][41] , \p[12][40] , \p[12][39] , 
        \p[12][38] , \p[12][37] , \p[12][36] , \p[12][35] , \p[12][34] , 
        \p[12][33] , \p[12][32] , \p[12][31] , \p[12][30] , \p[12][29] , 
        \p[12][28] , \p[12][27] , \p[12][26] , \p[12][25] , \p[12][24] , 
        \p[12][23] , \p[12][22] , \p[12][21] , \p[12][20] , \p[12][19] , 
        \p[12][18] , \p[12][17] , \p[12][16] , \p[12][15] , \p[12][14] , 
        \p[12][13] , \p[12][12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n394, n394, n394, n394, n394, n394, 
        n393, n393, n393, n393, n393, n393, n393, n392, n392, n392, n392, n392, 
        n392, n392, \p[13][43] , \p[13][42] , \p[13][41] , \p[13][40] , 
        \p[13][39] , \p[13][38] , \p[13][37] , \p[13][36] , \p[13][35] , 
        \p[13][34] , \p[13][33] , \p[13][32] , \p[13][31] , \p[13][30] , 
        \p[13][29] , \p[13][28] , \p[13][27] , \p[13][26] , \p[13][25] , 
        \p[13][24] , \p[13][23] , \p[13][22] , \p[13][21] , \p[13][20] , 
        \p[13][19] , \p[13][18] , \p[13][17] , \p[13][16] , \p[13][15] , 
        \p[13][14] , \p[13][13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n396, n396, n396, n396, 
        n396, n396, n396, n395, n395, n395, n395, n395, n395, n395, n395, n395, 
        n395, n395, n395, \p[14][44] , \p[14][43] , \p[14][42] , \p[14][41] , 
        \p[14][40] , \p[14][39] , \p[14][38] , \p[14][37] , \p[14][36] , 
        \p[14][35] , \p[14][34] , \p[14][33] , \p[14][32] , \p[14][31] , 
        \p[14][30] , \p[14][29] , \p[14][28] , \p[14][27] , \p[14][26] , 
        \p[14][25] , \p[14][24] , \p[14][23] , \p[14][22] , \p[14][21] , 
        \p[14][20] , \p[14][19] , \p[14][18] , \p[14][17] , \p[14][16] , 
        \p[14][15] , \p[14][14] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[4][63] , 
        \g[4][62] , \g[4][61] , \g[4][60] , \g[4][59] , \g[4][58] , \g[4][57] , 
        \g[4][56] , \g[4][55] , \g[4][54] , \g[4][53] , \g[4][52] , \g[4][51] , 
        \g[4][50] , \g[4][49] , \g[4][48] , \g[4][47] , \g[4][46] , \g[4][45] , 
        \g[4][44] , \g[4][43] , \g[4][42] , \g[4][41] , \g[4][40] , \g[4][39] , 
        \g[4][38] , \g[4][37] , \g[4][36] , \g[4][35] , \g[4][34] , \g[4][33] , 
        \g[4][32] , \g[4][31] , \g[4][30] , \g[4][29] , \g[4][28] , \g[4][27] , 
        \g[4][26] , \g[4][25] , \g[4][24] , \g[4][23] , \g[4][22] , \g[4][21] , 
        \g[4][20] , \g[4][19] , \g[4][18] , \g[4][17] , \g[4][16] , \g[4][15] , 
        \g[4][14] , \g[4][13] , \g[4][12] , \g[4][11] , \g[4][10] , \g[4][9] , 
        \g[4][8] , \g[4][7] , \g[4][6] , \g[4][5] , \g[4][4] , \g[4][3] , 
        \g[4][2] , \g[4][1] , \g[4][0] }), .cout({\g[25][63] , \g[25][62] , 
        \g[25][61] , \g[25][60] , \g[25][59] , \g[25][58] , \g[25][57] , 
        \g[25][56] , \g[25][55] , \g[25][54] , \g[25][53] , \g[25][52] , 
        \g[25][51] , \g[25][50] , \g[25][49] , \g[25][48] , \g[25][47] , 
        \g[25][46] , \g[25][45] , \g[25][44] , \g[25][43] , \g[25][42] , 
        \g[25][41] , \g[25][40] , \g[25][39] , \g[25][38] , \g[25][37] , 
        \g[25][36] , \g[25][35] , \g[25][34] , \g[25][33] , \g[25][32] , 
        \g[25][31] , \g[25][30] , \g[25][29] , \g[25][28] , \g[25][27] , 
        \g[25][26] , \g[25][25] , \g[25][24] , \g[25][23] , \g[25][22] , 
        \g[25][21] , \g[25][20] , \g[25][19] , \g[25][18] , \g[25][17] , 
        \g[25][16] , \g[25][15] , \g[25][14] , \g[25][13] , \g[25][12] , 
        \g[25][11] , \g[25][10] , \g[25][9] , \g[25][8] , \g[25][7] , 
        \g[25][6] , \g[25][5] , \g[25][4] , \g[25][3] , \g[25][2] , \g[25][1] , 
        SYNOPSYS_UNCONNECTED__4}) );
  FullAdder_57 \level1[5].x6  ( .a({n399, n399, n399, n399, n399, n399, n398, 
        n398, n398, n398, n398, n398, n397, n397, n397, n397, n397, n397, 
        \p[15][45] , \p[15][44] , \p[15][43] , \p[15][42] , \p[15][41] , 
        \p[15][40] , \p[15][39] , \p[15][38] , \p[15][37] , \p[15][36] , 
        \p[15][35] , \p[15][34] , \p[15][33] , \p[15][32] , \p[15][31] , 
        \p[15][30] , \p[15][29] , \p[15][28] , \p[15][27] , \p[15][26] , 
        \p[15][25] , \p[15][24] , \p[15][23] , \p[15][22] , \p[15][21] , 
        \p[15][20] , \p[15][19] , \p[15][18] , \p[15][17] , \p[15][16] , 
        \p[15][15] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n402, n402, n402, n401, n401, 
        n401, n401, n401, n401, n401, n400, n400, n400, n400, n400, n400, n400, 
        \p[16][46] , \p[16][45] , \p[16][44] , \p[16][43] , \p[16][42] , 
        \p[16][41] , \p[16][40] , \p[16][39] , \p[16][38] , \p[16][37] , 
        \p[16][36] , \p[16][35] , \p[16][34] , \p[16][33] , \p[16][32] , 
        \p[16][31] , \p[16][30] , \p[16][29] , \p[16][28] , \p[16][27] , 
        \p[16][26] , \p[16][25] , \p[16][24] , \p[16][23] , \p[16][22] , 
        \p[16][21] , \p[16][20] , \p[16][19] , \p[16][18] , \p[16][17] , 
        \p[16][16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n405, n405, n405, 
        n405, n404, n404, n404, n404, n404, n404, n403, n403, n403, n403, n403, 
        n403, \p[17][47] , \p[17][46] , \p[17][45] , \p[17][44] , \p[17][43] , 
        \p[17][42] , \p[17][41] , \p[17][40] , \p[17][39] , \p[17][38] , 
        \p[17][37] , \p[17][36] , \p[17][35] , \p[17][34] , \p[17][33] , 
        \p[17][32] , \p[17][31] , \p[17][30] , \p[17][29] , \p[17][28] , 
        \p[17][27] , \p[17][26] , \p[17][25] , \p[17][24] , \p[17][23] , 
        \p[17][22] , \p[17][21] , \p[17][20] , \p[17][19] , \p[17][18] , 
        \p[17][17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[5][63] , 
        \g[5][62] , \g[5][61] , \g[5][60] , \g[5][59] , \g[5][58] , \g[5][57] , 
        \g[5][56] , \g[5][55] , \g[5][54] , \g[5][53] , \g[5][52] , \g[5][51] , 
        \g[5][50] , \g[5][49] , \g[5][48] , \g[5][47] , \g[5][46] , \g[5][45] , 
        \g[5][44] , \g[5][43] , \g[5][42] , \g[5][41] , \g[5][40] , \g[5][39] , 
        \g[5][38] , \g[5][37] , \g[5][36] , \g[5][35] , \g[5][34] , \g[5][33] , 
        \g[5][32] , \g[5][31] , \g[5][30] , \g[5][29] , \g[5][28] , \g[5][27] , 
        \g[5][26] , \g[5][25] , \g[5][24] , \g[5][23] , \g[5][22] , \g[5][21] , 
        \g[5][20] , \g[5][19] , \g[5][18] , \g[5][17] , \g[5][16] , \g[5][15] , 
        \g[5][14] , \g[5][13] , \g[5][12] , \g[5][11] , \g[5][10] , \g[5][9] , 
        \g[5][8] , \g[5][7] , \g[5][6] , \g[5][5] , \g[5][4] , \g[5][3] , 
        \g[5][2] , \g[5][1] , \g[5][0] }), .cout({\g[26][63] , \g[26][62] , 
        \g[26][61] , \g[26][60] , \g[26][59] , \g[26][58] , \g[26][57] , 
        \g[26][56] , \g[26][55] , \g[26][54] , \g[26][53] , \g[26][52] , 
        \g[26][51] , \g[26][50] , \g[26][49] , \g[26][48] , \g[26][47] , 
        \g[26][46] , \g[26][45] , \g[26][44] , \g[26][43] , \g[26][42] , 
        \g[26][41] , \g[26][40] , \g[26][39] , \g[26][38] , \g[26][37] , 
        \g[26][36] , \g[26][35] , \g[26][34] , \g[26][33] , \g[26][32] , 
        \g[26][31] , \g[26][30] , \g[26][29] , \g[26][28] , \g[26][27] , 
        \g[26][26] , \g[26][25] , \g[26][24] , \g[26][23] , \g[26][22] , 
        \g[26][21] , \g[26][20] , \g[26][19] , \g[26][18] , \g[26][17] , 
        \g[26][16] , \g[26][15] , \g[26][14] , \g[26][13] , \g[26][12] , 
        \g[26][11] , \g[26][10] , \g[26][9] , \g[26][8] , \g[26][7] , 
        \g[26][6] , \g[26][5] , \g[26][4] , \g[26][3] , \g[26][2] , \g[26][1] , 
        SYNOPSYS_UNCONNECTED__5}) );
  FullAdder_56 \level1[6].x6  ( .a({n408, n408, n408, n407, n407, n407, n407, 
        n407, n407, n406, n406, n406, n406, n406, n406, \p[18][48] , 
        \p[18][47] , \p[18][46] , \p[18][45] , \p[18][44] , \p[18][43] , 
        \p[18][42] , \p[18][41] , \p[18][40] , \p[18][39] , \p[18][38] , 
        \p[18][37] , \p[18][36] , \p[18][35] , \p[18][34] , \p[18][33] , 
        \p[18][32] , \p[18][31] , \p[18][30] , \p[18][29] , \p[18][28] , 
        \p[18][27] , \p[18][26] , \p[18][25] , \p[18][24] , \p[18][23] , 
        \p[18][22] , \p[18][21] , \p[18][20] , \p[18][19] , \p[18][18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n410, n410, n410, n410, n410, n410, 
        n410, n409, n409, n409, n409, n409, n409, n409, \p[19][49] , 
        \p[19][48] , \p[19][47] , \p[19][46] , \p[19][45] , \p[19][44] , 
        \p[19][43] , \p[19][42] , \p[19][41] , \p[19][40] , \p[19][39] , 
        \p[19][38] , \p[19][37] , \p[19][36] , \p[19][35] , \p[19][34] , 
        \p[19][33] , \p[19][32] , \p[19][31] , \p[19][30] , \p[19][29] , 
        \p[19][28] , \p[19][27] , \p[19][26] , \p[19][25] , \p[19][24] , 
        \p[19][23] , \p[19][22] , \p[19][21] , \p[19][20] , \p[19][19] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({n412, n412, n412, n412, 
        n412, n411, n411, n411, n411, n411, n411, n411, n411, \p[20][50] , 
        \p[20][49] , \p[20][48] , \p[20][47] , \p[20][46] , \p[20][45] , 
        \p[20][44] , \p[20][43] , \p[20][42] , \p[20][41] , \p[20][40] , 
        \p[20][39] , \p[20][38] , \p[20][37] , \p[20][36] , \p[20][35] , 
        \p[20][34] , \p[20][33] , \p[20][32] , \p[20][31] , \p[20][30] , 
        \p[20][29] , \p[20][28] , \p[20][27] , \p[20][26] , \p[20][25] , 
        \p[20][24] , \p[20][23] , \p[20][22] , \p[20][21] , \p[20][20] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[6][63] , 
        \g[6][62] , \g[6][61] , \g[6][60] , \g[6][59] , \g[6][58] , \g[6][57] , 
        \g[6][56] , \g[6][55] , \g[6][54] , \g[6][53] , \g[6][52] , \g[6][51] , 
        \g[6][50] , \g[6][49] , \g[6][48] , \g[6][47] , \g[6][46] , \g[6][45] , 
        \g[6][44] , \g[6][43] , \g[6][42] , \g[6][41] , \g[6][40] , \g[6][39] , 
        \g[6][38] , \g[6][37] , \g[6][36] , \g[6][35] , \g[6][34] , \g[6][33] , 
        \g[6][32] , \g[6][31] , \g[6][30] , \g[6][29] , \g[6][28] , \g[6][27] , 
        \g[6][26] , \g[6][25] , \g[6][24] , \g[6][23] , \g[6][22] , \g[6][21] , 
        \g[6][20] , \g[6][19] , \g[6][18] , \g[6][17] , \g[6][16] , \g[6][15] , 
        \g[6][14] , \g[6][13] , \g[6][12] , \g[6][11] , \g[6][10] , \g[6][9] , 
        \g[6][8] , \g[6][7] , \g[6][6] , \g[6][5] , \g[6][4] , \g[6][3] , 
        \g[6][2] , \g[6][1] , \g[6][0] }), .cout({\g[27][63] , \g[27][62] , 
        \g[27][61] , \g[27][60] , \g[27][59] , \g[27][58] , \g[27][57] , 
        \g[27][56] , \g[27][55] , \g[27][54] , \g[27][53] , \g[27][52] , 
        \g[27][51] , \g[27][50] , \g[27][49] , \g[27][48] , \g[27][47] , 
        \g[27][46] , \g[27][45] , \g[27][44] , \g[27][43] , \g[27][42] , 
        \g[27][41] , \g[27][40] , \g[27][39] , \g[27][38] , \g[27][37] , 
        \g[27][36] , \g[27][35] , \g[27][34] , \g[27][33] , \g[27][32] , 
        \g[27][31] , \g[27][30] , \g[27][29] , \g[27][28] , \g[27][27] , 
        \g[27][26] , \g[27][25] , \g[27][24] , \g[27][23] , \g[27][22] , 
        \g[27][21] , \g[27][20] , \g[27][19] , \g[27][18] , \g[27][17] , 
        \g[27][16] , \g[27][15] , \g[27][14] , \g[27][13] , \g[27][12] , 
        \g[27][11] , \g[27][10] , \g[27][9] , \g[27][8] , \g[27][7] , 
        \g[27][6] , \g[27][5] , \g[27][4] , \g[27][3] , \g[27][2] , \g[27][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  FullAdder_55 \level1[7].x6  ( .a({n154, n155, n154, n155, n154, n155, n154, 
        n155, n153, n153, n153, n153, \p[21][51] , \p[21][50] , \p[21][49] , 
        \p[21][48] , \p[21][47] , \p[21][46] , \p[21][45] , \p[21][44] , 
        \p[21][43] , \p[21][42] , \p[21][41] , \p[21][40] , \p[21][39] , 
        \p[21][38] , \p[21][37] , \p[21][36] , \p[21][35] , \p[21][34] , 
        \p[21][33] , \p[21][32] , \p[21][31] , \p[21][30] , \p[21][29] , 
        \p[21][28] , \p[21][27] , \p[21][26] , \p[21][25] , \p[21][24] , 
        \p[21][23] , \p[21][22] , \p[21][21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .b({\p[22][63] , \p[22][63] , \p[22][63] , 
        \p[22][63] , \p[22][63] , \p[22][63] , \p[22][63] , \p[22][63] , 
        \p[22][63] , \p[22][63] , \p[22][63] , \p[22][52] , \p[22][51] , 
        \p[22][50] , \p[22][49] , \p[22][48] , \p[22][47] , \p[22][46] , 
        \p[22][45] , \p[22][44] , \p[22][43] , \p[22][42] , \p[22][41] , 
        \p[22][40] , \p[22][39] , \p[22][38] , \p[22][37] , \p[22][36] , 
        \p[22][35] , \p[22][34] , \p[22][33] , \p[22][32] , \p[22][31] , 
        \p[22][30] , \p[22][29] , \p[22][28] , \p[22][27] , \p[22][26] , 
        \p[22][25] , \p[22][24] , \p[22][23] , \p[22][22] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[23][63] , 
        \p[23][63] , \p[23][63] , \p[23][63] , \p[23][63] , \p[23][63] , 
        \p[23][63] , \p[23][63] , \p[23][63] , \p[23][63] , \p[23][53] , 
        \p[23][52] , \p[23][51] , \p[23][50] , \p[23][49] , \p[23][48] , 
        \p[23][47] , \p[23][46] , \p[23][45] , \p[23][44] , \p[23][43] , 
        \p[23][42] , \p[23][41] , \p[23][40] , \p[23][39] , \p[23][38] , 
        \p[23][37] , \p[23][36] , \p[23][35] , \p[23][34] , \p[23][33] , 
        \p[23][32] , \p[23][31] , \p[23][30] , \p[23][29] , \p[23][28] , 
        \p[23][27] , \p[23][26] , \p[23][25] , \p[23][24] , \p[23][23] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({
        \g[7][63] , \g[7][62] , \g[7][61] , \g[7][60] , \g[7][59] , \g[7][58] , 
        \g[7][57] , \g[7][56] , \g[7][55] , \g[7][54] , \g[7][53] , \g[7][52] , 
        \g[7][51] , \g[7][50] , \g[7][49] , \g[7][48] , \g[7][47] , \g[7][46] , 
        \g[7][45] , \g[7][44] , \g[7][43] , \g[7][42] , \g[7][41] , \g[7][40] , 
        \g[7][39] , \g[7][38] , \g[7][37] , \g[7][36] , \g[7][35] , \g[7][34] , 
        \g[7][33] , \g[7][32] , \g[7][31] , \g[7][30] , \g[7][29] , \g[7][28] , 
        \g[7][27] , \g[7][26] , \g[7][25] , \g[7][24] , \g[7][23] , \g[7][22] , 
        \g[7][21] , \g[7][20] , \g[7][19] , \g[7][18] , \g[7][17] , \g[7][16] , 
        \g[7][15] , \g[7][14] , \g[7][13] , \g[7][12] , \g[7][11] , \g[7][10] , 
        \g[7][9] , \g[7][8] , \g[7][7] , \g[7][6] , \g[7][5] , \g[7][4] , 
        \g[7][3] , \g[7][2] , \g[7][1] , \g[7][0] }), .cout({\g[28][63] , 
        \g[28][62] , \g[28][61] , \g[28][60] , \g[28][59] , \g[28][58] , 
        \g[28][57] , \g[28][56] , \g[28][55] , \g[28][54] , \g[28][53] , 
        \g[28][52] , \g[28][51] , \g[28][50] , \g[28][49] , \g[28][48] , 
        \g[28][47] , \g[28][46] , \g[28][45] , \g[28][44] , \g[28][43] , 
        \g[28][42] , \g[28][41] , \g[28][40] , \g[28][39] , \g[28][38] , 
        \g[28][37] , \g[28][36] , \g[28][35] , \g[28][34] , \g[28][33] , 
        \g[28][32] , \g[28][31] , \g[28][30] , \g[28][29] , \g[28][28] , 
        \g[28][27] , \g[28][26] , \g[28][25] , \g[28][24] , \g[28][23] , 
        \g[28][22] , \g[28][21] , \g[28][20] , \g[28][19] , \g[28][18] , 
        \g[28][17] , \g[28][16] , \g[28][15] , \g[28][14] , \g[28][13] , 
        \g[28][12] , \g[28][11] , \g[28][10] , \g[28][9] , \g[28][8] , 
        \g[28][7] , \g[28][6] , \g[28][5] , \g[28][4] , \g[28][3] , \g[28][2] , 
        \g[28][1] , SYNOPSYS_UNCONNECTED__7}) );
  FullAdder_54 \level1[8].x6  ( .a({\p[24][63] , \p[24][63] , \p[24][63] , 
        \p[24][63] , \p[24][63] , \p[24][63] , \p[24][63] , \p[24][63] , 
        \p[24][63] , \p[24][54] , \p[24][53] , \p[24][52] , \p[24][51] , 
        \p[24][50] , \p[24][49] , \p[24][48] , \p[24][47] , \p[24][46] , 
        \p[24][45] , \p[24][44] , \p[24][43] , \p[24][42] , \p[24][41] , 
        \p[24][40] , \p[24][39] , \p[24][38] , \p[24][37] , \p[24][36] , 
        \p[24][35] , \p[24][34] , \p[24][33] , \p[24][32] , \p[24][31] , 
        \p[24][30] , \p[24][29] , \p[24][28] , \p[24][27] , \p[24][26] , 
        \p[24][25] , \p[24][24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({\p[25][63] , \p[25][63] , 
        \p[25][63] , \p[25][63] , \p[25][63] , \p[25][63] , \p[25][63] , 
        \p[25][63] , \p[25][55] , \p[25][54] , \p[25][53] , \p[25][52] , 
        \p[25][51] , \p[25][50] , \p[25][49] , \p[25][48] , \p[25][47] , 
        \p[25][46] , \p[25][45] , \p[25][44] , \p[25][43] , \p[25][42] , 
        \p[25][41] , \p[25][40] , \p[25][39] , \p[25][38] , \p[25][37] , 
        \p[25][36] , \p[25][35] , \p[25][34] , \p[25][33] , \p[25][32] , 
        \p[25][31] , \p[25][30] , \p[25][29] , \p[25][28] , \p[25][27] , 
        \p[25][26] , \p[25][25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[26][63] , \p[26][63] , 
        \p[26][63] , \p[26][63] , \p[26][63] , \p[26][63] , \p[26][63] , 
        \p[26][56] , \p[26][55] , \p[26][54] , \p[26][53] , \p[26][52] , 
        \p[26][51] , \p[26][50] , \p[26][49] , \p[26][48] , \p[26][47] , 
        \p[26][46] , \p[26][45] , \p[26][44] , \p[26][43] , \p[26][42] , 
        \p[26][41] , \p[26][40] , \p[26][39] , \p[26][38] , \p[26][37] , 
        \p[26][36] , \p[26][35] , \p[26][34] , \p[26][33] , \p[26][32] , 
        \p[26][31] , \p[26][30] , \p[26][29] , \p[26][28] , \p[26][27] , 
        \p[26][26] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[8][63] , \g[8][62] , 
        \g[8][61] , \g[8][60] , \g[8][59] , \g[8][58] , \g[8][57] , \g[8][56] , 
        \g[8][55] , \g[8][54] , \g[8][53] , \g[8][52] , \g[8][51] , \g[8][50] , 
        \g[8][49] , \g[8][48] , \g[8][47] , \g[8][46] , \g[8][45] , \g[8][44] , 
        \g[8][43] , \g[8][42] , \g[8][41] , \g[8][40] , \g[8][39] , \g[8][38] , 
        \g[8][37] , \g[8][36] , \g[8][35] , \g[8][34] , \g[8][33] , \g[8][32] , 
        \g[8][31] , \g[8][30] , \g[8][29] , \g[8][28] , \g[8][27] , \g[8][26] , 
        \g[8][25] , \g[8][24] , \g[8][23] , \g[8][22] , \g[8][21] , \g[8][20] , 
        \g[8][19] , \g[8][18] , \g[8][17] , \g[8][16] , \g[8][15] , \g[8][14] , 
        \g[8][13] , \g[8][12] , \g[8][11] , \g[8][10] , \g[8][9] , \g[8][8] , 
        \g[8][7] , \g[8][6] , \g[8][5] , \g[8][4] , \g[8][3] , \g[8][2] , 
        \g[8][1] , \g[8][0] }), .cout({\g[29][63] , \g[29][62] , \g[29][61] , 
        \g[29][60] , \g[29][59] , \g[29][58] , \g[29][57] , \g[29][56] , 
        \g[29][55] , \g[29][54] , \g[29][53] , \g[29][52] , \g[29][51] , 
        \g[29][50] , \g[29][49] , \g[29][48] , \g[29][47] , \g[29][46] , 
        \g[29][45] , \g[29][44] , \g[29][43] , \g[29][42] , \g[29][41] , 
        \g[29][40] , \g[29][39] , \g[29][38] , \g[29][37] , \g[29][36] , 
        \g[29][35] , \g[29][34] , \g[29][33] , \g[29][32] , \g[29][31] , 
        \g[29][30] , \g[29][29] , \g[29][28] , \g[29][27] , \g[29][26] , 
        \g[29][25] , \g[29][24] , \g[29][23] , \g[29][22] , \g[29][21] , 
        \g[29][20] , \g[29][19] , \g[29][18] , \g[29][17] , \g[29][16] , 
        \g[29][15] , \g[29][14] , \g[29][13] , \g[29][12] , \g[29][11] , 
        \g[29][10] , \g[29][9] , \g[29][8] , \g[29][7] , \g[29][6] , 
        \g[29][5] , \g[29][4] , \g[29][3] , \g[29][2] , \g[29][1] , 
        SYNOPSYS_UNCONNECTED__8}) );
  FullAdder_53 \level1[9].x6  ( .a({\p[27][63] , \p[27][63] , \p[27][63] , 
        \p[27][63] , \p[27][63] , \p[27][63] , \p[27][57] , \p[27][56] , 
        \p[27][55] , \p[27][54] , \p[27][53] , \p[27][52] , \p[27][51] , 
        \p[27][50] , \p[27][49] , \p[27][48] , \p[27][47] , \p[27][46] , 
        \p[27][45] , \p[27][44] , \p[27][43] , \p[27][42] , \p[27][41] , 
        \p[27][40] , \p[27][39] , \p[27][38] , \p[27][37] , \p[27][36] , 
        \p[27][35] , \p[27][34] , \p[27][33] , \p[27][32] , \p[27][31] , 
        \p[27][30] , \p[27][29] , \p[27][28] , \p[27][27] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({\p[28][63] , \p[28][63] , \p[28][63] , \p[28][63] , \p[28][63] , 
        \p[28][58] , \p[28][57] , \p[28][56] , \p[28][55] , \p[28][54] , 
        \p[28][53] , \p[28][52] , \p[28][51] , \p[28][50] , \p[28][49] , 
        \p[28][48] , \p[28][47] , \p[28][46] , \p[28][45] , \p[28][44] , 
        \p[28][43] , \p[28][42] , \p[28][41] , \p[28][40] , \p[28][39] , 
        \p[28][38] , \p[28][37] , \p[28][36] , \p[28][35] , \p[28][34] , 
        \p[28][33] , \p[28][32] , \p[28][31] , \p[28][30] , \p[28][29] , 
        \p[28][28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[29][63] , 
        \p[29][63] , \p[29][63] , \p[29][63] , \p[29][59] , \p[29][58] , 
        \p[29][57] , \p[29][56] , \p[29][55] , \p[29][54] , \p[29][53] , 
        \p[29][52] , \p[29][51] , \p[29][50] , \p[29][49] , \p[29][48] , 
        \p[29][47] , \p[29][46] , \p[29][45] , \p[29][44] , \p[29][43] , 
        \p[29][42] , \p[29][41] , \p[29][40] , \p[29][39] , \p[29][38] , 
        \p[29][37] , \p[29][36] , \p[29][35] , \p[29][34] , \p[29][33] , 
        \p[29][32] , \p[29][31] , \p[29][30] , \p[29][29] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .sum({\g[9][63] , \g[9][62] , \g[9][61] , \g[9][60] , 
        \g[9][59] , \g[9][58] , \g[9][57] , \g[9][56] , \g[9][55] , \g[9][54] , 
        \g[9][53] , \g[9][52] , \g[9][51] , \g[9][50] , \g[9][49] , \g[9][48] , 
        \g[9][47] , \g[9][46] , \g[9][45] , \g[9][44] , \g[9][43] , \g[9][42] , 
        \g[9][41] , \g[9][40] , \g[9][39] , \g[9][38] , \g[9][37] , \g[9][36] , 
        \g[9][35] , \g[9][34] , \g[9][33] , \g[9][32] , \g[9][31] , \g[9][30] , 
        \g[9][29] , \g[9][28] , \g[9][27] , \g[9][26] , \g[9][25] , \g[9][24] , 
        \g[9][23] , \g[9][22] , \g[9][21] , \g[9][20] , \g[9][19] , \g[9][18] , 
        \g[9][17] , \g[9][16] , \g[9][15] , \g[9][14] , \g[9][13] , \g[9][12] , 
        \g[9][11] , \g[9][10] , \g[9][9] , \g[9][8] , \g[9][7] , \g[9][6] , 
        \g[9][5] , \g[9][4] , \g[9][3] , \g[9][2] , \g[9][1] , \g[9][0] }), 
        .cout({\g[30][63] , \g[30][62] , \g[30][61] , \g[30][60] , \g[30][59] , 
        \g[30][58] , \g[30][57] , \g[30][56] , \g[30][55] , \g[30][54] , 
        \g[30][53] , \g[30][52] , \g[30][51] , \g[30][50] , \g[30][49] , 
        \g[30][48] , \g[30][47] , \g[30][46] , \g[30][45] , \g[30][44] , 
        \g[30][43] , \g[30][42] , \g[30][41] , \g[30][40] , \g[30][39] , 
        \g[30][38] , \g[30][37] , \g[30][36] , \g[30][35] , \g[30][34] , 
        \g[30][33] , \g[30][32] , \g[30][31] , \g[30][30] , \g[30][29] , 
        \g[30][28] , \g[30][27] , \g[30][26] , \g[30][25] , \g[30][24] , 
        \g[30][23] , \g[30][22] , \g[30][21] , \g[30][20] , \g[30][19] , 
        \g[30][18] , \g[30][17] , \g[30][16] , \g[30][15] , \g[30][14] , 
        \g[30][13] , \g[30][12] , \g[30][11] , \g[30][10] , \g[30][9] , 
        \g[30][8] , \g[30][7] , \g[30][6] , \g[30][5] , \g[30][4] , \g[30][3] , 
        \g[30][2] , \g[30][1] , SYNOPSYS_UNCONNECTED__9}) );
  FullAdder_52 \level1[10].x6  ( .a({\p[30][63] , \p[30][63] , \p[30][63] , 
        \p[30][60] , \p[30][59] , \p[30][58] , \p[30][57] , \p[30][56] , 
        \p[30][55] , \p[30][54] , \p[30][53] , \p[30][52] , \p[30][51] , 
        \p[30][50] , \p[30][49] , \p[30][48] , \p[30][47] , \p[30][46] , 
        \p[30][45] , \p[30][44] , \p[30][43] , \p[30][42] , \p[30][41] , 
        \p[30][40] , \p[30][39] , \p[30][38] , \p[30][37] , \p[30][36] , 
        \p[30][35] , \p[30][34] , \p[30][33] , \p[30][32] , \p[30][31] , 
        \p[30][30] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({
        \p[32][63] , \p[32][63] , \p[33][63] , \p[34][63] , \p[35][63] , 
        \p[36][63] , \p[37][63] , \p[38][63] , \p[39][63] , \p[40][63] , 
        \p[41][63] , n157, n414, n416, n421, n424, n427, n430, n433, n436, 
        n443, n447, n451, n454, n458, n463, n472, n476, n482, n487, n491, n497, 
        n502, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[32][63] , 
        \p[33][63] , \p[34][63] , \p[35][63] , \p[36][63] , \p[37][63] , 
        \p[38][63] , \p[39][63] , \p[40][63] , \p[41][63] , n156, n413, n415, 
        n418, n422, n425, n428, n431, n434, n438, n444, n449, n453, n457, n460, 
        n466, n474, n478, n483, n488, n493, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .sum({\g[10][63] , \g[10][62] , \g[10][61] , 
        \g[10][60] , \g[10][59] , \g[10][58] , \g[10][57] , \g[10][56] , 
        \g[10][55] , \g[10][54] , \g[10][53] , \g[10][52] , \g[10][51] , 
        \g[10][50] , \g[10][49] , \g[10][48] , \g[10][47] , \g[10][46] , 
        \g[10][45] , \g[10][44] , \g[10][43] , \g[10][42] , \g[10][41] , 
        \g[10][40] , \g[10][39] , \g[10][38] , \g[10][37] , \g[10][36] , 
        \g[10][35] , \g[10][34] , \g[10][33] , \g[10][32] , \g[10][31] , 
        \g[10][30] , \g[10][29] , \g[10][28] , \g[10][27] , \g[10][26] , 
        \g[10][25] , \g[10][24] , \g[10][23] , \g[10][22] , \g[10][21] , 
        \g[10][20] , \g[10][19] , \g[10][18] , \g[10][17] , \g[10][16] , 
        \g[10][15] , \g[10][14] , \g[10][13] , \g[10][12] , \g[10][11] , 
        \g[10][10] , \g[10][9] , \g[10][8] , \g[10][7] , \g[10][6] , 
        \g[10][5] , \g[10][4] , \g[10][3] , \g[10][2] , \g[10][1] , \g[10][0] }), .cout({\g[31][63] , \g[31][62] , \g[31][61] , \g[31][60] , \g[31][59] , 
        \g[31][58] , \g[31][57] , \g[31][56] , \g[31][55] , \g[31][54] , 
        \g[31][53] , \g[31][52] , \g[31][51] , \g[31][50] , \g[31][49] , 
        \g[31][48] , \g[31][47] , \g[31][46] , \g[31][45] , \g[31][44] , 
        \g[31][43] , \g[31][42] , \g[31][41] , \g[31][40] , \g[31][39] , 
        \g[31][38] , \g[31][37] , \g[31][36] , \g[31][35] , \g[31][34] , 
        \g[31][33] , \g[31][32] , \g[31][31] , \g[31][30] , \g[31][29] , 
        \g[31][28] , \g[31][27] , \g[31][26] , \g[31][25] , \g[31][24] , 
        \g[31][23] , \g[31][22] , \g[31][21] , \g[31][20] , \g[31][19] , 
        \g[31][18] , \g[31][17] , \g[31][16] , \g[31][15] , \g[31][14] , 
        \g[31][13] , \g[31][12] , \g[31][11] , \g[31][10] , \g[31][9] , 
        \g[31][8] , \g[31][7] , \g[31][6] , \g[31][5] , \g[31][4] , \g[31][3] , 
        \g[31][2] , \g[31][1] , SYNOPSYS_UNCONNECTED__10}) );
  FullAdder_51 \level1[11].x6  ( .a({\p[33][63] , \p[34][63] , \p[35][63] , 
        \p[36][63] , \p[37][63] , \p[38][63] , \p[39][63] , \p[40][63] , 
        \p[41][63] , n158, n413, n415, n418, n423, n426, n429, n432, n435, 
        n439, n445, n449, n453, n458, n461, n467, n475, n479, n485, n489, n496, 
        n501, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({
        \p[34][63] , \p[35][63] , \p[36][63] , \p[37][63] , \p[38][63] , 
        \p[39][63] , \p[40][63] , \p[41][63] , n158, n414, n416, n421, n424, 
        n427, n430, n433, n436, n442, n446, n451, n454, n458, n463, n471, n476, 
        n482, n486, n492, n497, n502, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .cin({\p[35][63] , \p[36][63] , \p[37][63] , 
        \p[38][63] , \p[39][63] , \p[40][63] , \p[41][63] , n156, n413, n415, 
        n417, n422, n425, n428, n431, n434, n437, n444, n448, n452, n456, n460, 
        n464, n473, n478, n484, n488, n493, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[11][63] , \g[11][62] , 
        \g[11][61] , \g[11][60] , \g[11][59] , \g[11][58] , \g[11][57] , 
        \g[11][56] , \g[11][55] , \g[11][54] , \g[11][53] , \g[11][52] , 
        \g[11][51] , \g[11][50] , \g[11][49] , \g[11][48] , \g[11][47] , 
        \g[11][46] , \g[11][45] , \g[11][44] , \g[11][43] , \g[11][42] , 
        \g[11][41] , \g[11][40] , \g[11][39] , \g[11][38] , \g[11][37] , 
        \g[11][36] , \g[11][35] , \g[11][34] , \g[11][33] , \g[11][32] , 
        \g[11][31] , \g[11][30] , \g[11][29] , \g[11][28] , \g[11][27] , 
        \g[11][26] , \g[11][25] , \g[11][24] , \g[11][23] , \g[11][22] , 
        \g[11][21] , \g[11][20] , \g[11][19] , \g[11][18] , \g[11][17] , 
        \g[11][16] , \g[11][15] , \g[11][14] , \g[11][13] , \g[11][12] , 
        \g[11][11] , \g[11][10] , \g[11][9] , \g[11][8] , \g[11][7] , 
        \g[11][6] , \g[11][5] , \g[11][4] , \g[11][3] , \g[11][2] , \g[11][1] , 
        \g[11][0] }), .cout({\g[32][63] , \g[32][62] , \g[32][61] , 
        \g[32][60] , \g[32][59] , \g[32][58] , \g[32][57] , \g[32][56] , 
        \g[32][55] , \g[32][54] , \g[32][53] , \g[32][52] , \g[32][51] , 
        \g[32][50] , \g[32][49] , \g[32][48] , \g[32][47] , \g[32][46] , 
        \g[32][45] , \g[32][44] , \g[32][43] , \g[32][42] , \g[32][41] , 
        \g[32][40] , \g[32][39] , \g[32][38] , \g[32][37] , \g[32][36] , 
        \g[32][35] , \g[32][34] , \g[32][33] , \g[32][32] , \g[32][31] , 
        \g[32][30] , \g[32][29] , \g[32][28] , \g[32][27] , \g[32][26] , 
        \g[32][25] , \g[32][24] , \g[32][23] , \g[32][22] , \g[32][21] , 
        \g[32][20] , \g[32][19] , \g[32][18] , \g[32][17] , \g[32][16] , 
        \g[32][15] , \g[32][14] , \g[32][13] , \g[32][12] , \g[32][11] , 
        \g[32][10] , \g[32][9] , \g[32][8] , \g[32][7] , \g[32][6] , 
        \g[32][5] , \g[32][4] , \g[32][3] , \g[32][2] , \g[32][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  FullAdder_50 \level1[12].x6  ( .a({\p[36][63] , \p[37][63] , \p[38][63] , 
        \p[39][63] , \p[40][63] , \p[41][63] , n157, n414, n416, n419, n422, 
        n426, n429, n432, n435, n439, n445, n449, n454, n458, n461, n467, n475, 
        n479, n484, n490, n496, n501, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({\p[37][63] , \p[38][63] , 
        \p[39][63] , \p[40][63] , \p[41][63] , n157, n414, n416, n420, n423, 
        n426, n430, n433, n436, n442, n446, n450, n454, n459, n463, n471, n476, 
        n481, n486, n492, n497, n502, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({\p[38][63] , \p[39][63] , 
        \p[40][63] , \p[41][63] , n156, n413, n415, n417, n422, n425, n428, 
        n431, n434, n437, n444, n448, n452, n456, n460, n464, n474, n478, n484, 
        n488, n493, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[12][63] , \g[12][62] , 
        \g[12][61] , \g[12][60] , \g[12][59] , \g[12][58] , \g[12][57] , 
        \g[12][56] , \g[12][55] , \g[12][54] , \g[12][53] , \g[12][52] , 
        \g[12][51] , \g[12][50] , \g[12][49] , \g[12][48] , \g[12][47] , 
        \g[12][46] , \g[12][45] , \g[12][44] , \g[12][43] , \g[12][42] , 
        \g[12][41] , \g[12][40] , \g[12][39] , \g[12][38] , \g[12][37] , 
        \g[12][36] , \g[12][35] , \g[12][34] , \g[12][33] , \g[12][32] , 
        \g[12][31] , \g[12][30] , \g[12][29] , \g[12][28] , \g[12][27] , 
        \g[12][26] , \g[12][25] , \g[12][24] , \g[12][23] , \g[12][22] , 
        \g[12][21] , \g[12][20] , \g[12][19] , \g[12][18] , \g[12][17] , 
        \g[12][16] , \g[12][15] , \g[12][14] , \g[12][13] , \g[12][12] , 
        \g[12][11] , \g[12][10] , \g[12][9] , \g[12][8] , \g[12][7] , 
        \g[12][6] , \g[12][5] , \g[12][4] , \g[12][3] , \g[12][2] , \g[12][1] , 
        \g[12][0] }), .cout({\g[33][63] , \g[33][62] , \g[33][61] , 
        \g[33][60] , \g[33][59] , \g[33][58] , \g[33][57] , \g[33][56] , 
        \g[33][55] , \g[33][54] , \g[33][53] , \g[33][52] , \g[33][51] , 
        \g[33][50] , \g[33][49] , \g[33][48] , \g[33][47] , \g[33][46] , 
        \g[33][45] , \g[33][44] , \g[33][43] , \g[33][42] , \g[33][41] , 
        \g[33][40] , \g[33][39] , \g[33][38] , \g[33][37] , \g[33][36] , 
        \g[33][35] , \g[33][34] , \g[33][33] , \g[33][32] , \g[33][31] , 
        \g[33][30] , \g[33][29] , \g[33][28] , \g[33][27] , \g[33][26] , 
        \g[33][25] , \g[33][24] , \g[33][23] , \g[33][22] , \g[33][21] , 
        \g[33][20] , \g[33][19] , \g[33][18] , \g[33][17] , \g[33][16] , 
        \g[33][15] , \g[33][14] , \g[33][13] , \g[33][12] , \g[33][11] , 
        \g[33][10] , \g[33][9] , \g[33][8] , \g[33][7] , \g[33][6] , 
        \g[33][5] , \g[33][4] , \g[33][3] , \g[33][2] , \g[33][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  FullAdder_49 \level1[13].x6  ( .a({\p[39][63] , \p[40][63] , \p[41][63] , 
        n158, n414, n416, n419, n423, n426, n429, n432, n435, n440, n445, n449, 
        n454, n458, n461, n467, n475, n480, n484, n490, n495, n501, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .b({\p[40][63] , \p[41][63] , n158, n414, n416, n420, n423, 
        n426, n429, n433, n436, n441, n446, n450, n454, n459, n462, n470, n476, 
        n481, n486, n492, n496, n502, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .cin({
        \p[41][63] , n156, n413, n415, n418, n422, n425, n428, n431, n434, 
        n438, n444, n448, n453, n457, n460, n465, n473, n478, n484, n488, n493, 
        n499, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[13][63] , \g[13][62] , 
        \g[13][61] , \g[13][60] , \g[13][59] , \g[13][58] , \g[13][57] , 
        \g[13][56] , \g[13][55] , \g[13][54] , \g[13][53] , \g[13][52] , 
        \g[13][51] , \g[13][50] , \g[13][49] , \g[13][48] , \g[13][47] , 
        \g[13][46] , \g[13][45] , \g[13][44] , \g[13][43] , \g[13][42] , 
        \g[13][41] , \g[13][40] , \g[13][39] , \g[13][38] , \g[13][37] , 
        \g[13][36] , \g[13][35] , \g[13][34] , \g[13][33] , \g[13][32] , 
        \g[13][31] , \g[13][30] , \g[13][29] , \g[13][28] , \g[13][27] , 
        \g[13][26] , \g[13][25] , \g[13][24] , \g[13][23] , \g[13][22] , 
        \g[13][21] , \g[13][20] , \g[13][19] , \g[13][18] , \g[13][17] , 
        \g[13][16] , \g[13][15] , \g[13][14] , \g[13][13] , \g[13][12] , 
        \g[13][11] , \g[13][10] , \g[13][9] , \g[13][8] , \g[13][7] , 
        \g[13][6] , \g[13][5] , \g[13][4] , \g[13][3] , \g[13][2] , \g[13][1] , 
        \g[13][0] }), .cout({\g[34][63] , \g[34][62] , \g[34][61] , 
        \g[34][60] , \g[34][59] , \g[34][58] , \g[34][57] , \g[34][56] , 
        \g[34][55] , \g[34][54] , \g[34][53] , \g[34][52] , \g[34][51] , 
        \g[34][50] , \g[34][49] , \g[34][48] , \g[34][47] , \g[34][46] , 
        \g[34][45] , \g[34][44] , \g[34][43] , \g[34][42] , \g[34][41] , 
        \g[34][40] , \g[34][39] , \g[34][38] , \g[34][37] , \g[34][36] , 
        \g[34][35] , \g[34][34] , \g[34][33] , \g[34][32] , \g[34][31] , 
        \g[34][30] , \g[34][29] , \g[34][28] , \g[34][27] , \g[34][26] , 
        \g[34][25] , \g[34][24] , \g[34][23] , \g[34][22] , \g[34][21] , 
        \g[34][20] , \g[34][19] , \g[34][18] , \g[34][17] , \g[34][16] , 
        \g[34][15] , \g[34][14] , \g[34][13] , \g[34][12] , \g[34][11] , 
        \g[34][10] , \g[34][9] , \g[34][8] , \g[34][7] , \g[34][6] , 
        \g[34][5] , \g[34][4] , \g[34][3] , \g[34][2] , \g[34][1] , 
        SYNOPSYS_UNCONNECTED__13}) );
  FullAdder_48 \level1[14].x6  ( .a({n157, n413, n415, n419, n423, n426, n429, 
        n432, n435, n440, n446, n449, n454, n458, n461, n468, n475, n479, n485, 
        n490, n495, n500, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n413, n416, 
        n420, n424, n427, n430, n433, n436, n442, n446, n450, n455, n459, n463, 
        n470, n476, n481, n486, n492, n496, n501, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n415, n417, n422, n425, n428, n431, n434, n439, 
        n444, n448, n452, n456, n460, n466, n474, n479, n483, n489, n494, n499, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[14][63] , 
        \g[14][62] , \g[14][61] , \g[14][60] , \g[14][59] , \g[14][58] , 
        \g[14][57] , \g[14][56] , \g[14][55] , \g[14][54] , \g[14][53] , 
        \g[14][52] , \g[14][51] , \g[14][50] , \g[14][49] , \g[14][48] , 
        \g[14][47] , \g[14][46] , \g[14][45] , \g[14][44] , \g[14][43] , 
        \g[14][42] , \g[14][41] , \g[14][40] , \g[14][39] , \g[14][38] , 
        \g[14][37] , \g[14][36] , \g[14][35] , \g[14][34] , \g[14][33] , 
        \g[14][32] , \g[14][31] , \g[14][30] , \g[14][29] , \g[14][28] , 
        \g[14][27] , \g[14][26] , \g[14][25] , \g[14][24] , \g[14][23] , 
        \g[14][22] , \g[14][21] , \g[14][20] , \g[14][19] , \g[14][18] , 
        \g[14][17] , \g[14][16] , \g[14][15] , \g[14][14] , \g[14][13] , 
        \g[14][12] , \g[14][11] , \g[14][10] , \g[14][9] , \g[14][8] , 
        \g[14][7] , \g[14][6] , \g[14][5] , \g[14][4] , \g[14][3] , \g[14][2] , 
        \g[14][1] , \g[14][0] }), .cout({\g[35][63] , \g[35][62] , \g[35][61] , 
        \g[35][60] , \g[35][59] , \g[35][58] , \g[35][57] , \g[35][56] , 
        \g[35][55] , \g[35][54] , \g[35][53] , \g[35][52] , \g[35][51] , 
        \g[35][50] , \g[35][49] , \g[35][48] , \g[35][47] , \g[35][46] , 
        \g[35][45] , \g[35][44] , \g[35][43] , \g[35][42] , \g[35][41] , 
        \g[35][40] , \g[35][39] , \g[35][38] , \g[35][37] , \g[35][36] , 
        \g[35][35] , \g[35][34] , \g[35][33] , \g[35][32] , \g[35][31] , 
        \g[35][30] , \g[35][29] , \g[35][28] , \g[35][27] , \g[35][26] , 
        \g[35][25] , \g[35][24] , \g[35][23] , \g[35][22] , \g[35][21] , 
        \g[35][20] , \g[35][19] , \g[35][18] , \g[35][17] , \g[35][16] , 
        \g[35][15] , \g[35][14] , \g[35][13] , \g[35][12] , \g[35][11] , 
        \g[35][10] , \g[35][9] , \g[35][8] , \g[35][7] , \g[35][6] , 
        \g[35][5] , \g[35][4] , \g[35][3] , \g[35][2] , \g[35][1] , 
        SYNOPSYS_UNCONNECTED__14}) );
  FullAdder_47 \level1[15].x6  ( .a({n420, n423, n425, n429, n432, n435, n440, 
        n445, n450, n453, n457, n462, n468, n475, n480, n485, n490, n495, n500, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n423, n427, 
        n430, n433, n436, n441, n446, n450, n455, n459, n462, n469, n476, n481, 
        n486, n492, n496, n501, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n425, n428, n431, n434, n438, n445, n448, n452, 
        n456, n461, n465, n473, n478, n484, n489, n494, n499, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[15][63] , 
        \g[15][62] , \g[15][61] , \g[15][60] , \g[15][59] , \g[15][58] , 
        \g[15][57] , \g[15][56] , \g[15][55] , \g[15][54] , \g[15][53] , 
        \g[15][52] , \g[15][51] , \g[15][50] , \g[15][49] , \g[15][48] , 
        \g[15][47] , \g[15][46] , \g[15][45] , \g[15][44] , \g[15][43] , 
        \g[15][42] , \g[15][41] , \g[15][40] , \g[15][39] , \g[15][38] , 
        \g[15][37] , \g[15][36] , \g[15][35] , \g[15][34] , \g[15][33] , 
        \g[15][32] , \g[15][31] , \g[15][30] , \g[15][29] , \g[15][28] , 
        \g[15][27] , \g[15][26] , \g[15][25] , \g[15][24] , \g[15][23] , 
        \g[15][22] , \g[15][21] , \g[15][20] , \g[15][19] , \g[15][18] , 
        \g[15][17] , \g[15][16] , \g[15][15] , \g[15][14] , \g[15][13] , 
        \g[15][12] , \g[15][11] , \g[15][10] , \g[15][9] , \g[15][8] , 
        \g[15][7] , \g[15][6] , \g[15][5] , \g[15][4] , \g[15][3] , \g[15][2] , 
        \g[15][1] , \g[15][0] }), .cout({\g[36][63] , \g[36][62] , \g[36][61] , 
        \g[36][60] , \g[36][59] , \g[36][58] , \g[36][57] , \g[36][56] , 
        \g[36][55] , \g[36][54] , \g[36][53] , \g[36][52] , \g[36][51] , 
        \g[36][50] , \g[36][49] , \g[36][48] , \g[36][47] , \g[36][46] , 
        \g[36][45] , \g[36][44] , \g[36][43] , \g[36][42] , \g[36][41] , 
        \g[36][40] , \g[36][39] , \g[36][38] , \g[36][37] , \g[36][36] , 
        \g[36][35] , \g[36][34] , \g[36][33] , \g[36][32] , \g[36][31] , 
        \g[36][30] , \g[36][29] , \g[36][28] , \g[36][27] , \g[36][26] , 
        \g[36][25] , \g[36][24] , \g[36][23] , \g[36][22] , \g[36][21] , 
        \g[36][20] , \g[36][19] , \g[36][18] , \g[36][17] , \g[36][16] , 
        \g[36][15] , \g[36][14] , \g[36][13] , \g[36][12] , \g[36][11] , 
        \g[36][10] , \g[36][9] , \g[36][8] , \g[36][7] , \g[36][6] , 
        \g[36][5] , \g[36][4] , \g[36][3] , \g[36][2] , \g[36][1] , 
        SYNOPSYS_UNCONNECTED__15}) );
  FullAdder_46 \level1[16].x6  ( .a({n429, n432, n435, n441, n446, n450, n453, 
        n457, n462, n468, n475, n480, n485, n491, n495, n500, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n432, n436, 
        n443, n447, n450, n455, n459, n463, n471, n476, n481, n486, n491, n496, 
        n501, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n435, n437, n444, n448, n452, n456, n461, n466, 
        n473, n479, n483, n488, n494, n499, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[16][63] , 
        \g[16][62] , \g[16][61] , \g[16][60] , \g[16][59] , \g[16][58] , 
        \g[16][57] , \g[16][56] , \g[16][55] , \g[16][54] , \g[16][53] , 
        \g[16][52] , \g[16][51] , \g[16][50] , \g[16][49] , \g[16][48] , 
        \g[16][47] , \g[16][46] , \g[16][45] , \g[16][44] , \g[16][43] , 
        \g[16][42] , \g[16][41] , \g[16][40] , \g[16][39] , \g[16][38] , 
        \g[16][37] , \g[16][36] , \g[16][35] , \g[16][34] , \g[16][33] , 
        \g[16][32] , \g[16][31] , \g[16][30] , \g[16][29] , \g[16][28] , 
        \g[16][27] , \g[16][26] , \g[16][25] , \g[16][24] , \g[16][23] , 
        \g[16][22] , \g[16][21] , \g[16][20] , \g[16][19] , \g[16][18] , 
        \g[16][17] , \g[16][16] , \g[16][15] , \g[16][14] , \g[16][13] , 
        \g[16][12] , \g[16][11] , \g[16][10] , \g[16][9] , \g[16][8] , 
        \g[16][7] , \g[16][6] , \g[16][5] , \g[16][4] , \g[16][3] , \g[16][2] , 
        \g[16][1] , \g[16][0] }), .cout({\g[37][63] , \g[37][62] , \g[37][61] , 
        \g[37][60] , \g[37][59] , \g[37][58] , \g[37][57] , \g[37][56] , 
        \g[37][55] , \g[37][54] , \g[37][53] , \g[37][52] , \g[37][51] , 
        \g[37][50] , \g[37][49] , \g[37][48] , \g[37][47] , \g[37][46] , 
        \g[37][45] , \g[37][44] , \g[37][43] , \g[37][42] , \g[37][41] , 
        \g[37][40] , \g[37][39] , \g[37][38] , \g[37][37] , \g[37][36] , 
        \g[37][35] , \g[37][34] , \g[37][33] , \g[37][32] , \g[37][31] , 
        \g[37][30] , \g[37][29] , \g[37][28] , \g[37][27] , \g[37][26] , 
        \g[37][25] , \g[37][24] , \g[37][23] , \g[37][22] , \g[37][21] , 
        \g[37][20] , \g[37][19] , \g[37][18] , \g[37][17] , \g[37][16] , 
        \g[37][15] , \g[37][14] , \g[37][13] , \g[37][12] , \g[37][11] , 
        \g[37][10] , \g[37][9] , \g[37][8] , \g[37][7] , \g[37][6] , 
        \g[37][5] , \g[37][4] , \g[37][3] , \g[37][2] , \g[37][1] , 
        SYNOPSYS_UNCONNECTED__16}) );
  FullAdder_45 \level1[17].x6  ( .a({n441, n445, n449, n453, n457, n462, n469, 
        n474, n480, n485, n491, n494, n500, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n445, n451, 
        n455, n459, n463, n470, n477, n481, n487, n491, n496, n501, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n449, n452, n456, n460, n464, n473, n479, n483, 
        n489, n494, n499, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[17][63] , 
        \g[17][62] , \g[17][61] , \g[17][60] , \g[17][59] , \g[17][58] , 
        \g[17][57] , \g[17][56] , \g[17][55] , \g[17][54] , \g[17][53] , 
        \g[17][52] , \g[17][51] , \g[17][50] , \g[17][49] , \g[17][48] , 
        \g[17][47] , \g[17][46] , \g[17][45] , \g[17][44] , \g[17][43] , 
        \g[17][42] , \g[17][41] , \g[17][40] , \g[17][39] , \g[17][38] , 
        \g[17][37] , \g[17][36] , \g[17][35] , \g[17][34] , \g[17][33] , 
        \g[17][32] , \g[17][31] , \g[17][30] , \g[17][29] , \g[17][28] , 
        \g[17][27] , \g[17][26] , \g[17][25] , \g[17][24] , \g[17][23] , 
        \g[17][22] , \g[17][21] , \g[17][20] , \g[17][19] , \g[17][18] , 
        \g[17][17] , \g[17][16] , \g[17][15] , \g[17][14] , \g[17][13] , 
        \g[17][12] , \g[17][11] , \g[17][10] , \g[17][9] , \g[17][8] , 
        \g[17][7] , \g[17][6] , \g[17][5] , \g[17][4] , \g[17][3] , \g[17][2] , 
        \g[17][1] , \g[17][0] }), .cout({\g[38][63] , \g[38][62] , \g[38][61] , 
        \g[38][60] , \g[38][59] , \g[38][58] , \g[38][57] , \g[38][56] , 
        \g[38][55] , \g[38][54] , \g[38][53] , \g[38][52] , \g[38][51] , 
        \g[38][50] , \g[38][49] , \g[38][48] , \g[38][47] , \g[38][46] , 
        \g[38][45] , \g[38][44] , \g[38][43] , \g[38][42] , \g[38][41] , 
        \g[38][40] , \g[38][39] , \g[38][38] , \g[38][37] , \g[38][36] , 
        \g[38][35] , \g[38][34] , \g[38][33] , \g[38][32] , \g[38][31] , 
        \g[38][30] , \g[38][29] , \g[38][28] , \g[38][27] , \g[38][26] , 
        \g[38][25] , \g[38][24] , \g[38][23] , \g[38][22] , \g[38][21] , 
        \g[38][20] , \g[38][19] , \g[38][18] , \g[38][17] , \g[38][16] , 
        \g[38][15] , \g[38][14] , \g[38][13] , \g[38][12] , \g[38][11] , 
        \g[38][10] , \g[38][9] , \g[38][8] , \g[38][7] , \g[38][6] , 
        \g[38][5] , \g[38][4] , \g[38][3] , \g[38][2] , \g[38][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  FullAdder_44 \level1[18].x6  ( .a({n453, n457, n462, n469, n474, n480, n485, 
        n490, n495, n500, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n457, n463, 
        n472, n477, n481, n487, n491, n497, n502, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n461, n465, n473, n478, n483, n489, n493, n498, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[18][63] , 
        \g[18][62] , \g[18][61] , \g[18][60] , \g[18][59] , \g[18][58] , 
        \g[18][57] , \g[18][56] , \g[18][55] , \g[18][54] , \g[18][53] , 
        \g[18][52] , \g[18][51] , \g[18][50] , \g[18][49] , \g[18][48] , 
        \g[18][47] , \g[18][46] , \g[18][45] , \g[18][44] , \g[18][43] , 
        \g[18][42] , \g[18][41] , \g[18][40] , \g[18][39] , \g[18][38] , 
        \g[18][37] , \g[18][36] , \g[18][35] , \g[18][34] , \g[18][33] , 
        \g[18][32] , \g[18][31] , \g[18][30] , \g[18][29] , \g[18][28] , 
        \g[18][27] , \g[18][26] , \g[18][25] , \g[18][24] , \g[18][23] , 
        \g[18][22] , \g[18][21] , \g[18][20] , \g[18][19] , \g[18][18] , 
        \g[18][17] , \g[18][16] , \g[18][15] , \g[18][14] , \g[18][13] , 
        \g[18][12] , \g[18][11] , \g[18][10] , \g[18][9] , \g[18][8] , 
        \g[18][7] , \g[18][6] , \g[18][5] , \g[18][4] , \g[18][3] , \g[18][2] , 
        \g[18][1] , \g[18][0] }), .cout({\g[39][63] , \g[39][62] , \g[39][61] , 
        \g[39][60] , \g[39][59] , \g[39][58] , \g[39][57] , \g[39][56] , 
        \g[39][55] , \g[39][54] , \g[39][53] , \g[39][52] , \g[39][51] , 
        \g[39][50] , \g[39][49] , \g[39][48] , \g[39][47] , \g[39][46] , 
        \g[39][45] , \g[39][44] , \g[39][43] , \g[39][42] , \g[39][41] , 
        \g[39][40] , \g[39][39] , \g[39][38] , \g[39][37] , \g[39][36] , 
        \g[39][35] , \g[39][34] , \g[39][33] , \g[39][32] , \g[39][31] , 
        \g[39][30] , \g[39][29] , \g[39][28] , \g[39][27] , \g[39][26] , 
        \g[39][25] , \g[39][24] , \g[39][23] , \g[39][22] , \g[39][21] , 
        \g[39][20] , \g[39][19] , \g[39][18] , \g[39][17] , \g[39][16] , 
        \g[39][15] , \g[39][14] , \g[39][13] , \g[39][12] , \g[39][11] , 
        \g[39][10] , \g[39][9] , \g[39][8] , \g[39][7] , \g[39][6] , 
        \g[39][5] , \g[39][4] , \g[39][3] , \g[39][2] , \g[39][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  FullAdder_43 \level1[19].x6  ( .a({n470, n474, n480, n486, n489, n494, n499, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n474, n482, 
        n487, n491, n497, n502, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n479, n483, n488, n493, n498, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[19][63] , 
        \g[19][62] , \g[19][61] , \g[19][60] , \g[19][59] , \g[19][58] , 
        \g[19][57] , \g[19][56] , \g[19][55] , \g[19][54] , \g[19][53] , 
        \g[19][52] , \g[19][51] , \g[19][50] , \g[19][49] , \g[19][48] , 
        \g[19][47] , \g[19][46] , \g[19][45] , \g[19][44] , \g[19][43] , 
        \g[19][42] , \g[19][41] , \g[19][40] , \g[19][39] , \g[19][38] , 
        \g[19][37] , \g[19][36] , \g[19][35] , \g[19][34] , \g[19][33] , 
        \g[19][32] , \g[19][31] , \g[19][30] , \g[19][29] , \g[19][28] , 
        \g[19][27] , \g[19][26] , \g[19][25] , \g[19][24] , \g[19][23] , 
        \g[19][22] , \g[19][21] , \g[19][20] , \g[19][19] , \g[19][18] , 
        \g[19][17] , \g[19][16] , \g[19][15] , \g[19][14] , \g[19][13] , 
        \g[19][12] , \g[19][11] , \g[19][10] , \g[19][9] , \g[19][8] , 
        \g[19][7] , \g[19][6] , \g[19][5] , \g[19][4] , \g[19][3] , \g[19][2] , 
        \g[19][1] , \g[19][0] }), .cout({\g[40][63] , \g[40][62] , \g[40][61] , 
        \g[40][60] , \g[40][59] , \g[40][58] , \g[40][57] , \g[40][56] , 
        \g[40][55] , \g[40][54] , \g[40][53] , \g[40][52] , \g[40][51] , 
        \g[40][50] , \g[40][49] , \g[40][48] , \g[40][47] , \g[40][46] , 
        \g[40][45] , \g[40][44] , \g[40][43] , \g[40][42] , \g[40][41] , 
        \g[40][40] , \g[40][39] , \g[40][38] , \g[40][37] , \g[40][36] , 
        \g[40][35] , \g[40][34] , \g[40][33] , \g[40][32] , \g[40][31] , 
        \g[40][30] , \g[40][29] , \g[40][28] , \g[40][27] , \g[40][26] , 
        \g[40][25] , \g[40][24] , \g[40][23] , \g[40][22] , \g[40][21] , 
        \g[40][20] , \g[40][19] , \g[40][18] , \g[40][17] , \g[40][16] , 
        \g[40][15] , \g[40][14] , \g[40][13] , \g[40][12] , \g[40][11] , 
        \g[40][10] , \g[40][9] , \g[40][8] , \g[40][7] , \g[40][6] , 
        \g[40][5] , \g[40][4] , \g[40][3] , \g[40][2] , \g[40][1] , 
        SYNOPSYS_UNCONNECTED__19}) );
  FullAdder_42 \level1[20].x6  ( .a({n484, n490, n495, n500, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n489, n497, 
        n502, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .cin({n494, n498, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({\g[20][63] , 
        \g[20][62] , \g[20][61] , \g[20][60] , \g[20][59] , \g[20][58] , 
        \g[20][57] , \g[20][56] , \g[20][55] , \g[20][54] , \g[20][53] , 
        \g[20][52] , \g[20][51] , \g[20][50] , \g[20][49] , \g[20][48] , 
        \g[20][47] , \g[20][46] , \g[20][45] , \g[20][44] , \g[20][43] , 
        \g[20][42] , \g[20][41] , \g[20][40] , \g[20][39] , \g[20][38] , 
        \g[20][37] , \g[20][36] , \g[20][35] , \g[20][34] , \g[20][33] , 
        \g[20][32] , \g[20][31] , \g[20][30] , \g[20][29] , \g[20][28] , 
        \g[20][27] , \g[20][26] , \g[20][25] , \g[20][24] , \g[20][23] , 
        \g[20][22] , \g[20][21] , \g[20][20] , \g[20][19] , \g[20][18] , 
        \g[20][17] , \g[20][16] , \g[20][15] , \g[20][14] , \g[20][13] , 
        \g[20][12] , \g[20][11] , \g[20][10] , \g[20][9] , \g[20][8] , 
        \g[20][7] , \g[20][6] , \g[20][5] , \g[20][4] , \g[20][3] , \g[20][2] , 
        \g[20][1] , \g[20][0] }), .cout({\g[41][63] , \g[41][62] , \g[41][61] , 
        \g[41][60] , \g[41][59] , \g[41][58] , \g[41][57] , \g[41][56] , 
        \g[41][55] , \g[41][54] , \g[41][53] , \g[41][52] , \g[41][51] , 
        \g[41][50] , \g[41][49] , \g[41][48] , \g[41][47] , \g[41][46] , 
        \g[41][45] , \g[41][44] , \g[41][43] , \g[41][42] , \g[41][41] , 
        \g[41][40] , \g[41][39] , \g[41][38] , \g[41][37] , \g[41][36] , 
        \g[41][35] , \g[41][34] , \g[41][33] , \g[41][32] , \g[41][31] , 
        \g[41][30] , \g[41][29] , \g[41][28] , \g[41][27] , \g[41][26] , 
        \g[41][25] , \g[41][24] , \g[41][23] , \g[41][22] , \g[41][21] , 
        \g[41][20] , \g[41][19] , \g[41][18] , \g[41][17] , \g[41][16] , 
        \g[41][15] , \g[41][14] , \g[41][13] , \g[41][12] , \g[41][11] , 
        \g[41][10] , \g[41][9] , \g[41][8] , \g[41][7] , \g[41][6] , 
        \g[41][5] , \g[41][4] , \g[41][3] , \g[41][2] , \g[41][1] , 
        SYNOPSYS_UNCONNECTED__20}) );
  FullAdder_41 \level2[0].x5  ( .a({\g[0][63] , \g[0][62] , \g[0][61] , 
        \g[0][60] , \g[0][59] , \g[0][58] , \g[0][57] , \g[0][56] , \g[0][55] , 
        \g[0][54] , \g[0][53] , \g[0][52] , \g[0][51] , \g[0][50] , \g[0][49] , 
        \g[0][48] , \g[0][47] , \g[0][46] , \g[0][45] , \g[0][44] , \g[0][43] , 
        \g[0][42] , \g[0][41] , \g[0][40] , \g[0][39] , \g[0][38] , \g[0][37] , 
        \g[0][36] , \g[0][35] , \g[0][34] , \g[0][33] , \g[0][32] , \g[0][31] , 
        \g[0][30] , \g[0][29] , \g[0][28] , \g[0][27] , \g[0][26] , \g[0][25] , 
        \g[0][24] , \g[0][23] , \g[0][22] , \g[0][21] , \g[0][20] , \g[0][19] , 
        \g[0][18] , \g[0][17] , \g[0][16] , \g[0][15] , \g[0][14] , \g[0][13] , 
        \g[0][12] , \g[0][11] , \g[0][10] , \g[0][9] , \g[0][8] , \g[0][7] , 
        \g[0][6] , \g[0][5] , \g[0][4] , \g[0][3] , \g[0][2] , \g[0][1] , 
        \g[0][0] }), .b({\g[1][63] , \g[1][62] , \g[1][61] , \g[1][60] , 
        \g[1][59] , \g[1][58] , \g[1][57] , \g[1][56] , \g[1][55] , \g[1][54] , 
        \g[1][53] , \g[1][52] , \g[1][51] , \g[1][50] , \g[1][49] , \g[1][48] , 
        \g[1][47] , \g[1][46] , \g[1][45] , \g[1][44] , \g[1][43] , \g[1][42] , 
        \g[1][41] , \g[1][40] , \g[1][39] , \g[1][38] , \g[1][37] , \g[1][36] , 
        \g[1][35] , \g[1][34] , \g[1][33] , \g[1][32] , \g[1][31] , \g[1][30] , 
        \g[1][29] , \g[1][28] , \g[1][27] , \g[1][26] , \g[1][25] , \g[1][24] , 
        \g[1][23] , \g[1][22] , \g[1][21] , \g[1][20] , \g[1][19] , \g[1][18] , 
        \g[1][17] , \g[1][16] , \g[1][15] , \g[1][14] , \g[1][13] , \g[1][12] , 
        \g[1][11] , \g[1][10] , \g[1][9] , \g[1][8] , \g[1][7] , \g[1][6] , 
        \g[1][5] , \g[1][4] , \g[1][3] , \g[1][2] , \g[1][1] , \g[1][0] }), 
        .cin({\g[2][63] , \g[2][62] , \g[2][61] , \g[2][60] , \g[2][59] , 
        \g[2][58] , \g[2][57] , \g[2][56] , \g[2][55] , \g[2][54] , \g[2][53] , 
        \g[2][52] , \g[2][51] , \g[2][50] , \g[2][49] , \g[2][48] , \g[2][47] , 
        \g[2][46] , \g[2][45] , \g[2][44] , \g[2][43] , \g[2][42] , \g[2][41] , 
        \g[2][40] , \g[2][39] , \g[2][38] , \g[2][37] , \g[2][36] , \g[2][35] , 
        \g[2][34] , \g[2][33] , \g[2][32] , \g[2][31] , \g[2][30] , \g[2][29] , 
        \g[2][28] , \g[2][27] , \g[2][26] , \g[2][25] , \g[2][24] , \g[2][23] , 
        \g[2][22] , \g[2][21] , \g[2][20] , \g[2][19] , \g[2][18] , \g[2][17] , 
        \g[2][16] , \g[2][15] , \g[2][14] , \g[2][13] , \g[2][12] , \g[2][11] , 
        \g[2][10] , \g[2][9] , \g[2][8] , \g[2][7] , \g[2][6] , \g[2][5] , 
        \g[2][4] , \g[2][3] , \g[2][2] , \g[2][1] , \g[2][0] }), .sum({
        \g2[0][63] , \g2[0][62] , \g2[0][61] , \g2[0][60] , \g2[0][59] , 
        \g2[0][58] , \g2[0][57] , \g2[0][56] , \g2[0][55] , \g2[0][54] , 
        \g2[0][53] , \g2[0][52] , \g2[0][51] , \g2[0][50] , \g2[0][49] , 
        \g2[0][48] , \g2[0][47] , \g2[0][46] , \g2[0][45] , \g2[0][44] , 
        \g2[0][43] , \g2[0][42] , \g2[0][41] , \g2[0][40] , \g2[0][39] , 
        \g2[0][38] , \g2[0][37] , \g2[0][36] , \g2[0][35] , \g2[0][34] , 
        \g2[0][33] , \g2[0][32] , \g2[0][31] , \g2[0][30] , \g2[0][29] , 
        \g2[0][28] , \g2[0][27] , \g2[0][26] , \g2[0][25] , \g2[0][24] , 
        \g2[0][23] , \g2[0][22] , \g2[0][21] , \g2[0][20] , \g2[0][19] , 
        \g2[0][18] , \g2[0][17] , \g2[0][16] , \g2[0][15] , \g2[0][14] , 
        \g2[0][13] , \g2[0][12] , \g2[0][11] , \g2[0][10] , \g2[0][9] , 
        \g2[0][8] , \g2[0][7] , \g2[0][6] , \g2[0][5] , \g2[0][4] , \g2[0][3] , 
        \g2[0][2] , \g2[0][1] , \g2[0][0] }), .cout({\g2[14][63] , 
        \g2[14][62] , \g2[14][61] , \g2[14][60] , \g2[14][59] , \g2[14][58] , 
        \g2[14][57] , \g2[14][56] , \g2[14][55] , \g2[14][54] , \g2[14][53] , 
        \g2[14][52] , \g2[14][51] , \g2[14][50] , \g2[14][49] , \g2[14][48] , 
        \g2[14][47] , \g2[14][46] , \g2[14][45] , \g2[14][44] , \g2[14][43] , 
        \g2[14][42] , \g2[14][41] , \g2[14][40] , \g2[14][39] , \g2[14][38] , 
        \g2[14][37] , \g2[14][36] , \g2[14][35] , \g2[14][34] , \g2[14][33] , 
        \g2[14][32] , \g2[14][31] , \g2[14][30] , \g2[14][29] , \g2[14][28] , 
        \g2[14][27] , \g2[14][26] , \g2[14][25] , \g2[14][24] , \g2[14][23] , 
        \g2[14][22] , \g2[14][21] , \g2[14][20] , \g2[14][19] , \g2[14][18] , 
        \g2[14][17] , \g2[14][16] , \g2[14][15] , \g2[14][14] , \g2[14][13] , 
        \g2[14][12] , \g2[14][11] , \g2[14][10] , \g2[14][9] , \g2[14][8] , 
        \g2[14][7] , \g2[14][6] , \g2[14][5] , \g2[14][4] , \g2[14][3] , 
        \g2[14][2] , \g2[14][1] , SYNOPSYS_UNCONNECTED__21}) );
  FullAdder_40 \level2[1].x5  ( .a({\g[3][63] , \g[3][62] , \g[3][61] , 
        \g[3][60] , \g[3][59] , \g[3][58] , \g[3][57] , \g[3][56] , \g[3][55] , 
        \g[3][54] , \g[3][53] , \g[3][52] , \g[3][51] , \g[3][50] , \g[3][49] , 
        \g[3][48] , \g[3][47] , \g[3][46] , \g[3][45] , \g[3][44] , \g[3][43] , 
        \g[3][42] , \g[3][41] , \g[3][40] , \g[3][39] , \g[3][38] , \g[3][37] , 
        \g[3][36] , \g[3][35] , \g[3][34] , \g[3][33] , \g[3][32] , \g[3][31] , 
        \g[3][30] , \g[3][29] , \g[3][28] , \g[3][27] , \g[3][26] , \g[3][25] , 
        \g[3][24] , \g[3][23] , \g[3][22] , \g[3][21] , \g[3][20] , \g[3][19] , 
        \g[3][18] , \g[3][17] , \g[3][16] , \g[3][15] , \g[3][14] , \g[3][13] , 
        \g[3][12] , \g[3][11] , \g[3][10] , \g[3][9] , \g[3][8] , \g[3][7] , 
        \g[3][6] , \g[3][5] , \g[3][4] , \g[3][3] , \g[3][2] , \g[3][1] , 
        \g[3][0] }), .b({\g[4][63] , \g[4][62] , \g[4][61] , \g[4][60] , 
        \g[4][59] , \g[4][58] , \g[4][57] , \g[4][56] , \g[4][55] , \g[4][54] , 
        \g[4][53] , \g[4][52] , \g[4][51] , \g[4][50] , \g[4][49] , \g[4][48] , 
        \g[4][47] , \g[4][46] , \g[4][45] , \g[4][44] , \g[4][43] , \g[4][42] , 
        \g[4][41] , \g[4][40] , \g[4][39] , \g[4][38] , \g[4][37] , \g[4][36] , 
        \g[4][35] , \g[4][34] , \g[4][33] , \g[4][32] , \g[4][31] , \g[4][30] , 
        \g[4][29] , \g[4][28] , \g[4][27] , \g[4][26] , \g[4][25] , \g[4][24] , 
        \g[4][23] , \g[4][22] , \g[4][21] , \g[4][20] , \g[4][19] , \g[4][18] , 
        \g[4][17] , \g[4][16] , \g[4][15] , \g[4][14] , \g[4][13] , \g[4][12] , 
        \g[4][11] , \g[4][10] , \g[4][9] , \g[4][8] , \g[4][7] , \g[4][6] , 
        \g[4][5] , \g[4][4] , \g[4][3] , \g[4][2] , \g[4][1] , \g[4][0] }), 
        .cin({\g[5][63] , \g[5][62] , \g[5][61] , \g[5][60] , \g[5][59] , 
        \g[5][58] , \g[5][57] , \g[5][56] , \g[5][55] , \g[5][54] , \g[5][53] , 
        \g[5][52] , \g[5][51] , \g[5][50] , \g[5][49] , \g[5][48] , \g[5][47] , 
        \g[5][46] , \g[5][45] , \g[5][44] , \g[5][43] , \g[5][42] , \g[5][41] , 
        \g[5][40] , \g[5][39] , \g[5][38] , \g[5][37] , \g[5][36] , \g[5][35] , 
        \g[5][34] , \g[5][33] , \g[5][32] , \g[5][31] , \g[5][30] , \g[5][29] , 
        \g[5][28] , \g[5][27] , \g[5][26] , \g[5][25] , \g[5][24] , \g[5][23] , 
        \g[5][22] , \g[5][21] , \g[5][20] , \g[5][19] , \g[5][18] , \g[5][17] , 
        \g[5][16] , \g[5][15] , \g[5][14] , \g[5][13] , \g[5][12] , \g[5][11] , 
        \g[5][10] , \g[5][9] , \g[5][8] , \g[5][7] , \g[5][6] , \g[5][5] , 
        \g[5][4] , \g[5][3] , \g[5][2] , \g[5][1] , \g[5][0] }), .sum({
        \g2[1][63] , \g2[1][62] , \g2[1][61] , \g2[1][60] , \g2[1][59] , 
        \g2[1][58] , \g2[1][57] , \g2[1][56] , \g2[1][55] , \g2[1][54] , 
        \g2[1][53] , \g2[1][52] , \g2[1][51] , \g2[1][50] , \g2[1][49] , 
        \g2[1][48] , \g2[1][47] , \g2[1][46] , \g2[1][45] , \g2[1][44] , 
        \g2[1][43] , \g2[1][42] , \g2[1][41] , \g2[1][40] , \g2[1][39] , 
        \g2[1][38] , \g2[1][37] , \g2[1][36] , \g2[1][35] , \g2[1][34] , 
        \g2[1][33] , \g2[1][32] , \g2[1][31] , \g2[1][30] , \g2[1][29] , 
        \g2[1][28] , \g2[1][27] , \g2[1][26] , \g2[1][25] , \g2[1][24] , 
        \g2[1][23] , \g2[1][22] , \g2[1][21] , \g2[1][20] , \g2[1][19] , 
        \g2[1][18] , \g2[1][17] , \g2[1][16] , \g2[1][15] , \g2[1][14] , 
        \g2[1][13] , \g2[1][12] , \g2[1][11] , \g2[1][10] , \g2[1][9] , 
        \g2[1][8] , \g2[1][7] , \g2[1][6] , \g2[1][5] , \g2[1][4] , \g2[1][3] , 
        \g2[1][2] , \g2[1][1] , \g2[1][0] }), .cout({\g2[15][63] , 
        \g2[15][62] , \g2[15][61] , \g2[15][60] , \g2[15][59] , \g2[15][58] , 
        \g2[15][57] , \g2[15][56] , \g2[15][55] , \g2[15][54] , \g2[15][53] , 
        \g2[15][52] , \g2[15][51] , \g2[15][50] , \g2[15][49] , \g2[15][48] , 
        \g2[15][47] , \g2[15][46] , \g2[15][45] , \g2[15][44] , \g2[15][43] , 
        \g2[15][42] , \g2[15][41] , \g2[15][40] , \g2[15][39] , \g2[15][38] , 
        \g2[15][37] , \g2[15][36] , \g2[15][35] , \g2[15][34] , \g2[15][33] , 
        \g2[15][32] , \g2[15][31] , \g2[15][30] , \g2[15][29] , \g2[15][28] , 
        \g2[15][27] , \g2[15][26] , \g2[15][25] , \g2[15][24] , \g2[15][23] , 
        \g2[15][22] , \g2[15][21] , \g2[15][20] , \g2[15][19] , \g2[15][18] , 
        \g2[15][17] , \g2[15][16] , \g2[15][15] , \g2[15][14] , \g2[15][13] , 
        \g2[15][12] , \g2[15][11] , \g2[15][10] , \g2[15][9] , \g2[15][8] , 
        \g2[15][7] , \g2[15][6] , \g2[15][5] , \g2[15][4] , \g2[15][3] , 
        \g2[15][2] , \g2[15][1] , SYNOPSYS_UNCONNECTED__22}) );
  FullAdder_39 \level2[2].x5  ( .a({\g[6][63] , \g[6][62] , \g[6][61] , 
        \g[6][60] , \g[6][59] , \g[6][58] , \g[6][57] , \g[6][56] , \g[6][55] , 
        \g[6][54] , \g[6][53] , \g[6][52] , \g[6][51] , \g[6][50] , \g[6][49] , 
        \g[6][48] , \g[6][47] , \g[6][46] , \g[6][45] , \g[6][44] , \g[6][43] , 
        \g[6][42] , \g[6][41] , \g[6][40] , \g[6][39] , \g[6][38] , \g[6][37] , 
        \g[6][36] , \g[6][35] , \g[6][34] , \g[6][33] , \g[6][32] , \g[6][31] , 
        \g[6][30] , \g[6][29] , \g[6][28] , \g[6][27] , \g[6][26] , \g[6][25] , 
        \g[6][24] , \g[6][23] , \g[6][22] , \g[6][21] , \g[6][20] , \g[6][19] , 
        \g[6][18] , \g[6][17] , \g[6][16] , \g[6][15] , \g[6][14] , \g[6][13] , 
        \g[6][12] , \g[6][11] , \g[6][10] , \g[6][9] , \g[6][8] , \g[6][7] , 
        \g[6][6] , \g[6][5] , \g[6][4] , \g[6][3] , \g[6][2] , \g[6][1] , 
        \g[6][0] }), .b({\g[7][63] , \g[7][62] , \g[7][61] , \g[7][60] , 
        \g[7][59] , \g[7][58] , \g[7][57] , \g[7][56] , \g[7][55] , \g[7][54] , 
        \g[7][53] , \g[7][52] , \g[7][51] , \g[7][50] , \g[7][49] , \g[7][48] , 
        \g[7][47] , \g[7][46] , \g[7][45] , \g[7][44] , \g[7][43] , \g[7][42] , 
        \g[7][41] , \g[7][40] , \g[7][39] , \g[7][38] , \g[7][37] , \g[7][36] , 
        \g[7][35] , \g[7][34] , \g[7][33] , \g[7][32] , \g[7][31] , \g[7][30] , 
        \g[7][29] , \g[7][28] , \g[7][27] , \g[7][26] , \g[7][25] , \g[7][24] , 
        \g[7][23] , \g[7][22] , \g[7][21] , \g[7][20] , \g[7][19] , \g[7][18] , 
        \g[7][17] , \g[7][16] , \g[7][15] , \g[7][14] , \g[7][13] , \g[7][12] , 
        \g[7][11] , \g[7][10] , \g[7][9] , \g[7][8] , \g[7][7] , \g[7][6] , 
        \g[7][5] , \g[7][4] , \g[7][3] , \g[7][2] , \g[7][1] , \g[7][0] }), 
        .cin({\g[8][63] , \g[8][62] , \g[8][61] , \g[8][60] , \g[8][59] , 
        \g[8][58] , \g[8][57] , \g[8][56] , \g[8][55] , \g[8][54] , \g[8][53] , 
        \g[8][52] , \g[8][51] , \g[8][50] , \g[8][49] , \g[8][48] , \g[8][47] , 
        \g[8][46] , \g[8][45] , \g[8][44] , \g[8][43] , \g[8][42] , \g[8][41] , 
        \g[8][40] , \g[8][39] , \g[8][38] , \g[8][37] , \g[8][36] , \g[8][35] , 
        \g[8][34] , \g[8][33] , \g[8][32] , \g[8][31] , \g[8][30] , \g[8][29] , 
        \g[8][28] , \g[8][27] , \g[8][26] , \g[8][25] , \g[8][24] , \g[8][23] , 
        \g[8][22] , \g[8][21] , \g[8][20] , \g[8][19] , \g[8][18] , \g[8][17] , 
        \g[8][16] , \g[8][15] , \g[8][14] , \g[8][13] , \g[8][12] , \g[8][11] , 
        \g[8][10] , \g[8][9] , \g[8][8] , \g[8][7] , \g[8][6] , \g[8][5] , 
        \g[8][4] , \g[8][3] , \g[8][2] , \g[8][1] , \g[8][0] }), .sum({
        \g2[2][63] , \g2[2][62] , \g2[2][61] , \g2[2][60] , \g2[2][59] , 
        \g2[2][58] , \g2[2][57] , \g2[2][56] , \g2[2][55] , \g2[2][54] , 
        \g2[2][53] , \g2[2][52] , \g2[2][51] , \g2[2][50] , \g2[2][49] , 
        \g2[2][48] , \g2[2][47] , \g2[2][46] , \g2[2][45] , \g2[2][44] , 
        \g2[2][43] , \g2[2][42] , \g2[2][41] , \g2[2][40] , \g2[2][39] , 
        \g2[2][38] , \g2[2][37] , \g2[2][36] , \g2[2][35] , \g2[2][34] , 
        \g2[2][33] , \g2[2][32] , \g2[2][31] , \g2[2][30] , \g2[2][29] , 
        \g2[2][28] , \g2[2][27] , \g2[2][26] , \g2[2][25] , \g2[2][24] , 
        \g2[2][23] , \g2[2][22] , \g2[2][21] , \g2[2][20] , \g2[2][19] , 
        \g2[2][18] , \g2[2][17] , \g2[2][16] , \g2[2][15] , \g2[2][14] , 
        \g2[2][13] , \g2[2][12] , \g2[2][11] , \g2[2][10] , \g2[2][9] , 
        \g2[2][8] , \g2[2][7] , \g2[2][6] , \g2[2][5] , \g2[2][4] , \g2[2][3] , 
        \g2[2][2] , \g2[2][1] , \g2[2][0] }), .cout({\g2[16][63] , 
        \g2[16][62] , \g2[16][61] , \g2[16][60] , \g2[16][59] , \g2[16][58] , 
        \g2[16][57] , \g2[16][56] , \g2[16][55] , \g2[16][54] , \g2[16][53] , 
        \g2[16][52] , \g2[16][51] , \g2[16][50] , \g2[16][49] , \g2[16][48] , 
        \g2[16][47] , \g2[16][46] , \g2[16][45] , \g2[16][44] , \g2[16][43] , 
        \g2[16][42] , \g2[16][41] , \g2[16][40] , \g2[16][39] , \g2[16][38] , 
        \g2[16][37] , \g2[16][36] , \g2[16][35] , \g2[16][34] , \g2[16][33] , 
        \g2[16][32] , \g2[16][31] , \g2[16][30] , \g2[16][29] , \g2[16][28] , 
        \g2[16][27] , \g2[16][26] , \g2[16][25] , \g2[16][24] , \g2[16][23] , 
        \g2[16][22] , \g2[16][21] , \g2[16][20] , \g2[16][19] , \g2[16][18] , 
        \g2[16][17] , \g2[16][16] , \g2[16][15] , \g2[16][14] , \g2[16][13] , 
        \g2[16][12] , \g2[16][11] , \g2[16][10] , \g2[16][9] , \g2[16][8] , 
        \g2[16][7] , \g2[16][6] , \g2[16][5] , \g2[16][4] , \g2[16][3] , 
        \g2[16][2] , \g2[16][1] , SYNOPSYS_UNCONNECTED__23}) );
  FullAdder_38 \level2[3].x5  ( .a({\g[9][63] , \g[9][62] , \g[9][61] , 
        \g[9][60] , \g[9][59] , \g[9][58] , \g[9][57] , \g[9][56] , \g[9][55] , 
        \g[9][54] , \g[9][53] , \g[9][52] , \g[9][51] , \g[9][50] , \g[9][49] , 
        \g[9][48] , \g[9][47] , \g[9][46] , \g[9][45] , \g[9][44] , \g[9][43] , 
        \g[9][42] , \g[9][41] , \g[9][40] , \g[9][39] , \g[9][38] , \g[9][37] , 
        \g[9][36] , \g[9][35] , \g[9][34] , \g[9][33] , \g[9][32] , \g[9][31] , 
        \g[9][30] , \g[9][29] , \g[9][28] , \g[9][27] , \g[9][26] , \g[9][25] , 
        \g[9][24] , \g[9][23] , \g[9][22] , \g[9][21] , \g[9][20] , \g[9][19] , 
        \g[9][18] , \g[9][17] , \g[9][16] , \g[9][15] , \g[9][14] , \g[9][13] , 
        \g[9][12] , \g[9][11] , \g[9][10] , \g[9][9] , \g[9][8] , \g[9][7] , 
        \g[9][6] , \g[9][5] , \g[9][4] , \g[9][3] , \g[9][2] , \g[9][1] , 
        \g[9][0] }), .b({\g[10][63] , \g[10][62] , \g[10][61] , \g[10][60] , 
        \g[10][59] , \g[10][58] , \g[10][57] , \g[10][56] , \g[10][55] , 
        \g[10][54] , \g[10][53] , \g[10][52] , \g[10][51] , \g[10][50] , 
        \g[10][49] , \g[10][48] , \g[10][47] , \g[10][46] , \g[10][45] , 
        \g[10][44] , \g[10][43] , \g[10][42] , \g[10][41] , \g[10][40] , 
        \g[10][39] , \g[10][38] , \g[10][37] , \g[10][36] , \g[10][35] , 
        \g[10][34] , \g[10][33] , \g[10][32] , \g[10][31] , \g[10][30] , 
        \g[10][29] , \g[10][28] , \g[10][27] , \g[10][26] , \g[10][25] , 
        \g[10][24] , \g[10][23] , \g[10][22] , \g[10][21] , \g[10][20] , 
        \g[10][19] , \g[10][18] , \g[10][17] , \g[10][16] , \g[10][15] , 
        \g[10][14] , \g[10][13] , \g[10][12] , \g[10][11] , \g[10][10] , 
        \g[10][9] , \g[10][8] , \g[10][7] , \g[10][6] , \g[10][5] , \g[10][4] , 
        \g[10][3] , \g[10][2] , \g[10][1] , \g[10][0] }), .cin({\g[11][63] , 
        \g[11][62] , \g[11][61] , \g[11][60] , \g[11][59] , \g[11][58] , 
        \g[11][57] , \g[11][56] , \g[11][55] , \g[11][54] , \g[11][53] , 
        \g[11][52] , \g[11][51] , \g[11][50] , \g[11][49] , \g[11][48] , 
        \g[11][47] , \g[11][46] , \g[11][45] , \g[11][44] , \g[11][43] , 
        \g[11][42] , \g[11][41] , \g[11][40] , \g[11][39] , \g[11][38] , 
        \g[11][37] , \g[11][36] , \g[11][35] , \g[11][34] , \g[11][33] , 
        \g[11][32] , \g[11][31] , \g[11][30] , \g[11][29] , \g[11][28] , 
        \g[11][27] , \g[11][26] , \g[11][25] , \g[11][24] , \g[11][23] , 
        \g[11][22] , \g[11][21] , \g[11][20] , \g[11][19] , \g[11][18] , 
        \g[11][17] , \g[11][16] , \g[11][15] , \g[11][14] , \g[11][13] , 
        \g[11][12] , \g[11][11] , \g[11][10] , \g[11][9] , \g[11][8] , 
        \g[11][7] , \g[11][6] , \g[11][5] , \g[11][4] , \g[11][3] , \g[11][2] , 
        \g[11][1] , \g[11][0] }), .sum({\g2[3][63] , \g2[3][62] , \g2[3][61] , 
        \g2[3][60] , \g2[3][59] , \g2[3][58] , \g2[3][57] , \g2[3][56] , 
        \g2[3][55] , \g2[3][54] , \g2[3][53] , \g2[3][52] , \g2[3][51] , 
        \g2[3][50] , \g2[3][49] , \g2[3][48] , \g2[3][47] , \g2[3][46] , 
        \g2[3][45] , \g2[3][44] , \g2[3][43] , \g2[3][42] , \g2[3][41] , 
        \g2[3][40] , \g2[3][39] , \g2[3][38] , \g2[3][37] , \g2[3][36] , 
        \g2[3][35] , \g2[3][34] , \g2[3][33] , \g2[3][32] , \g2[3][31] , 
        \g2[3][30] , \g2[3][29] , \g2[3][28] , \g2[3][27] , \g2[3][26] , 
        \g2[3][25] , \g2[3][24] , \g2[3][23] , \g2[3][22] , \g2[3][21] , 
        \g2[3][20] , \g2[3][19] , \g2[3][18] , \g2[3][17] , \g2[3][16] , 
        \g2[3][15] , \g2[3][14] , \g2[3][13] , \g2[3][12] , \g2[3][11] , 
        \g2[3][10] , \g2[3][9] , \g2[3][8] , \g2[3][7] , \g2[3][6] , 
        \g2[3][5] , \g2[3][4] , \g2[3][3] , \g2[3][2] , \g2[3][1] , \g2[3][0] }), .cout({\g2[17][63] , \g2[17][62] , \g2[17][61] , \g2[17][60] , \g2[17][59] , 
        \g2[17][58] , \g2[17][57] , \g2[17][56] , \g2[17][55] , \g2[17][54] , 
        \g2[17][53] , \g2[17][52] , \g2[17][51] , \g2[17][50] , \g2[17][49] , 
        \g2[17][48] , \g2[17][47] , \g2[17][46] , \g2[17][45] , \g2[17][44] , 
        \g2[17][43] , \g2[17][42] , \g2[17][41] , \g2[17][40] , \g2[17][39] , 
        \g2[17][38] , \g2[17][37] , \g2[17][36] , \g2[17][35] , \g2[17][34] , 
        \g2[17][33] , \g2[17][32] , \g2[17][31] , \g2[17][30] , \g2[17][29] , 
        \g2[17][28] , \g2[17][27] , \g2[17][26] , \g2[17][25] , \g2[17][24] , 
        \g2[17][23] , \g2[17][22] , \g2[17][21] , \g2[17][20] , \g2[17][19] , 
        \g2[17][18] , \g2[17][17] , \g2[17][16] , \g2[17][15] , \g2[17][14] , 
        \g2[17][13] , \g2[17][12] , \g2[17][11] , \g2[17][10] , \g2[17][9] , 
        \g2[17][8] , \g2[17][7] , \g2[17][6] , \g2[17][5] , \g2[17][4] , 
        \g2[17][3] , \g2[17][2] , \g2[17][1] , SYNOPSYS_UNCONNECTED__24}) );
  FullAdder_37 \level2[4].x5  ( .a({\g[12][63] , \g[12][62] , \g[12][61] , 
        \g[12][60] , \g[12][59] , \g[12][58] , \g[12][57] , \g[12][56] , 
        \g[12][55] , \g[12][54] , \g[12][53] , \g[12][52] , \g[12][51] , 
        \g[12][50] , \g[12][49] , \g[12][48] , \g[12][47] , \g[12][46] , 
        \g[12][45] , \g[12][44] , \g[12][43] , \g[12][42] , \g[12][41] , 
        \g[12][40] , \g[12][39] , \g[12][38] , \g[12][37] , \g[12][36] , 
        \g[12][35] , \g[12][34] , \g[12][33] , \g[12][32] , \g[12][31] , 
        \g[12][30] , \g[12][29] , \g[12][28] , \g[12][27] , \g[12][26] , 
        \g[12][25] , \g[12][24] , \g[12][23] , \g[12][22] , \g[12][21] , 
        \g[12][20] , \g[12][19] , \g[12][18] , \g[12][17] , \g[12][16] , 
        \g[12][15] , \g[12][14] , \g[12][13] , \g[12][12] , \g[12][11] , 
        \g[12][10] , \g[12][9] , \g[12][8] , \g[12][7] , \g[12][6] , 
        \g[12][5] , \g[12][4] , \g[12][3] , \g[12][2] , \g[12][1] , \g[12][0] }), .b({\g[13][63] , \g[13][62] , \g[13][61] , \g[13][60] , \g[13][59] , 
        \g[13][58] , \g[13][57] , \g[13][56] , \g[13][55] , \g[13][54] , 
        \g[13][53] , \g[13][52] , \g[13][51] , \g[13][50] , \g[13][49] , 
        \g[13][48] , \g[13][47] , \g[13][46] , \g[13][45] , \g[13][44] , 
        \g[13][43] , \g[13][42] , \g[13][41] , \g[13][40] , \g[13][39] , 
        \g[13][38] , \g[13][37] , \g[13][36] , \g[13][35] , \g[13][34] , 
        \g[13][33] , \g[13][32] , \g[13][31] , \g[13][30] , \g[13][29] , 
        \g[13][28] , \g[13][27] , \g[13][26] , \g[13][25] , \g[13][24] , 
        \g[13][23] , \g[13][22] , \g[13][21] , \g[13][20] , \g[13][19] , 
        \g[13][18] , \g[13][17] , \g[13][16] , \g[13][15] , \g[13][14] , 
        \g[13][13] , \g[13][12] , \g[13][11] , \g[13][10] , \g[13][9] , 
        \g[13][8] , \g[13][7] , \g[13][6] , \g[13][5] , \g[13][4] , \g[13][3] , 
        \g[13][2] , \g[13][1] , \g[13][0] }), .cin({\g[14][63] , \g[14][62] , 
        \g[14][61] , \g[14][60] , \g[14][59] , \g[14][58] , \g[14][57] , 
        \g[14][56] , \g[14][55] , \g[14][54] , \g[14][53] , \g[14][52] , 
        \g[14][51] , \g[14][50] , \g[14][49] , \g[14][48] , \g[14][47] , 
        \g[14][46] , \g[14][45] , \g[14][44] , \g[14][43] , \g[14][42] , 
        \g[14][41] , \g[14][40] , \g[14][39] , \g[14][38] , \g[14][37] , 
        \g[14][36] , \g[14][35] , \g[14][34] , \g[14][33] , \g[14][32] , 
        \g[14][31] , \g[14][30] , \g[14][29] , \g[14][28] , \g[14][27] , 
        \g[14][26] , \g[14][25] , \g[14][24] , \g[14][23] , \g[14][22] , 
        \g[14][21] , \g[14][20] , \g[14][19] , \g[14][18] , \g[14][17] , 
        \g[14][16] , \g[14][15] , \g[14][14] , \g[14][13] , \g[14][12] , 
        \g[14][11] , \g[14][10] , \g[14][9] , \g[14][8] , \g[14][7] , 
        \g[14][6] , \g[14][5] , \g[14][4] , \g[14][3] , \g[14][2] , \g[14][1] , 
        \g[14][0] }), .sum({\g2[4][63] , \g2[4][62] , \g2[4][61] , \g2[4][60] , 
        \g2[4][59] , \g2[4][58] , \g2[4][57] , \g2[4][56] , \g2[4][55] , 
        \g2[4][54] , \g2[4][53] , \g2[4][52] , \g2[4][51] , \g2[4][50] , 
        \g2[4][49] , \g2[4][48] , \g2[4][47] , \g2[4][46] , \g2[4][45] , 
        \g2[4][44] , \g2[4][43] , \g2[4][42] , \g2[4][41] , \g2[4][40] , 
        \g2[4][39] , \g2[4][38] , \g2[4][37] , \g2[4][36] , \g2[4][35] , 
        \g2[4][34] , \g2[4][33] , \g2[4][32] , \g2[4][31] , \g2[4][30] , 
        \g2[4][29] , \g2[4][28] , \g2[4][27] , \g2[4][26] , \g2[4][25] , 
        \g2[4][24] , \g2[4][23] , \g2[4][22] , \g2[4][21] , \g2[4][20] , 
        \g2[4][19] , \g2[4][18] , \g2[4][17] , \g2[4][16] , \g2[4][15] , 
        \g2[4][14] , \g2[4][13] , \g2[4][12] , \g2[4][11] , \g2[4][10] , 
        \g2[4][9] , \g2[4][8] , \g2[4][7] , \g2[4][6] , \g2[4][5] , \g2[4][4] , 
        \g2[4][3] , \g2[4][2] , \g2[4][1] , \g2[4][0] }), .cout({\g2[18][63] , 
        \g2[18][62] , \g2[18][61] , \g2[18][60] , \g2[18][59] , \g2[18][58] , 
        \g2[18][57] , \g2[18][56] , \g2[18][55] , \g2[18][54] , \g2[18][53] , 
        \g2[18][52] , \g2[18][51] , \g2[18][50] , \g2[18][49] , \g2[18][48] , 
        \g2[18][47] , \g2[18][46] , \g2[18][45] , \g2[18][44] , \g2[18][43] , 
        \g2[18][42] , \g2[18][41] , \g2[18][40] , \g2[18][39] , \g2[18][38] , 
        \g2[18][37] , \g2[18][36] , \g2[18][35] , \g2[18][34] , \g2[18][33] , 
        \g2[18][32] , \g2[18][31] , \g2[18][30] , \g2[18][29] , \g2[18][28] , 
        \g2[18][27] , \g2[18][26] , \g2[18][25] , \g2[18][24] , \g2[18][23] , 
        \g2[18][22] , \g2[18][21] , \g2[18][20] , \g2[18][19] , \g2[18][18] , 
        \g2[18][17] , \g2[18][16] , \g2[18][15] , \g2[18][14] , \g2[18][13] , 
        \g2[18][12] , \g2[18][11] , \g2[18][10] , \g2[18][9] , \g2[18][8] , 
        \g2[18][7] , \g2[18][6] , \g2[18][5] , \g2[18][4] , \g2[18][3] , 
        \g2[18][2] , \g2[18][1] , SYNOPSYS_UNCONNECTED__25}) );
  FullAdder_36 \level2[5].x5  ( .a({\g[15][63] , \g[15][62] , \g[15][61] , 
        \g[15][60] , \g[15][59] , \g[15][58] , \g[15][57] , \g[15][56] , 
        \g[15][55] , \g[15][54] , \g[15][53] , \g[15][52] , \g[15][51] , 
        \g[15][50] , \g[15][49] , \g[15][48] , \g[15][47] , \g[15][46] , 
        \g[15][45] , \g[15][44] , \g[15][43] , \g[15][42] , \g[15][41] , 
        \g[15][40] , \g[15][39] , \g[15][38] , \g[15][37] , \g[15][36] , 
        \g[15][35] , \g[15][34] , \g[15][33] , \g[15][32] , \g[15][31] , 
        \g[15][30] , \g[15][29] , \g[15][28] , \g[15][27] , \g[15][26] , 
        \g[15][25] , \g[15][24] , \g[15][23] , \g[15][22] , \g[15][21] , 
        \g[15][20] , \g[15][19] , \g[15][18] , \g[15][17] , \g[15][16] , 
        \g[15][15] , \g[15][14] , \g[15][13] , \g[15][12] , \g[15][11] , 
        \g[15][10] , \g[15][9] , \g[15][8] , \g[15][7] , \g[15][6] , 
        \g[15][5] , \g[15][4] , \g[15][3] , \g[15][2] , \g[15][1] , \g[15][0] }), .b({\g[16][63] , \g[16][62] , \g[16][61] , \g[16][60] , \g[16][59] , 
        \g[16][58] , \g[16][57] , \g[16][56] , \g[16][55] , \g[16][54] , 
        \g[16][53] , \g[16][52] , \g[16][51] , \g[16][50] , \g[16][49] , 
        \g[16][48] , \g[16][47] , \g[16][46] , \g[16][45] , \g[16][44] , 
        \g[16][43] , \g[16][42] , \g[16][41] , \g[16][40] , \g[16][39] , 
        \g[16][38] , \g[16][37] , \g[16][36] , \g[16][35] , \g[16][34] , 
        \g[16][33] , \g[16][32] , \g[16][31] , \g[16][30] , \g[16][29] , 
        \g[16][28] , \g[16][27] , \g[16][26] , \g[16][25] , \g[16][24] , 
        \g[16][23] , \g[16][22] , \g[16][21] , \g[16][20] , \g[16][19] , 
        \g[16][18] , \g[16][17] , \g[16][16] , \g[16][15] , \g[16][14] , 
        \g[16][13] , \g[16][12] , \g[16][11] , \g[16][10] , \g[16][9] , 
        \g[16][8] , \g[16][7] , \g[16][6] , \g[16][5] , \g[16][4] , \g[16][3] , 
        \g[16][2] , \g[16][1] , \g[16][0] }), .cin({\g[17][63] , \g[17][62] , 
        \g[17][61] , \g[17][60] , \g[17][59] , \g[17][58] , \g[17][57] , 
        \g[17][56] , \g[17][55] , \g[17][54] , \g[17][53] , \g[17][52] , 
        \g[17][51] , \g[17][50] , \g[17][49] , \g[17][48] , \g[17][47] , 
        \g[17][46] , \g[17][45] , \g[17][44] , \g[17][43] , \g[17][42] , 
        \g[17][41] , \g[17][40] , \g[17][39] , \g[17][38] , \g[17][37] , 
        \g[17][36] , \g[17][35] , \g[17][34] , \g[17][33] , \g[17][32] , 
        \g[17][31] , \g[17][30] , \g[17][29] , \g[17][28] , \g[17][27] , 
        \g[17][26] , \g[17][25] , \g[17][24] , \g[17][23] , \g[17][22] , 
        \g[17][21] , \g[17][20] , \g[17][19] , \g[17][18] , \g[17][17] , 
        \g[17][16] , \g[17][15] , \g[17][14] , \g[17][13] , \g[17][12] , 
        \g[17][11] , \g[17][10] , \g[17][9] , \g[17][8] , \g[17][7] , 
        \g[17][6] , \g[17][5] , \g[17][4] , \g[17][3] , \g[17][2] , \g[17][1] , 
        \g[17][0] }), .sum({\g2[5][63] , \g2[5][62] , \g2[5][61] , \g2[5][60] , 
        \g2[5][59] , \g2[5][58] , \g2[5][57] , \g2[5][56] , \g2[5][55] , 
        \g2[5][54] , \g2[5][53] , \g2[5][52] , \g2[5][51] , \g2[5][50] , 
        \g2[5][49] , \g2[5][48] , \g2[5][47] , \g2[5][46] , \g2[5][45] , 
        \g2[5][44] , \g2[5][43] , \g2[5][42] , \g2[5][41] , \g2[5][40] , 
        \g2[5][39] , \g2[5][38] , \g2[5][37] , \g2[5][36] , \g2[5][35] , 
        \g2[5][34] , \g2[5][33] , \g2[5][32] , \g2[5][31] , \g2[5][30] , 
        \g2[5][29] , \g2[5][28] , \g2[5][27] , \g2[5][26] , \g2[5][25] , 
        \g2[5][24] , \g2[5][23] , \g2[5][22] , \g2[5][21] , \g2[5][20] , 
        \g2[5][19] , \g2[5][18] , \g2[5][17] , \g2[5][16] , \g2[5][15] , 
        \g2[5][14] , \g2[5][13] , \g2[5][12] , \g2[5][11] , \g2[5][10] , 
        \g2[5][9] , \g2[5][8] , \g2[5][7] , \g2[5][6] , \g2[5][5] , \g2[5][4] , 
        \g2[5][3] , \g2[5][2] , \g2[5][1] , \g2[5][0] }), .cout({\g2[19][63] , 
        \g2[19][62] , \g2[19][61] , \g2[19][60] , \g2[19][59] , \g2[19][58] , 
        \g2[19][57] , \g2[19][56] , \g2[19][55] , \g2[19][54] , \g2[19][53] , 
        \g2[19][52] , \g2[19][51] , \g2[19][50] , \g2[19][49] , \g2[19][48] , 
        \g2[19][47] , \g2[19][46] , \g2[19][45] , \g2[19][44] , \g2[19][43] , 
        \g2[19][42] , \g2[19][41] , \g2[19][40] , \g2[19][39] , \g2[19][38] , 
        \g2[19][37] , \g2[19][36] , \g2[19][35] , \g2[19][34] , \g2[19][33] , 
        \g2[19][32] , \g2[19][31] , \g2[19][30] , \g2[19][29] , \g2[19][28] , 
        \g2[19][27] , \g2[19][26] , \g2[19][25] , \g2[19][24] , \g2[19][23] , 
        \g2[19][22] , \g2[19][21] , \g2[19][20] , \g2[19][19] , \g2[19][18] , 
        \g2[19][17] , \g2[19][16] , \g2[19][15] , \g2[19][14] , \g2[19][13] , 
        \g2[19][12] , \g2[19][11] , \g2[19][10] , \g2[19][9] , \g2[19][8] , 
        \g2[19][7] , \g2[19][6] , \g2[19][5] , \g2[19][4] , \g2[19][3] , 
        \g2[19][2] , \g2[19][1] , SYNOPSYS_UNCONNECTED__26}) );
  FullAdder_35 \level2[6].x5  ( .a({\g[18][63] , \g[18][62] , \g[18][61] , 
        \g[18][60] , \g[18][59] , \g[18][58] , \g[18][57] , \g[18][56] , 
        \g[18][55] , \g[18][54] , \g[18][53] , \g[18][52] , \g[18][51] , 
        \g[18][50] , \g[18][49] , \g[18][48] , \g[18][47] , \g[18][46] , 
        \g[18][45] , \g[18][44] , \g[18][43] , \g[18][42] , \g[18][41] , 
        \g[18][40] , \g[18][39] , \g[18][38] , \g[18][37] , \g[18][36] , 
        \g[18][35] , \g[18][34] , \g[18][33] , \g[18][32] , \g[18][31] , 
        \g[18][30] , \g[18][29] , \g[18][28] , \g[18][27] , \g[18][26] , 
        \g[18][25] , \g[18][24] , \g[18][23] , \g[18][22] , \g[18][21] , 
        \g[18][20] , \g[18][19] , \g[18][18] , \g[18][17] , \g[18][16] , 
        \g[18][15] , \g[18][14] , \g[18][13] , \g[18][12] , \g[18][11] , 
        \g[18][10] , \g[18][9] , \g[18][8] , \g[18][7] , \g[18][6] , 
        \g[18][5] , \g[18][4] , \g[18][3] , \g[18][2] , \g[18][1] , \g[18][0] }), .b({\g[19][63] , \g[19][62] , \g[19][61] , \g[19][60] , \g[19][59] , 
        \g[19][58] , \g[19][57] , \g[19][56] , \g[19][55] , \g[19][54] , 
        \g[19][53] , \g[19][52] , \g[19][51] , \g[19][50] , \g[19][49] , 
        \g[19][48] , \g[19][47] , \g[19][46] , \g[19][45] , \g[19][44] , 
        \g[19][43] , \g[19][42] , \g[19][41] , \g[19][40] , \g[19][39] , 
        \g[19][38] , \g[19][37] , \g[19][36] , \g[19][35] , \g[19][34] , 
        \g[19][33] , \g[19][32] , \g[19][31] , \g[19][30] , \g[19][29] , 
        \g[19][28] , \g[19][27] , \g[19][26] , \g[19][25] , \g[19][24] , 
        \g[19][23] , \g[19][22] , \g[19][21] , \g[19][20] , \g[19][19] , 
        \g[19][18] , \g[19][17] , \g[19][16] , \g[19][15] , \g[19][14] , 
        \g[19][13] , \g[19][12] , \g[19][11] , \g[19][10] , \g[19][9] , 
        \g[19][8] , \g[19][7] , \g[19][6] , \g[19][5] , \g[19][4] , \g[19][3] , 
        \g[19][2] , \g[19][1] , \g[19][0] }), .cin({\g[20][63] , \g[20][62] , 
        \g[20][61] , \g[20][60] , \g[20][59] , \g[20][58] , \g[20][57] , 
        \g[20][56] , \g[20][55] , \g[20][54] , \g[20][53] , \g[20][52] , 
        \g[20][51] , \g[20][50] , \g[20][49] , \g[20][48] , \g[20][47] , 
        \g[20][46] , \g[20][45] , \g[20][44] , \g[20][43] , \g[20][42] , 
        \g[20][41] , \g[20][40] , \g[20][39] , \g[20][38] , \g[20][37] , 
        \g[20][36] , \g[20][35] , \g[20][34] , \g[20][33] , \g[20][32] , 
        \g[20][31] , \g[20][30] , \g[20][29] , \g[20][28] , \g[20][27] , 
        \g[20][26] , \g[20][25] , \g[20][24] , \g[20][23] , \g[20][22] , 
        \g[20][21] , \g[20][20] , \g[20][19] , \g[20][18] , \g[20][17] , 
        \g[20][16] , \g[20][15] , \g[20][14] , \g[20][13] , \g[20][12] , 
        \g[20][11] , \g[20][10] , \g[20][9] , \g[20][8] , \g[20][7] , 
        \g[20][6] , \g[20][5] , \g[20][4] , \g[20][3] , \g[20][2] , \g[20][1] , 
        \g[20][0] }), .sum({\g2[6][63] , \g2[6][62] , \g2[6][61] , \g2[6][60] , 
        \g2[6][59] , \g2[6][58] , \g2[6][57] , \g2[6][56] , \g2[6][55] , 
        \g2[6][54] , \g2[6][53] , \g2[6][52] , \g2[6][51] , \g2[6][50] , 
        \g2[6][49] , \g2[6][48] , \g2[6][47] , \g2[6][46] , \g2[6][45] , 
        \g2[6][44] , \g2[6][43] , \g2[6][42] , \g2[6][41] , \g2[6][40] , 
        \g2[6][39] , \g2[6][38] , \g2[6][37] , \g2[6][36] , \g2[6][35] , 
        \g2[6][34] , \g2[6][33] , \g2[6][32] , \g2[6][31] , \g2[6][30] , 
        \g2[6][29] , \g2[6][28] , \g2[6][27] , \g2[6][26] , \g2[6][25] , 
        \g2[6][24] , \g2[6][23] , \g2[6][22] , \g2[6][21] , \g2[6][20] , 
        \g2[6][19] , \g2[6][18] , \g2[6][17] , \g2[6][16] , \g2[6][15] , 
        \g2[6][14] , \g2[6][13] , \g2[6][12] , \g2[6][11] , \g2[6][10] , 
        \g2[6][9] , \g2[6][8] , \g2[6][7] , \g2[6][6] , \g2[6][5] , \g2[6][4] , 
        \g2[6][3] , \g2[6][2] , \g2[6][1] , \g2[6][0] }), .cout({\g2[20][63] , 
        \g2[20][62] , \g2[20][61] , \g2[20][60] , \g2[20][59] , \g2[20][58] , 
        \g2[20][57] , \g2[20][56] , \g2[20][55] , \g2[20][54] , \g2[20][53] , 
        \g2[20][52] , \g2[20][51] , \g2[20][50] , \g2[20][49] , \g2[20][48] , 
        \g2[20][47] , \g2[20][46] , \g2[20][45] , \g2[20][44] , \g2[20][43] , 
        \g2[20][42] , \g2[20][41] , \g2[20][40] , \g2[20][39] , \g2[20][38] , 
        \g2[20][37] , \g2[20][36] , \g2[20][35] , \g2[20][34] , \g2[20][33] , 
        \g2[20][32] , \g2[20][31] , \g2[20][30] , \g2[20][29] , \g2[20][28] , 
        \g2[20][27] , \g2[20][26] , \g2[20][25] , \g2[20][24] , \g2[20][23] , 
        \g2[20][22] , \g2[20][21] , \g2[20][20] , \g2[20][19] , \g2[20][18] , 
        \g2[20][17] , \g2[20][16] , \g2[20][15] , \g2[20][14] , \g2[20][13] , 
        \g2[20][12] , \g2[20][11] , \g2[20][10] , \g2[20][9] , \g2[20][8] , 
        \g2[20][7] , \g2[20][6] , \g2[20][5] , \g2[20][4] , \g2[20][3] , 
        \g2[20][2] , \g2[20][1] , SYNOPSYS_UNCONNECTED__27}) );
  FullAdder_34 \level2[7].x5  ( .a({\g[21][63] , \g[21][62] , \g[21][61] , 
        \g[21][60] , \g[21][59] , \g[21][58] , \g[21][57] , \g[21][56] , 
        \g[21][55] , \g[21][54] , \g[21][53] , \g[21][52] , \g[21][51] , 
        \g[21][50] , \g[21][49] , \g[21][48] , \g[21][47] , \g[21][46] , 
        \g[21][45] , \g[21][44] , \g[21][43] , \g[21][42] , \g[21][41] , 
        \g[21][40] , \g[21][39] , \g[21][38] , \g[21][37] , \g[21][36] , 
        \g[21][35] , \g[21][34] , \g[21][33] , \g[21][32] , \g[21][31] , 
        \g[21][30] , \g[21][29] , \g[21][28] , \g[21][27] , \g[21][26] , 
        \g[21][25] , \g[21][24] , \g[21][23] , \g[21][22] , \g[21][21] , 
        \g[21][20] , \g[21][19] , \g[21][18] , \g[21][17] , \g[21][16] , 
        \g[21][15] , \g[21][14] , \g[21][13] , \g[21][12] , \g[21][11] , 
        \g[21][10] , \g[21][9] , \g[21][8] , \g[21][7] , \g[21][6] , 
        \g[21][5] , \g[21][4] , \g[21][3] , \g[21][2] , \g[21][1] , 1'b0}), 
        .b({\g[22][63] , \g[22][62] , \g[22][61] , \g[22][60] , \g[22][59] , 
        \g[22][58] , \g[22][57] , \g[22][56] , \g[22][55] , \g[22][54] , 
        \g[22][53] , \g[22][52] , \g[22][51] , \g[22][50] , \g[22][49] , 
        \g[22][48] , \g[22][47] , \g[22][46] , \g[22][45] , \g[22][44] , 
        \g[22][43] , \g[22][42] , \g[22][41] , \g[22][40] , \g[22][39] , 
        \g[22][38] , \g[22][37] , \g[22][36] , \g[22][35] , \g[22][34] , 
        \g[22][33] , \g[22][32] , \g[22][31] , \g[22][30] , \g[22][29] , 
        \g[22][28] , \g[22][27] , \g[22][26] , \g[22][25] , \g[22][24] , 
        \g[22][23] , \g[22][22] , \g[22][21] , \g[22][20] , \g[22][19] , 
        \g[22][18] , \g[22][17] , \g[22][16] , \g[22][15] , \g[22][14] , 
        \g[22][13] , \g[22][12] , \g[22][11] , \g[22][10] , \g[22][9] , 
        \g[22][8] , \g[22][7] , \g[22][6] , \g[22][5] , \g[22][4] , \g[22][3] , 
        \g[22][2] , \g[22][1] , 1'b0}), .cin({\g[23][63] , \g[23][62] , 
        \g[23][61] , \g[23][60] , \g[23][59] , \g[23][58] , \g[23][57] , 
        \g[23][56] , \g[23][55] , \g[23][54] , \g[23][53] , \g[23][52] , 
        \g[23][51] , \g[23][50] , \g[23][49] , \g[23][48] , \g[23][47] , 
        \g[23][46] , \g[23][45] , \g[23][44] , \g[23][43] , \g[23][42] , 
        \g[23][41] , \g[23][40] , \g[23][39] , \g[23][38] , \g[23][37] , 
        \g[23][36] , \g[23][35] , \g[23][34] , \g[23][33] , \g[23][32] , 
        \g[23][31] , \g[23][30] , \g[23][29] , \g[23][28] , \g[23][27] , 
        \g[23][26] , \g[23][25] , \g[23][24] , \g[23][23] , \g[23][22] , 
        \g[23][21] , \g[23][20] , \g[23][19] , \g[23][18] , \g[23][17] , 
        \g[23][16] , \g[23][15] , \g[23][14] , \g[23][13] , \g[23][12] , 
        \g[23][11] , \g[23][10] , \g[23][9] , \g[23][8] , \g[23][7] , 
        \g[23][6] , \g[23][5] , \g[23][4] , \g[23][3] , \g[23][2] , \g[23][1] , 
        1'b0}), .sum({\g2[7][63] , \g2[7][62] , \g2[7][61] , \g2[7][60] , 
        \g2[7][59] , \g2[7][58] , \g2[7][57] , \g2[7][56] , \g2[7][55] , 
        \g2[7][54] , \g2[7][53] , \g2[7][52] , \g2[7][51] , \g2[7][50] , 
        \g2[7][49] , \g2[7][48] , \g2[7][47] , \g2[7][46] , \g2[7][45] , 
        \g2[7][44] , \g2[7][43] , \g2[7][42] , \g2[7][41] , \g2[7][40] , 
        \g2[7][39] , \g2[7][38] , \g2[7][37] , \g2[7][36] , \g2[7][35] , 
        \g2[7][34] , \g2[7][33] , \g2[7][32] , \g2[7][31] , \g2[7][30] , 
        \g2[7][29] , \g2[7][28] , \g2[7][27] , \g2[7][26] , \g2[7][25] , 
        \g2[7][24] , \g2[7][23] , \g2[7][22] , \g2[7][21] , \g2[7][20] , 
        \g2[7][19] , \g2[7][18] , \g2[7][17] , \g2[7][16] , \g2[7][15] , 
        \g2[7][14] , \g2[7][13] , \g2[7][12] , \g2[7][11] , \g2[7][10] , 
        \g2[7][9] , \g2[7][8] , \g2[7][7] , \g2[7][6] , \g2[7][5] , \g2[7][4] , 
        \g2[7][3] , \g2[7][2] , \g2[7][1] , \g2[7][0] }), .cout({\g2[21][63] , 
        \g2[21][62] , \g2[21][61] , \g2[21][60] , \g2[21][59] , \g2[21][58] , 
        \g2[21][57] , \g2[21][56] , \g2[21][55] , \g2[21][54] , \g2[21][53] , 
        \g2[21][52] , \g2[21][51] , \g2[21][50] , \g2[21][49] , \g2[21][48] , 
        \g2[21][47] , \g2[21][46] , \g2[21][45] , \g2[21][44] , \g2[21][43] , 
        \g2[21][42] , \g2[21][41] , \g2[21][40] , \g2[21][39] , \g2[21][38] , 
        \g2[21][37] , \g2[21][36] , \g2[21][35] , \g2[21][34] , \g2[21][33] , 
        \g2[21][32] , \g2[21][31] , \g2[21][30] , \g2[21][29] , \g2[21][28] , 
        \g2[21][27] , \g2[21][26] , \g2[21][25] , \g2[21][24] , \g2[21][23] , 
        \g2[21][22] , \g2[21][21] , \g2[21][20] , \g2[21][19] , \g2[21][18] , 
        \g2[21][17] , \g2[21][16] , \g2[21][15] , \g2[21][14] , \g2[21][13] , 
        \g2[21][12] , \g2[21][11] , \g2[21][10] , \g2[21][9] , \g2[21][8] , 
        \g2[21][7] , \g2[21][6] , \g2[21][5] , \g2[21][4] , \g2[21][3] , 
        \g2[21][2] , \g2[21][1] , SYNOPSYS_UNCONNECTED__28}) );
  FullAdder_33 \level2[8].x5  ( .a({\g[24][63] , \g[24][62] , \g[24][61] , 
        \g[24][60] , \g[24][59] , \g[24][58] , \g[24][57] , \g[24][56] , 
        \g[24][55] , \g[24][54] , \g[24][53] , \g[24][52] , \g[24][51] , 
        \g[24][50] , \g[24][49] , \g[24][48] , \g[24][47] , \g[24][46] , 
        \g[24][45] , \g[24][44] , \g[24][43] , \g[24][42] , \g[24][41] , 
        \g[24][40] , \g[24][39] , \g[24][38] , \g[24][37] , \g[24][36] , 
        \g[24][35] , \g[24][34] , \g[24][33] , \g[24][32] , \g[24][31] , 
        \g[24][30] , \g[24][29] , \g[24][28] , \g[24][27] , \g[24][26] , 
        \g[24][25] , \g[24][24] , \g[24][23] , \g[24][22] , \g[24][21] , 
        \g[24][20] , \g[24][19] , \g[24][18] , \g[24][17] , \g[24][16] , 
        \g[24][15] , \g[24][14] , \g[24][13] , \g[24][12] , \g[24][11] , 
        \g[24][10] , \g[24][9] , \g[24][8] , \g[24][7] , \g[24][6] , 
        \g[24][5] , \g[24][4] , \g[24][3] , \g[24][2] , \g[24][1] , 1'b0}), 
        .b({\g[25][63] , \g[25][62] , \g[25][61] , \g[25][60] , \g[25][59] , 
        \g[25][58] , \g[25][57] , \g[25][56] , \g[25][55] , \g[25][54] , 
        \g[25][53] , \g[25][52] , \g[25][51] , \g[25][50] , \g[25][49] , 
        \g[25][48] , \g[25][47] , \g[25][46] , \g[25][45] , \g[25][44] , 
        \g[25][43] , \g[25][42] , \g[25][41] , \g[25][40] , \g[25][39] , 
        \g[25][38] , \g[25][37] , \g[25][36] , \g[25][35] , \g[25][34] , 
        \g[25][33] , \g[25][32] , \g[25][31] , \g[25][30] , \g[25][29] , 
        \g[25][28] , \g[25][27] , \g[25][26] , \g[25][25] , \g[25][24] , 
        \g[25][23] , \g[25][22] , \g[25][21] , \g[25][20] , \g[25][19] , 
        \g[25][18] , \g[25][17] , \g[25][16] , \g[25][15] , \g[25][14] , 
        \g[25][13] , \g[25][12] , \g[25][11] , \g[25][10] , \g[25][9] , 
        \g[25][8] , \g[25][7] , \g[25][6] , \g[25][5] , \g[25][4] , \g[25][3] , 
        \g[25][2] , \g[25][1] , 1'b0}), .cin({\g[26][63] , \g[26][62] , 
        \g[26][61] , \g[26][60] , \g[26][59] , \g[26][58] , \g[26][57] , 
        \g[26][56] , \g[26][55] , \g[26][54] , \g[26][53] , \g[26][52] , 
        \g[26][51] , \g[26][50] , \g[26][49] , \g[26][48] , \g[26][47] , 
        \g[26][46] , \g[26][45] , \g[26][44] , \g[26][43] , \g[26][42] , 
        \g[26][41] , \g[26][40] , \g[26][39] , \g[26][38] , \g[26][37] , 
        \g[26][36] , \g[26][35] , \g[26][34] , \g[26][33] , \g[26][32] , 
        \g[26][31] , \g[26][30] , \g[26][29] , \g[26][28] , \g[26][27] , 
        \g[26][26] , \g[26][25] , \g[26][24] , \g[26][23] , \g[26][22] , 
        \g[26][21] , \g[26][20] , \g[26][19] , \g[26][18] , \g[26][17] , 
        \g[26][16] , \g[26][15] , \g[26][14] , \g[26][13] , \g[26][12] , 
        \g[26][11] , \g[26][10] , \g[26][9] , \g[26][8] , \g[26][7] , 
        \g[26][6] , \g[26][5] , \g[26][4] , \g[26][3] , \g[26][2] , \g[26][1] , 
        1'b0}), .sum({\g2[8][63] , \g2[8][62] , \g2[8][61] , \g2[8][60] , 
        \g2[8][59] , \g2[8][58] , \g2[8][57] , \g2[8][56] , \g2[8][55] , 
        \g2[8][54] , \g2[8][53] , \g2[8][52] , \g2[8][51] , \g2[8][50] , 
        \g2[8][49] , \g2[8][48] , \g2[8][47] , \g2[8][46] , \g2[8][45] , 
        \g2[8][44] , \g2[8][43] , \g2[8][42] , \g2[8][41] , \g2[8][40] , 
        \g2[8][39] , \g2[8][38] , \g2[8][37] , \g2[8][36] , \g2[8][35] , 
        \g2[8][34] , \g2[8][33] , \g2[8][32] , \g2[8][31] , \g2[8][30] , 
        \g2[8][29] , \g2[8][28] , \g2[8][27] , \g2[8][26] , \g2[8][25] , 
        \g2[8][24] , \g2[8][23] , \g2[8][22] , \g2[8][21] , \g2[8][20] , 
        \g2[8][19] , \g2[8][18] , \g2[8][17] , \g2[8][16] , \g2[8][15] , 
        \g2[8][14] , \g2[8][13] , \g2[8][12] , \g2[8][11] , \g2[8][10] , 
        \g2[8][9] , \g2[8][8] , \g2[8][7] , \g2[8][6] , \g2[8][5] , \g2[8][4] , 
        \g2[8][3] , \g2[8][2] , \g2[8][1] , \g2[8][0] }), .cout({\g2[22][63] , 
        \g2[22][62] , \g2[22][61] , \g2[22][60] , \g2[22][59] , \g2[22][58] , 
        \g2[22][57] , \g2[22][56] , \g2[22][55] , \g2[22][54] , \g2[22][53] , 
        \g2[22][52] , \g2[22][51] , \g2[22][50] , \g2[22][49] , \g2[22][48] , 
        \g2[22][47] , \g2[22][46] , \g2[22][45] , \g2[22][44] , \g2[22][43] , 
        \g2[22][42] , \g2[22][41] , \g2[22][40] , \g2[22][39] , \g2[22][38] , 
        \g2[22][37] , \g2[22][36] , \g2[22][35] , \g2[22][34] , \g2[22][33] , 
        \g2[22][32] , \g2[22][31] , \g2[22][30] , \g2[22][29] , \g2[22][28] , 
        \g2[22][27] , \g2[22][26] , \g2[22][25] , \g2[22][24] , \g2[22][23] , 
        \g2[22][22] , \g2[22][21] , \g2[22][20] , \g2[22][19] , \g2[22][18] , 
        \g2[22][17] , \g2[22][16] , \g2[22][15] , \g2[22][14] , \g2[22][13] , 
        \g2[22][12] , \g2[22][11] , \g2[22][10] , \g2[22][9] , \g2[22][8] , 
        \g2[22][7] , \g2[22][6] , \g2[22][5] , \g2[22][4] , \g2[22][3] , 
        \g2[22][2] , \g2[22][1] , SYNOPSYS_UNCONNECTED__29}) );
  FullAdder_32 \level2[9].x5  ( .a({\g[27][63] , \g[27][62] , \g[27][61] , 
        \g[27][60] , \g[27][59] , \g[27][58] , \g[27][57] , \g[27][56] , 
        \g[27][55] , \g[27][54] , \g[27][53] , \g[27][52] , \g[27][51] , 
        \g[27][50] , \g[27][49] , \g[27][48] , \g[27][47] , \g[27][46] , 
        \g[27][45] , \g[27][44] , \g[27][43] , \g[27][42] , \g[27][41] , 
        \g[27][40] , \g[27][39] , \g[27][38] , \g[27][37] , \g[27][36] , 
        \g[27][35] , \g[27][34] , \g[27][33] , \g[27][32] , \g[27][31] , 
        \g[27][30] , \g[27][29] , \g[27][28] , \g[27][27] , \g[27][26] , 
        \g[27][25] , \g[27][24] , \g[27][23] , \g[27][22] , \g[27][21] , 
        \g[27][20] , \g[27][19] , \g[27][18] , \g[27][17] , \g[27][16] , 
        \g[27][15] , \g[27][14] , \g[27][13] , \g[27][12] , \g[27][11] , 
        \g[27][10] , \g[27][9] , \g[27][8] , \g[27][7] , \g[27][6] , 
        \g[27][5] , \g[27][4] , \g[27][3] , \g[27][2] , \g[27][1] , 1'b0}), 
        .b({\g[28][63] , \g[28][62] , \g[28][61] , \g[28][60] , \g[28][59] , 
        \g[28][58] , \g[28][57] , \g[28][56] , \g[28][55] , \g[28][54] , 
        \g[28][53] , \g[28][52] , \g[28][51] , \g[28][50] , \g[28][49] , 
        \g[28][48] , \g[28][47] , \g[28][46] , \g[28][45] , \g[28][44] , 
        \g[28][43] , \g[28][42] , \g[28][41] , \g[28][40] , \g[28][39] , 
        \g[28][38] , \g[28][37] , \g[28][36] , \g[28][35] , \g[28][34] , 
        \g[28][33] , \g[28][32] , \g[28][31] , \g[28][30] , \g[28][29] , 
        \g[28][28] , \g[28][27] , \g[28][26] , \g[28][25] , \g[28][24] , 
        \g[28][23] , \g[28][22] , \g[28][21] , \g[28][20] , \g[28][19] , 
        \g[28][18] , \g[28][17] , \g[28][16] , \g[28][15] , \g[28][14] , 
        \g[28][13] , \g[28][12] , \g[28][11] , \g[28][10] , \g[28][9] , 
        \g[28][8] , \g[28][7] , \g[28][6] , \g[28][5] , \g[28][4] , \g[28][3] , 
        \g[28][2] , \g[28][1] , 1'b0}), .cin({\g[29][63] , \g[29][62] , 
        \g[29][61] , \g[29][60] , \g[29][59] , \g[29][58] , \g[29][57] , 
        \g[29][56] , \g[29][55] , \g[29][54] , \g[29][53] , \g[29][52] , 
        \g[29][51] , \g[29][50] , \g[29][49] , \g[29][48] , \g[29][47] , 
        \g[29][46] , \g[29][45] , \g[29][44] , \g[29][43] , \g[29][42] , 
        \g[29][41] , \g[29][40] , \g[29][39] , \g[29][38] , \g[29][37] , 
        \g[29][36] , \g[29][35] , \g[29][34] , \g[29][33] , \g[29][32] , 
        \g[29][31] , \g[29][30] , \g[29][29] , \g[29][28] , \g[29][27] , 
        \g[29][26] , \g[29][25] , \g[29][24] , \g[29][23] , \g[29][22] , 
        \g[29][21] , \g[29][20] , \g[29][19] , \g[29][18] , \g[29][17] , 
        \g[29][16] , \g[29][15] , \g[29][14] , \g[29][13] , \g[29][12] , 
        \g[29][11] , \g[29][10] , \g[29][9] , \g[29][8] , \g[29][7] , 
        \g[29][6] , \g[29][5] , \g[29][4] , \g[29][3] , \g[29][2] , \g[29][1] , 
        1'b0}), .sum({\g2[9][63] , \g2[9][62] , \g2[9][61] , \g2[9][60] , 
        \g2[9][59] , \g2[9][58] , \g2[9][57] , \g2[9][56] , \g2[9][55] , 
        \g2[9][54] , \g2[9][53] , \g2[9][52] , \g2[9][51] , \g2[9][50] , 
        \g2[9][49] , \g2[9][48] , \g2[9][47] , \g2[9][46] , \g2[9][45] , 
        \g2[9][44] , \g2[9][43] , \g2[9][42] , \g2[9][41] , \g2[9][40] , 
        \g2[9][39] , \g2[9][38] , \g2[9][37] , \g2[9][36] , \g2[9][35] , 
        \g2[9][34] , \g2[9][33] , \g2[9][32] , \g2[9][31] , \g2[9][30] , 
        \g2[9][29] , \g2[9][28] , \g2[9][27] , \g2[9][26] , \g2[9][25] , 
        \g2[9][24] , \g2[9][23] , \g2[9][22] , \g2[9][21] , \g2[9][20] , 
        \g2[9][19] , \g2[9][18] , \g2[9][17] , \g2[9][16] , \g2[9][15] , 
        \g2[9][14] , \g2[9][13] , \g2[9][12] , \g2[9][11] , \g2[9][10] , 
        \g2[9][9] , \g2[9][8] , \g2[9][7] , \g2[9][6] , \g2[9][5] , \g2[9][4] , 
        \g2[9][3] , \g2[9][2] , \g2[9][1] , \g2[9][0] }), .cout({\g2[23][63] , 
        \g2[23][62] , \g2[23][61] , \g2[23][60] , \g2[23][59] , \g2[23][58] , 
        \g2[23][57] , \g2[23][56] , \g2[23][55] , \g2[23][54] , \g2[23][53] , 
        \g2[23][52] , \g2[23][51] , \g2[23][50] , \g2[23][49] , \g2[23][48] , 
        \g2[23][47] , \g2[23][46] , \g2[23][45] , \g2[23][44] , \g2[23][43] , 
        \g2[23][42] , \g2[23][41] , \g2[23][40] , \g2[23][39] , \g2[23][38] , 
        \g2[23][37] , \g2[23][36] , \g2[23][35] , \g2[23][34] , \g2[23][33] , 
        \g2[23][32] , \g2[23][31] , \g2[23][30] , \g2[23][29] , \g2[23][28] , 
        \g2[23][27] , \g2[23][26] , \g2[23][25] , \g2[23][24] , \g2[23][23] , 
        \g2[23][22] , \g2[23][21] , \g2[23][20] , \g2[23][19] , \g2[23][18] , 
        \g2[23][17] , \g2[23][16] , \g2[23][15] , \g2[23][14] , \g2[23][13] , 
        \g2[23][12] , \g2[23][11] , \g2[23][10] , \g2[23][9] , \g2[23][8] , 
        \g2[23][7] , \g2[23][6] , \g2[23][5] , \g2[23][4] , \g2[23][3] , 
        \g2[23][2] , \g2[23][1] , SYNOPSYS_UNCONNECTED__30}) );
  FullAdder_31 \level2[10].x5  ( .a({\g[30][63] , \g[30][62] , \g[30][61] , 
        \g[30][60] , \g[30][59] , \g[30][58] , \g[30][57] , \g[30][56] , 
        \g[30][55] , \g[30][54] , \g[30][53] , \g[30][52] , \g[30][51] , 
        \g[30][50] , \g[30][49] , \g[30][48] , \g[30][47] , \g[30][46] , 
        \g[30][45] , \g[30][44] , \g[30][43] , \g[30][42] , \g[30][41] , 
        \g[30][40] , \g[30][39] , \g[30][38] , \g[30][37] , \g[30][36] , 
        \g[30][35] , \g[30][34] , \g[30][33] , \g[30][32] , \g[30][31] , 
        \g[30][30] , \g[30][29] , \g[30][28] , \g[30][27] , \g[30][26] , 
        \g[30][25] , \g[30][24] , \g[30][23] , \g[30][22] , \g[30][21] , 
        \g[30][20] , \g[30][19] , \g[30][18] , \g[30][17] , \g[30][16] , 
        \g[30][15] , \g[30][14] , \g[30][13] , \g[30][12] , \g[30][11] , 
        \g[30][10] , \g[30][9] , \g[30][8] , \g[30][7] , \g[30][6] , 
        \g[30][5] , \g[30][4] , \g[30][3] , \g[30][2] , \g[30][1] , 1'b0}), 
        .b({\g[31][63] , \g[31][62] , \g[31][61] , \g[31][60] , \g[31][59] , 
        \g[31][58] , \g[31][57] , \g[31][56] , \g[31][55] , \g[31][54] , 
        \g[31][53] , \g[31][52] , \g[31][51] , \g[31][50] , \g[31][49] , 
        \g[31][48] , \g[31][47] , \g[31][46] , \g[31][45] , \g[31][44] , 
        \g[31][43] , \g[31][42] , \g[31][41] , \g[31][40] , \g[31][39] , 
        \g[31][38] , \g[31][37] , \g[31][36] , \g[31][35] , \g[31][34] , 
        \g[31][33] , \g[31][32] , \g[31][31] , \g[31][30] , \g[31][29] , 
        \g[31][28] , \g[31][27] , \g[31][26] , \g[31][25] , \g[31][24] , 
        \g[31][23] , \g[31][22] , \g[31][21] , \g[31][20] , \g[31][19] , 
        \g[31][18] , \g[31][17] , \g[31][16] , \g[31][15] , \g[31][14] , 
        \g[31][13] , \g[31][12] , \g[31][11] , \g[31][10] , \g[31][9] , 
        \g[31][8] , \g[31][7] , \g[31][6] , \g[31][5] , \g[31][4] , \g[31][3] , 
        \g[31][2] , \g[31][1] , 1'b0}), .cin({\g[32][63] , \g[32][62] , 
        \g[32][61] , \g[32][60] , \g[32][59] , \g[32][58] , \g[32][57] , 
        \g[32][56] , \g[32][55] , \g[32][54] , \g[32][53] , \g[32][52] , 
        \g[32][51] , \g[32][50] , \g[32][49] , \g[32][48] , \g[32][47] , 
        \g[32][46] , \g[32][45] , \g[32][44] , \g[32][43] , \g[32][42] , 
        \g[32][41] , \g[32][40] , \g[32][39] , \g[32][38] , \g[32][37] , 
        \g[32][36] , \g[32][35] , \g[32][34] , \g[32][33] , \g[32][32] , 
        \g[32][31] , \g[32][30] , \g[32][29] , \g[32][28] , \g[32][27] , 
        \g[32][26] , \g[32][25] , \g[32][24] , \g[32][23] , \g[32][22] , 
        \g[32][21] , \g[32][20] , \g[32][19] , \g[32][18] , \g[32][17] , 
        \g[32][16] , \g[32][15] , \g[32][14] , \g[32][13] , \g[32][12] , 
        \g[32][11] , \g[32][10] , \g[32][9] , \g[32][8] , \g[32][7] , 
        \g[32][6] , \g[32][5] , \g[32][4] , \g[32][3] , \g[32][2] , \g[32][1] , 
        1'b0}), .sum({\g2[10][63] , \g2[10][62] , \g2[10][61] , \g2[10][60] , 
        \g2[10][59] , \g2[10][58] , \g2[10][57] , \g2[10][56] , \g2[10][55] , 
        \g2[10][54] , \g2[10][53] , \g2[10][52] , \g2[10][51] , \g2[10][50] , 
        \g2[10][49] , \g2[10][48] , \g2[10][47] , \g2[10][46] , \g2[10][45] , 
        \g2[10][44] , \g2[10][43] , \g2[10][42] , \g2[10][41] , \g2[10][40] , 
        \g2[10][39] , \g2[10][38] , \g2[10][37] , \g2[10][36] , \g2[10][35] , 
        \g2[10][34] , \g2[10][33] , \g2[10][32] , \g2[10][31] , \g2[10][30] , 
        \g2[10][29] , \g2[10][28] , \g2[10][27] , \g2[10][26] , \g2[10][25] , 
        \g2[10][24] , \g2[10][23] , \g2[10][22] , \g2[10][21] , \g2[10][20] , 
        \g2[10][19] , \g2[10][18] , \g2[10][17] , \g2[10][16] , \g2[10][15] , 
        \g2[10][14] , \g2[10][13] , \g2[10][12] , \g2[10][11] , \g2[10][10] , 
        \g2[10][9] , \g2[10][8] , \g2[10][7] , \g2[10][6] , \g2[10][5] , 
        \g2[10][4] , \g2[10][3] , \g2[10][2] , \g2[10][1] , \g2[10][0] }), 
        .cout({\g2[24][63] , \g2[24][62] , \g2[24][61] , \g2[24][60] , 
        \g2[24][59] , \g2[24][58] , \g2[24][57] , \g2[24][56] , \g2[24][55] , 
        \g2[24][54] , \g2[24][53] , \g2[24][52] , \g2[24][51] , \g2[24][50] , 
        \g2[24][49] , \g2[24][48] , \g2[24][47] , \g2[24][46] , \g2[24][45] , 
        \g2[24][44] , \g2[24][43] , \g2[24][42] , \g2[24][41] , \g2[24][40] , 
        \g2[24][39] , \g2[24][38] , \g2[24][37] , \g2[24][36] , \g2[24][35] , 
        \g2[24][34] , \g2[24][33] , \g2[24][32] , \g2[24][31] , \g2[24][30] , 
        \g2[24][29] , \g2[24][28] , \g2[24][27] , \g2[24][26] , \g2[24][25] , 
        \g2[24][24] , \g2[24][23] , \g2[24][22] , \g2[24][21] , \g2[24][20] , 
        \g2[24][19] , \g2[24][18] , \g2[24][17] , \g2[24][16] , \g2[24][15] , 
        \g2[24][14] , \g2[24][13] , \g2[24][12] , \g2[24][11] , \g2[24][10] , 
        \g2[24][9] , \g2[24][8] , \g2[24][7] , \g2[24][6] , \g2[24][5] , 
        \g2[24][4] , \g2[24][3] , \g2[24][2] , \g2[24][1] , 
        SYNOPSYS_UNCONNECTED__31}) );
  FullAdder_30 \level2[11].x5  ( .a({\g[33][63] , \g[33][62] , \g[33][61] , 
        \g[33][60] , \g[33][59] , \g[33][58] , \g[33][57] , \g[33][56] , 
        \g[33][55] , \g[33][54] , \g[33][53] , \g[33][52] , \g[33][51] , 
        \g[33][50] , \g[33][49] , \g[33][48] , \g[33][47] , \g[33][46] , 
        \g[33][45] , \g[33][44] , \g[33][43] , \g[33][42] , \g[33][41] , 
        \g[33][40] , \g[33][39] , \g[33][38] , \g[33][37] , \g[33][36] , 
        \g[33][35] , \g[33][34] , \g[33][33] , \g[33][32] , \g[33][31] , 
        \g[33][30] , \g[33][29] , \g[33][28] , \g[33][27] , \g[33][26] , 
        \g[33][25] , \g[33][24] , \g[33][23] , \g[33][22] , \g[33][21] , 
        \g[33][20] , \g[33][19] , \g[33][18] , \g[33][17] , \g[33][16] , 
        \g[33][15] , \g[33][14] , \g[33][13] , \g[33][12] , \g[33][11] , 
        \g[33][10] , \g[33][9] , \g[33][8] , \g[33][7] , \g[33][6] , 
        \g[33][5] , \g[33][4] , \g[33][3] , \g[33][2] , \g[33][1] , 1'b0}), 
        .b({\g[34][63] , \g[34][62] , \g[34][61] , \g[34][60] , \g[34][59] , 
        \g[34][58] , \g[34][57] , \g[34][56] , \g[34][55] , \g[34][54] , 
        \g[34][53] , \g[34][52] , \g[34][51] , \g[34][50] , \g[34][49] , 
        \g[34][48] , \g[34][47] , \g[34][46] , \g[34][45] , \g[34][44] , 
        \g[34][43] , \g[34][42] , \g[34][41] , \g[34][40] , \g[34][39] , 
        \g[34][38] , \g[34][37] , \g[34][36] , \g[34][35] , \g[34][34] , 
        \g[34][33] , \g[34][32] , \g[34][31] , \g[34][30] , \g[34][29] , 
        \g[34][28] , \g[34][27] , \g[34][26] , \g[34][25] , \g[34][24] , 
        \g[34][23] , \g[34][22] , \g[34][21] , \g[34][20] , \g[34][19] , 
        \g[34][18] , \g[34][17] , \g[34][16] , \g[34][15] , \g[34][14] , 
        \g[34][13] , \g[34][12] , \g[34][11] , \g[34][10] , \g[34][9] , 
        \g[34][8] , \g[34][7] , \g[34][6] , \g[34][5] , \g[34][4] , \g[34][3] , 
        \g[34][2] , \g[34][1] , 1'b0}), .cin({\g[35][63] , \g[35][62] , 
        \g[35][61] , \g[35][60] , \g[35][59] , \g[35][58] , \g[35][57] , 
        \g[35][56] , \g[35][55] , \g[35][54] , \g[35][53] , \g[35][52] , 
        \g[35][51] , \g[35][50] , \g[35][49] , \g[35][48] , \g[35][47] , 
        \g[35][46] , \g[35][45] , \g[35][44] , \g[35][43] , \g[35][42] , 
        \g[35][41] , \g[35][40] , \g[35][39] , \g[35][38] , \g[35][37] , 
        \g[35][36] , \g[35][35] , \g[35][34] , \g[35][33] , \g[35][32] , 
        \g[35][31] , \g[35][30] , \g[35][29] , \g[35][28] , \g[35][27] , 
        \g[35][26] , \g[35][25] , \g[35][24] , \g[35][23] , \g[35][22] , 
        \g[35][21] , \g[35][20] , \g[35][19] , \g[35][18] , \g[35][17] , 
        \g[35][16] , \g[35][15] , \g[35][14] , \g[35][13] , \g[35][12] , 
        \g[35][11] , \g[35][10] , \g[35][9] , \g[35][8] , \g[35][7] , 
        \g[35][6] , \g[35][5] , \g[35][4] , \g[35][3] , \g[35][2] , \g[35][1] , 
        1'b0}), .sum({\g2[11][63] , \g2[11][62] , \g2[11][61] , \g2[11][60] , 
        \g2[11][59] , \g2[11][58] , \g2[11][57] , \g2[11][56] , \g2[11][55] , 
        \g2[11][54] , \g2[11][53] , \g2[11][52] , \g2[11][51] , \g2[11][50] , 
        \g2[11][49] , \g2[11][48] , \g2[11][47] , \g2[11][46] , \g2[11][45] , 
        \g2[11][44] , \g2[11][43] , \g2[11][42] , \g2[11][41] , \g2[11][40] , 
        \g2[11][39] , \g2[11][38] , \g2[11][37] , \g2[11][36] , \g2[11][35] , 
        \g2[11][34] , \g2[11][33] , \g2[11][32] , \g2[11][31] , \g2[11][30] , 
        \g2[11][29] , \g2[11][28] , \g2[11][27] , \g2[11][26] , \g2[11][25] , 
        \g2[11][24] , \g2[11][23] , \g2[11][22] , \g2[11][21] , \g2[11][20] , 
        \g2[11][19] , \g2[11][18] , \g2[11][17] , \g2[11][16] , \g2[11][15] , 
        \g2[11][14] , \g2[11][13] , \g2[11][12] , \g2[11][11] , \g2[11][10] , 
        \g2[11][9] , \g2[11][8] , \g2[11][7] , \g2[11][6] , \g2[11][5] , 
        \g2[11][4] , \g2[11][3] , \g2[11][2] , \g2[11][1] , \g2[11][0] }), 
        .cout({\g2[25][63] , \g2[25][62] , \g2[25][61] , \g2[25][60] , 
        \g2[25][59] , \g2[25][58] , \g2[25][57] , \g2[25][56] , \g2[25][55] , 
        \g2[25][54] , \g2[25][53] , \g2[25][52] , \g2[25][51] , \g2[25][50] , 
        \g2[25][49] , \g2[25][48] , \g2[25][47] , \g2[25][46] , \g2[25][45] , 
        \g2[25][44] , \g2[25][43] , \g2[25][42] , \g2[25][41] , \g2[25][40] , 
        \g2[25][39] , \g2[25][38] , \g2[25][37] , \g2[25][36] , \g2[25][35] , 
        \g2[25][34] , \g2[25][33] , \g2[25][32] , \g2[25][31] , \g2[25][30] , 
        \g2[25][29] , \g2[25][28] , \g2[25][27] , \g2[25][26] , \g2[25][25] , 
        \g2[25][24] , \g2[25][23] , \g2[25][22] , \g2[25][21] , \g2[25][20] , 
        \g2[25][19] , \g2[25][18] , \g2[25][17] , \g2[25][16] , \g2[25][15] , 
        \g2[25][14] , \g2[25][13] , \g2[25][12] , \g2[25][11] , \g2[25][10] , 
        \g2[25][9] , \g2[25][8] , \g2[25][7] , \g2[25][6] , \g2[25][5] , 
        \g2[25][4] , \g2[25][3] , \g2[25][2] , \g2[25][1] , 
        SYNOPSYS_UNCONNECTED__32}) );
  FullAdder_29 \level2[12].x5  ( .a({\g[36][63] , \g[36][62] , \g[36][61] , 
        \g[36][60] , \g[36][59] , \g[36][58] , \g[36][57] , \g[36][56] , 
        \g[36][55] , \g[36][54] , \g[36][53] , \g[36][52] , \g[36][51] , 
        \g[36][50] , \g[36][49] , \g[36][48] , \g[36][47] , \g[36][46] , 
        \g[36][45] , \g[36][44] , \g[36][43] , \g[36][42] , \g[36][41] , 
        \g[36][40] , \g[36][39] , \g[36][38] , \g[36][37] , \g[36][36] , 
        \g[36][35] , \g[36][34] , \g[36][33] , \g[36][32] , \g[36][31] , 
        \g[36][30] , \g[36][29] , \g[36][28] , \g[36][27] , \g[36][26] , 
        \g[36][25] , \g[36][24] , \g[36][23] , \g[36][22] , \g[36][21] , 
        \g[36][20] , \g[36][19] , \g[36][18] , \g[36][17] , \g[36][16] , 
        \g[36][15] , \g[36][14] , \g[36][13] , \g[36][12] , \g[36][11] , 
        \g[36][10] , \g[36][9] , \g[36][8] , \g[36][7] , \g[36][6] , 
        \g[36][5] , \g[36][4] , \g[36][3] , \g[36][2] , \g[36][1] , 1'b0}), 
        .b({\g[37][63] , \g[37][62] , \g[37][61] , \g[37][60] , \g[37][59] , 
        \g[37][58] , \g[37][57] , \g[37][56] , \g[37][55] , \g[37][54] , 
        \g[37][53] , \g[37][52] , \g[37][51] , \g[37][50] , \g[37][49] , 
        \g[37][48] , \g[37][47] , \g[37][46] , \g[37][45] , \g[37][44] , 
        \g[37][43] , \g[37][42] , \g[37][41] , \g[37][40] , \g[37][39] , 
        \g[37][38] , \g[37][37] , \g[37][36] , \g[37][35] , \g[37][34] , 
        \g[37][33] , \g[37][32] , \g[37][31] , \g[37][30] , \g[37][29] , 
        \g[37][28] , \g[37][27] , \g[37][26] , \g[37][25] , \g[37][24] , 
        \g[37][23] , \g[37][22] , \g[37][21] , \g[37][20] , \g[37][19] , 
        \g[37][18] , \g[37][17] , \g[37][16] , \g[37][15] , \g[37][14] , 
        \g[37][13] , \g[37][12] , \g[37][11] , \g[37][10] , \g[37][9] , 
        \g[37][8] , \g[37][7] , \g[37][6] , \g[37][5] , \g[37][4] , \g[37][3] , 
        \g[37][2] , \g[37][1] , 1'b0}), .cin({\g[38][63] , \g[38][62] , 
        \g[38][61] , \g[38][60] , \g[38][59] , \g[38][58] , \g[38][57] , 
        \g[38][56] , \g[38][55] , \g[38][54] , \g[38][53] , \g[38][52] , 
        \g[38][51] , \g[38][50] , \g[38][49] , \g[38][48] , \g[38][47] , 
        \g[38][46] , \g[38][45] , \g[38][44] , \g[38][43] , \g[38][42] , 
        \g[38][41] , \g[38][40] , \g[38][39] , \g[38][38] , \g[38][37] , 
        \g[38][36] , \g[38][35] , \g[38][34] , \g[38][33] , \g[38][32] , 
        \g[38][31] , \g[38][30] , \g[38][29] , \g[38][28] , \g[38][27] , 
        \g[38][26] , \g[38][25] , \g[38][24] , \g[38][23] , \g[38][22] , 
        \g[38][21] , \g[38][20] , \g[38][19] , \g[38][18] , \g[38][17] , 
        \g[38][16] , \g[38][15] , \g[38][14] , \g[38][13] , \g[38][12] , 
        \g[38][11] , \g[38][10] , \g[38][9] , \g[38][8] , \g[38][7] , 
        \g[38][6] , \g[38][5] , \g[38][4] , \g[38][3] , \g[38][2] , \g[38][1] , 
        1'b0}), .sum({\g2[12][63] , \g2[12][62] , \g2[12][61] , \g2[12][60] , 
        \g2[12][59] , \g2[12][58] , \g2[12][57] , \g2[12][56] , \g2[12][55] , 
        \g2[12][54] , \g2[12][53] , \g2[12][52] , \g2[12][51] , \g2[12][50] , 
        \g2[12][49] , \g2[12][48] , \g2[12][47] , \g2[12][46] , \g2[12][45] , 
        \g2[12][44] , \g2[12][43] , \g2[12][42] , \g2[12][41] , \g2[12][40] , 
        \g2[12][39] , \g2[12][38] , \g2[12][37] , \g2[12][36] , \g2[12][35] , 
        \g2[12][34] , \g2[12][33] , \g2[12][32] , \g2[12][31] , \g2[12][30] , 
        \g2[12][29] , \g2[12][28] , \g2[12][27] , \g2[12][26] , \g2[12][25] , 
        \g2[12][24] , \g2[12][23] , \g2[12][22] , \g2[12][21] , \g2[12][20] , 
        \g2[12][19] , \g2[12][18] , \g2[12][17] , \g2[12][16] , \g2[12][15] , 
        \g2[12][14] , \g2[12][13] , \g2[12][12] , \g2[12][11] , \g2[12][10] , 
        \g2[12][9] , \g2[12][8] , \g2[12][7] , \g2[12][6] , \g2[12][5] , 
        \g2[12][4] , \g2[12][3] , \g2[12][2] , \g2[12][1] , \g2[12][0] }), 
        .cout({\g2[26][63] , \g2[26][62] , \g2[26][61] , \g2[26][60] , 
        \g2[26][59] , \g2[26][58] , \g2[26][57] , \g2[26][56] , \g2[26][55] , 
        \g2[26][54] , \g2[26][53] , \g2[26][52] , \g2[26][51] , \g2[26][50] , 
        \g2[26][49] , \g2[26][48] , \g2[26][47] , \g2[26][46] , \g2[26][45] , 
        \g2[26][44] , \g2[26][43] , \g2[26][42] , \g2[26][41] , \g2[26][40] , 
        \g2[26][39] , \g2[26][38] , \g2[26][37] , \g2[26][36] , \g2[26][35] , 
        \g2[26][34] , \g2[26][33] , \g2[26][32] , \g2[26][31] , \g2[26][30] , 
        \g2[26][29] , \g2[26][28] , \g2[26][27] , \g2[26][26] , \g2[26][25] , 
        \g2[26][24] , \g2[26][23] , \g2[26][22] , \g2[26][21] , \g2[26][20] , 
        \g2[26][19] , \g2[26][18] , \g2[26][17] , \g2[26][16] , \g2[26][15] , 
        \g2[26][14] , \g2[26][13] , \g2[26][12] , \g2[26][11] , \g2[26][10] , 
        \g2[26][9] , \g2[26][8] , \g2[26][7] , \g2[26][6] , \g2[26][5] , 
        \g2[26][4] , \g2[26][3] , \g2[26][2] , \g2[26][1] , 
        SYNOPSYS_UNCONNECTED__33}) );
  FullAdder_28 \level2[13].x5  ( .a({\g[39][63] , \g[39][62] , \g[39][61] , 
        \g[39][60] , \g[39][59] , \g[39][58] , \g[39][57] , \g[39][56] , 
        \g[39][55] , \g[39][54] , \g[39][53] , \g[39][52] , \g[39][51] , 
        \g[39][50] , \g[39][49] , \g[39][48] , \g[39][47] , \g[39][46] , 
        \g[39][45] , \g[39][44] , \g[39][43] , \g[39][42] , \g[39][41] , 
        \g[39][40] , \g[39][39] , \g[39][38] , \g[39][37] , \g[39][36] , 
        \g[39][35] , \g[39][34] , \g[39][33] , \g[39][32] , \g[39][31] , 
        \g[39][30] , \g[39][29] , \g[39][28] , \g[39][27] , \g[39][26] , 
        \g[39][25] , \g[39][24] , \g[39][23] , \g[39][22] , \g[39][21] , 
        \g[39][20] , \g[39][19] , \g[39][18] , \g[39][17] , \g[39][16] , 
        \g[39][15] , \g[39][14] , \g[39][13] , \g[39][12] , \g[39][11] , 
        \g[39][10] , \g[39][9] , \g[39][8] , \g[39][7] , \g[39][6] , 
        \g[39][5] , \g[39][4] , \g[39][3] , \g[39][2] , \g[39][1] , 1'b0}), 
        .b({\g[40][63] , \g[40][62] , \g[40][61] , \g[40][60] , \g[40][59] , 
        \g[40][58] , \g[40][57] , \g[40][56] , \g[40][55] , \g[40][54] , 
        \g[40][53] , \g[40][52] , \g[40][51] , \g[40][50] , \g[40][49] , 
        \g[40][48] , \g[40][47] , \g[40][46] , \g[40][45] , \g[40][44] , 
        \g[40][43] , \g[40][42] , \g[40][41] , \g[40][40] , \g[40][39] , 
        \g[40][38] , \g[40][37] , \g[40][36] , \g[40][35] , \g[40][34] , 
        \g[40][33] , \g[40][32] , \g[40][31] , \g[40][30] , \g[40][29] , 
        \g[40][28] , \g[40][27] , \g[40][26] , \g[40][25] , \g[40][24] , 
        \g[40][23] , \g[40][22] , \g[40][21] , \g[40][20] , \g[40][19] , 
        \g[40][18] , \g[40][17] , \g[40][16] , \g[40][15] , \g[40][14] , 
        \g[40][13] , \g[40][12] , \g[40][11] , \g[40][10] , \g[40][9] , 
        \g[40][8] , \g[40][7] , \g[40][6] , \g[40][5] , \g[40][4] , \g[40][3] , 
        \g[40][2] , \g[40][1] , 1'b0}), .cin({\g[41][63] , \g[41][62] , 
        \g[41][61] , \g[41][60] , \g[41][59] , \g[41][58] , \g[41][57] , 
        \g[41][56] , \g[41][55] , \g[41][54] , \g[41][53] , \g[41][52] , 
        \g[41][51] , \g[41][50] , \g[41][49] , \g[41][48] , \g[41][47] , 
        \g[41][46] , \g[41][45] , \g[41][44] , \g[41][43] , \g[41][42] , 
        \g[41][41] , \g[41][40] , \g[41][39] , \g[41][38] , \g[41][37] , 
        \g[41][36] , \g[41][35] , \g[41][34] , \g[41][33] , \g[41][32] , 
        \g[41][31] , \g[41][30] , \g[41][29] , \g[41][28] , \g[41][27] , 
        \g[41][26] , \g[41][25] , \g[41][24] , \g[41][23] , \g[41][22] , 
        \g[41][21] , \g[41][20] , \g[41][19] , \g[41][18] , \g[41][17] , 
        \g[41][16] , \g[41][15] , \g[41][14] , \g[41][13] , \g[41][12] , 
        \g[41][11] , \g[41][10] , \g[41][9] , \g[41][8] , \g[41][7] , 
        \g[41][6] , \g[41][5] , \g[41][4] , \g[41][3] , \g[41][2] , \g[41][1] , 
        1'b0}), .sum({\g2[13][63] , \g2[13][62] , \g2[13][61] , \g2[13][60] , 
        \g2[13][59] , \g2[13][58] , \g2[13][57] , \g2[13][56] , \g2[13][55] , 
        \g2[13][54] , \g2[13][53] , \g2[13][52] , \g2[13][51] , \g2[13][50] , 
        \g2[13][49] , \g2[13][48] , \g2[13][47] , \g2[13][46] , \g2[13][45] , 
        \g2[13][44] , \g2[13][43] , \g2[13][42] , \g2[13][41] , \g2[13][40] , 
        \g2[13][39] , \g2[13][38] , \g2[13][37] , \g2[13][36] , \g2[13][35] , 
        \g2[13][34] , \g2[13][33] , \g2[13][32] , \g2[13][31] , \g2[13][30] , 
        \g2[13][29] , \g2[13][28] , \g2[13][27] , \g2[13][26] , \g2[13][25] , 
        \g2[13][24] , \g2[13][23] , \g2[13][22] , \g2[13][21] , \g2[13][20] , 
        \g2[13][19] , \g2[13][18] , \g2[13][17] , \g2[13][16] , \g2[13][15] , 
        \g2[13][14] , \g2[13][13] , \g2[13][12] , \g2[13][11] , \g2[13][10] , 
        \g2[13][9] , \g2[13][8] , \g2[13][7] , \g2[13][6] , \g2[13][5] , 
        \g2[13][4] , \g2[13][3] , \g2[13][2] , \g2[13][1] , \g2[13][0] }), 
        .cout({\g2[27][63] , \g2[27][62] , \g2[27][61] , \g2[27][60] , 
        \g2[27][59] , \g2[27][58] , \g2[27][57] , \g2[27][56] , \g2[27][55] , 
        \g2[27][54] , \g2[27][53] , \g2[27][52] , \g2[27][51] , \g2[27][50] , 
        \g2[27][49] , \g2[27][48] , \g2[27][47] , \g2[27][46] , \g2[27][45] , 
        \g2[27][44] , \g2[27][43] , \g2[27][42] , \g2[27][41] , \g2[27][40] , 
        \g2[27][39] , \g2[27][38] , \g2[27][37] , \g2[27][36] , \g2[27][35] , 
        \g2[27][34] , \g2[27][33] , \g2[27][32] , \g2[27][31] , \g2[27][30] , 
        \g2[27][29] , \g2[27][28] , \g2[27][27] , \g2[27][26] , \g2[27][25] , 
        \g2[27][24] , \g2[27][23] , \g2[27][22] , \g2[27][21] , \g2[27][20] , 
        \g2[27][19] , \g2[27][18] , \g2[27][17] , \g2[27][16] , \g2[27][15] , 
        \g2[27][14] , \g2[27][13] , \g2[27][12] , \g2[27][11] , \g2[27][10] , 
        \g2[27][9] , \g2[27][8] , \g2[27][7] , \g2[27][6] , \g2[27][5] , 
        \g2[27][4] , \g2[27][3] , \g2[27][2] , \g2[27][1] , 
        SYNOPSYS_UNCONNECTED__34}) );
  FullAdder_27 \level3[0].x0  ( .a({\g2[0][63] , \g2[0][62] , \g2[0][61] , 
        \g2[0][60] , \g2[0][59] , \g2[0][58] , \g2[0][57] , \g2[0][56] , 
        \g2[0][55] , \g2[0][54] , \g2[0][53] , \g2[0][52] , \g2[0][51] , 
        \g2[0][50] , \g2[0][49] , \g2[0][48] , \g2[0][47] , \g2[0][46] , 
        \g2[0][45] , \g2[0][44] , \g2[0][43] , \g2[0][42] , \g2[0][41] , 
        \g2[0][40] , \g2[0][39] , \g2[0][38] , \g2[0][37] , \g2[0][36] , 
        \g2[0][35] , \g2[0][34] , \g2[0][33] , \g2[0][32] , \g2[0][31] , 
        \g2[0][30] , \g2[0][29] , \g2[0][28] , \g2[0][27] , \g2[0][26] , 
        \g2[0][25] , \g2[0][24] , \g2[0][23] , \g2[0][22] , \g2[0][21] , 
        \g2[0][20] , \g2[0][19] , \g2[0][18] , \g2[0][17] , \g2[0][16] , 
        \g2[0][15] , \g2[0][14] , \g2[0][13] , \g2[0][12] , \g2[0][11] , 
        \g2[0][10] , \g2[0][9] , \g2[0][8] , \g2[0][7] , \g2[0][6] , 
        \g2[0][5] , \g2[0][4] , \g2[0][3] , \g2[0][2] , \g2[0][1] , \g2[0][0] }), .b({\g2[1][63] , \g2[1][62] , \g2[1][61] , \g2[1][60] , \g2[1][59] , 
        \g2[1][58] , \g2[1][57] , \g2[1][56] , \g2[1][55] , \g2[1][54] , 
        \g2[1][53] , \g2[1][52] , \g2[1][51] , \g2[1][50] , \g2[1][49] , 
        \g2[1][48] , \g2[1][47] , \g2[1][46] , \g2[1][45] , \g2[1][44] , 
        \g2[1][43] , \g2[1][42] , \g2[1][41] , \g2[1][40] , \g2[1][39] , 
        \g2[1][38] , \g2[1][37] , \g2[1][36] , \g2[1][35] , \g2[1][34] , 
        \g2[1][33] , \g2[1][32] , \g2[1][31] , \g2[1][30] , \g2[1][29] , 
        \g2[1][28] , \g2[1][27] , \g2[1][26] , \g2[1][25] , \g2[1][24] , 
        \g2[1][23] , \g2[1][22] , \g2[1][21] , \g2[1][20] , \g2[1][19] , 
        \g2[1][18] , \g2[1][17] , \g2[1][16] , \g2[1][15] , \g2[1][14] , 
        \g2[1][13] , \g2[1][12] , \g2[1][11] , \g2[1][10] , \g2[1][9] , 
        \g2[1][8] , \g2[1][7] , \g2[1][6] , \g2[1][5] , \g2[1][4] , \g2[1][3] , 
        \g2[1][2] , \g2[1][1] , \g2[1][0] }), .cin({\g2[2][63] , \g2[2][62] , 
        \g2[2][61] , \g2[2][60] , \g2[2][59] , \g2[2][58] , \g2[2][57] , 
        \g2[2][56] , \g2[2][55] , \g2[2][54] , \g2[2][53] , \g2[2][52] , 
        \g2[2][51] , \g2[2][50] , \g2[2][49] , \g2[2][48] , \g2[2][47] , 
        \g2[2][46] , \g2[2][45] , \g2[2][44] , \g2[2][43] , \g2[2][42] , 
        \g2[2][41] , \g2[2][40] , \g2[2][39] , \g2[2][38] , \g2[2][37] , 
        \g2[2][36] , \g2[2][35] , \g2[2][34] , \g2[2][33] , \g2[2][32] , 
        \g2[2][31] , \g2[2][30] , \g2[2][29] , \g2[2][28] , \g2[2][27] , 
        \g2[2][26] , \g2[2][25] , \g2[2][24] , \g2[2][23] , \g2[2][22] , 
        \g2[2][21] , \g2[2][20] , \g2[2][19] , \g2[2][18] , \g2[2][17] , 
        \g2[2][16] , \g2[2][15] , \g2[2][14] , \g2[2][13] , \g2[2][12] , 
        \g2[2][11] , \g2[2][10] , \g2[2][9] , \g2[2][8] , \g2[2][7] , 
        \g2[2][6] , \g2[2][5] , \g2[2][4] , \g2[2][3] , \g2[2][2] , \g2[2][1] , 
        \g2[2][0] }), .sum({\g3[0][63] , \g3[0][62] , \g3[0][61] , \g3[0][60] , 
        \g3[0][59] , \g3[0][58] , \g3[0][57] , \g3[0][56] , \g3[0][55] , 
        \g3[0][54] , \g3[0][53] , \g3[0][52] , \g3[0][51] , \g3[0][50] , 
        \g3[0][49] , \g3[0][48] , \g3[0][47] , \g3[0][46] , \g3[0][45] , 
        \g3[0][44] , \g3[0][43] , \g3[0][42] , \g3[0][41] , \g3[0][40] , 
        \g3[0][39] , \g3[0][38] , \g3[0][37] , \g3[0][36] , \g3[0][35] , 
        \g3[0][34] , \g3[0][33] , \g3[0][32] , \g3[0][31] , \g3[0][30] , 
        \g3[0][29] , \g3[0][28] , \g3[0][27] , \g3[0][26] , \g3[0][25] , 
        \g3[0][24] , \g3[0][23] , \g3[0][22] , \g3[0][21] , \g3[0][20] , 
        \g3[0][19] , \g3[0][18] , \g3[0][17] , \g3[0][16] , \g3[0][15] , 
        \g3[0][14] , \g3[0][13] , \g3[0][12] , \g3[0][11] , \g3[0][10] , 
        \g3[0][9] , \g3[0][8] , \g3[0][7] , \g3[0][6] , \g3[0][5] , \g3[0][4] , 
        \g3[0][3] , \g3[0][2] , \g3[0][1] , \g3[0][0] }), .cout({\g3[9][63] , 
        \g3[9][62] , \g3[9][61] , \g3[9][60] , \g3[9][59] , \g3[9][58] , 
        \g3[9][57] , \g3[9][56] , \g3[9][55] , \g3[9][54] , \g3[9][53] , 
        \g3[9][52] , \g3[9][51] , \g3[9][50] , \g3[9][49] , \g3[9][48] , 
        \g3[9][47] , \g3[9][46] , \g3[9][45] , \g3[9][44] , \g3[9][43] , 
        \g3[9][42] , \g3[9][41] , \g3[9][40] , \g3[9][39] , \g3[9][38] , 
        \g3[9][37] , \g3[9][36] , \g3[9][35] , \g3[9][34] , \g3[9][33] , 
        \g3[9][32] , \g3[9][31] , \g3[9][30] , \g3[9][29] , \g3[9][28] , 
        \g3[9][27] , \g3[9][26] , \g3[9][25] , \g3[9][24] , \g3[9][23] , 
        \g3[9][22] , \g3[9][21] , \g3[9][20] , \g3[9][19] , \g3[9][18] , 
        \g3[9][17] , \g3[9][16] , \g3[9][15] , \g3[9][14] , \g3[9][13] , 
        \g3[9][12] , \g3[9][11] , \g3[9][10] , \g3[9][9] , \g3[9][8] , 
        \g3[9][7] , \g3[9][6] , \g3[9][5] , \g3[9][4] , \g3[9][3] , \g3[9][2] , 
        \g3[9][1] , SYNOPSYS_UNCONNECTED__35}) );
  FullAdder_26 \level3[1].x0  ( .a({\g2[3][63] , \g2[3][62] , \g2[3][61] , 
        \g2[3][60] , \g2[3][59] , \g2[3][58] , \g2[3][57] , \g2[3][56] , 
        \g2[3][55] , \g2[3][54] , \g2[3][53] , \g2[3][52] , \g2[3][51] , 
        \g2[3][50] , \g2[3][49] , \g2[3][48] , \g2[3][47] , \g2[3][46] , 
        \g2[3][45] , \g2[3][44] , \g2[3][43] , \g2[3][42] , \g2[3][41] , 
        \g2[3][40] , \g2[3][39] , \g2[3][38] , \g2[3][37] , \g2[3][36] , 
        \g2[3][35] , \g2[3][34] , \g2[3][33] , \g2[3][32] , \g2[3][31] , 
        \g2[3][30] , \g2[3][29] , \g2[3][28] , \g2[3][27] , \g2[3][26] , 
        \g2[3][25] , \g2[3][24] , \g2[3][23] , \g2[3][22] , \g2[3][21] , 
        \g2[3][20] , \g2[3][19] , \g2[3][18] , \g2[3][17] , \g2[3][16] , 
        \g2[3][15] , \g2[3][14] , \g2[3][13] , \g2[3][12] , \g2[3][11] , 
        \g2[3][10] , \g2[3][9] , \g2[3][8] , \g2[3][7] , \g2[3][6] , 
        \g2[3][5] , \g2[3][4] , \g2[3][3] , \g2[3][2] , \g2[3][1] , \g2[3][0] }), .b({\g2[4][63] , \g2[4][62] , \g2[4][61] , \g2[4][60] , \g2[4][59] , 
        \g2[4][58] , \g2[4][57] , \g2[4][56] , \g2[4][55] , \g2[4][54] , 
        \g2[4][53] , \g2[4][52] , \g2[4][51] , \g2[4][50] , \g2[4][49] , 
        \g2[4][48] , \g2[4][47] , \g2[4][46] , \g2[4][45] , \g2[4][44] , 
        \g2[4][43] , \g2[4][42] , \g2[4][41] , \g2[4][40] , \g2[4][39] , 
        \g2[4][38] , \g2[4][37] , \g2[4][36] , \g2[4][35] , \g2[4][34] , 
        \g2[4][33] , \g2[4][32] , \g2[4][31] , \g2[4][30] , \g2[4][29] , 
        \g2[4][28] , \g2[4][27] , \g2[4][26] , \g2[4][25] , \g2[4][24] , 
        \g2[4][23] , \g2[4][22] , \g2[4][21] , \g2[4][20] , \g2[4][19] , 
        \g2[4][18] , \g2[4][17] , \g2[4][16] , \g2[4][15] , \g2[4][14] , 
        \g2[4][13] , \g2[4][12] , \g2[4][11] , \g2[4][10] , \g2[4][9] , 
        \g2[4][8] , \g2[4][7] , \g2[4][6] , \g2[4][5] , \g2[4][4] , \g2[4][3] , 
        \g2[4][2] , \g2[4][1] , \g2[4][0] }), .cin({\g2[5][63] , \g2[5][62] , 
        \g2[5][61] , \g2[5][60] , \g2[5][59] , \g2[5][58] , \g2[5][57] , 
        \g2[5][56] , \g2[5][55] , \g2[5][54] , \g2[5][53] , \g2[5][52] , 
        \g2[5][51] , \g2[5][50] , \g2[5][49] , \g2[5][48] , \g2[5][47] , 
        \g2[5][46] , \g2[5][45] , \g2[5][44] , \g2[5][43] , \g2[5][42] , 
        \g2[5][41] , \g2[5][40] , \g2[5][39] , \g2[5][38] , \g2[5][37] , 
        \g2[5][36] , \g2[5][35] , \g2[5][34] , \g2[5][33] , \g2[5][32] , 
        \g2[5][31] , \g2[5][30] , \g2[5][29] , \g2[5][28] , \g2[5][27] , 
        \g2[5][26] , \g2[5][25] , \g2[5][24] , \g2[5][23] , \g2[5][22] , 
        \g2[5][21] , \g2[5][20] , \g2[5][19] , \g2[5][18] , \g2[5][17] , 
        \g2[5][16] , \g2[5][15] , \g2[5][14] , \g2[5][13] , \g2[5][12] , 
        \g2[5][11] , \g2[5][10] , \g2[5][9] , \g2[5][8] , \g2[5][7] , 
        \g2[5][6] , \g2[5][5] , \g2[5][4] , \g2[5][3] , \g2[5][2] , \g2[5][1] , 
        \g2[5][0] }), .sum({\g3[1][63] , \g3[1][62] , \g3[1][61] , \g3[1][60] , 
        \g3[1][59] , \g3[1][58] , \g3[1][57] , \g3[1][56] , \g3[1][55] , 
        \g3[1][54] , \g3[1][53] , \g3[1][52] , \g3[1][51] , \g3[1][50] , 
        \g3[1][49] , \g3[1][48] , \g3[1][47] , \g3[1][46] , \g3[1][45] , 
        \g3[1][44] , \g3[1][43] , \g3[1][42] , \g3[1][41] , \g3[1][40] , 
        \g3[1][39] , \g3[1][38] , \g3[1][37] , \g3[1][36] , \g3[1][35] , 
        \g3[1][34] , \g3[1][33] , \g3[1][32] , \g3[1][31] , \g3[1][30] , 
        \g3[1][29] , \g3[1][28] , \g3[1][27] , \g3[1][26] , \g3[1][25] , 
        \g3[1][24] , \g3[1][23] , \g3[1][22] , \g3[1][21] , \g3[1][20] , 
        \g3[1][19] , \g3[1][18] , \g3[1][17] , \g3[1][16] , \g3[1][15] , 
        \g3[1][14] , \g3[1][13] , \g3[1][12] , \g3[1][11] , \g3[1][10] , 
        \g3[1][9] , \g3[1][8] , \g3[1][7] , \g3[1][6] , \g3[1][5] , \g3[1][4] , 
        \g3[1][3] , \g3[1][2] , \g3[1][1] , \g3[1][0] }), .cout({\g3[10][63] , 
        \g3[10][62] , \g3[10][61] , \g3[10][60] , \g3[10][59] , \g3[10][58] , 
        \g3[10][57] , \g3[10][56] , \g3[10][55] , \g3[10][54] , \g3[10][53] , 
        \g3[10][52] , \g3[10][51] , \g3[10][50] , \g3[10][49] , \g3[10][48] , 
        \g3[10][47] , \g3[10][46] , \g3[10][45] , \g3[10][44] , \g3[10][43] , 
        \g3[10][42] , \g3[10][41] , \g3[10][40] , \g3[10][39] , \g3[10][38] , 
        \g3[10][37] , \g3[10][36] , \g3[10][35] , \g3[10][34] , \g3[10][33] , 
        \g3[10][32] , \g3[10][31] , \g3[10][30] , \g3[10][29] , \g3[10][28] , 
        \g3[10][27] , \g3[10][26] , \g3[10][25] , \g3[10][24] , \g3[10][23] , 
        \g3[10][22] , \g3[10][21] , \g3[10][20] , \g3[10][19] , \g3[10][18] , 
        \g3[10][17] , \g3[10][16] , \g3[10][15] , \g3[10][14] , \g3[10][13] , 
        \g3[10][12] , \g3[10][11] , \g3[10][10] , \g3[10][9] , \g3[10][8] , 
        \g3[10][7] , \g3[10][6] , \g3[10][5] , \g3[10][4] , \g3[10][3] , 
        \g3[10][2] , \g3[10][1] , SYNOPSYS_UNCONNECTED__36}) );
  FullAdder_25 \level3[2].x0  ( .a({\g2[6][63] , \g2[6][62] , \g2[6][61] , 
        \g2[6][60] , \g2[6][59] , \g2[6][58] , \g2[6][57] , \g2[6][56] , 
        \g2[6][55] , \g2[6][54] , \g2[6][53] , \g2[6][52] , \g2[6][51] , 
        \g2[6][50] , \g2[6][49] , \g2[6][48] , \g2[6][47] , \g2[6][46] , 
        \g2[6][45] , \g2[6][44] , \g2[6][43] , \g2[6][42] , \g2[6][41] , 
        \g2[6][40] , \g2[6][39] , \g2[6][38] , \g2[6][37] , \g2[6][36] , 
        \g2[6][35] , \g2[6][34] , \g2[6][33] , \g2[6][32] , \g2[6][31] , 
        \g2[6][30] , \g2[6][29] , \g2[6][28] , \g2[6][27] , \g2[6][26] , 
        \g2[6][25] , \g2[6][24] , \g2[6][23] , \g2[6][22] , \g2[6][21] , 
        \g2[6][20] , \g2[6][19] , \g2[6][18] , \g2[6][17] , \g2[6][16] , 
        \g2[6][15] , \g2[6][14] , \g2[6][13] , \g2[6][12] , \g2[6][11] , 
        \g2[6][10] , \g2[6][9] , \g2[6][8] , \g2[6][7] , \g2[6][6] , 
        \g2[6][5] , \g2[6][4] , \g2[6][3] , \g2[6][2] , \g2[6][1] , \g2[6][0] }), .b({\g2[7][63] , \g2[7][62] , \g2[7][61] , \g2[7][60] , \g2[7][59] , 
        \g2[7][58] , \g2[7][57] , \g2[7][56] , \g2[7][55] , \g2[7][54] , 
        \g2[7][53] , \g2[7][52] , \g2[7][51] , \g2[7][50] , \g2[7][49] , 
        \g2[7][48] , \g2[7][47] , \g2[7][46] , \g2[7][45] , \g2[7][44] , 
        \g2[7][43] , \g2[7][42] , \g2[7][41] , \g2[7][40] , \g2[7][39] , 
        \g2[7][38] , \g2[7][37] , \g2[7][36] , \g2[7][35] , \g2[7][34] , 
        \g2[7][33] , \g2[7][32] , \g2[7][31] , \g2[7][30] , \g2[7][29] , 
        \g2[7][28] , \g2[7][27] , \g2[7][26] , \g2[7][25] , \g2[7][24] , 
        \g2[7][23] , \g2[7][22] , \g2[7][21] , \g2[7][20] , \g2[7][19] , 
        \g2[7][18] , \g2[7][17] , \g2[7][16] , \g2[7][15] , \g2[7][14] , 
        \g2[7][13] , \g2[7][12] , \g2[7][11] , \g2[7][10] , \g2[7][9] , 
        \g2[7][8] , \g2[7][7] , \g2[7][6] , \g2[7][5] , \g2[7][4] , \g2[7][3] , 
        \g2[7][2] , \g2[7][1] , \g2[7][0] }), .cin({\g2[8][63] , \g2[8][62] , 
        \g2[8][61] , \g2[8][60] , \g2[8][59] , \g2[8][58] , \g2[8][57] , 
        \g2[8][56] , \g2[8][55] , \g2[8][54] , \g2[8][53] , \g2[8][52] , 
        \g2[8][51] , \g2[8][50] , \g2[8][49] , \g2[8][48] , \g2[8][47] , 
        \g2[8][46] , \g2[8][45] , \g2[8][44] , \g2[8][43] , \g2[8][42] , 
        \g2[8][41] , \g2[8][40] , \g2[8][39] , \g2[8][38] , \g2[8][37] , 
        \g2[8][36] , \g2[8][35] , \g2[8][34] , \g2[8][33] , \g2[8][32] , 
        \g2[8][31] , \g2[8][30] , \g2[8][29] , \g2[8][28] , \g2[8][27] , 
        \g2[8][26] , \g2[8][25] , \g2[8][24] , \g2[8][23] , \g2[8][22] , 
        \g2[8][21] , \g2[8][20] , \g2[8][19] , \g2[8][18] , \g2[8][17] , 
        \g2[8][16] , \g2[8][15] , \g2[8][14] , \g2[8][13] , \g2[8][12] , 
        \g2[8][11] , \g2[8][10] , \g2[8][9] , \g2[8][8] , \g2[8][7] , 
        \g2[8][6] , \g2[8][5] , \g2[8][4] , \g2[8][3] , \g2[8][2] , \g2[8][1] , 
        \g2[8][0] }), .sum({\g3[2][63] , \g3[2][62] , \g3[2][61] , \g3[2][60] , 
        \g3[2][59] , \g3[2][58] , \g3[2][57] , \g3[2][56] , \g3[2][55] , 
        \g3[2][54] , \g3[2][53] , \g3[2][52] , \g3[2][51] , \g3[2][50] , 
        \g3[2][49] , \g3[2][48] , \g3[2][47] , \g3[2][46] , \g3[2][45] , 
        \g3[2][44] , \g3[2][43] , \g3[2][42] , \g3[2][41] , \g3[2][40] , 
        \g3[2][39] , \g3[2][38] , \g3[2][37] , \g3[2][36] , \g3[2][35] , 
        \g3[2][34] , \g3[2][33] , \g3[2][32] , \g3[2][31] , \g3[2][30] , 
        \g3[2][29] , \g3[2][28] , \g3[2][27] , \g3[2][26] , \g3[2][25] , 
        \g3[2][24] , \g3[2][23] , \g3[2][22] , \g3[2][21] , \g3[2][20] , 
        \g3[2][19] , \g3[2][18] , \g3[2][17] , \g3[2][16] , \g3[2][15] , 
        \g3[2][14] , \g3[2][13] , \g3[2][12] , \g3[2][11] , \g3[2][10] , 
        \g3[2][9] , \g3[2][8] , \g3[2][7] , \g3[2][6] , \g3[2][5] , \g3[2][4] , 
        \g3[2][3] , \g3[2][2] , \g3[2][1] , \g3[2][0] }), .cout({\g3[11][63] , 
        \g3[11][62] , \g3[11][61] , \g3[11][60] , \g3[11][59] , \g3[11][58] , 
        \g3[11][57] , \g3[11][56] , \g3[11][55] , \g3[11][54] , \g3[11][53] , 
        \g3[11][52] , \g3[11][51] , \g3[11][50] , \g3[11][49] , \g3[11][48] , 
        \g3[11][47] , \g3[11][46] , \g3[11][45] , \g3[11][44] , \g3[11][43] , 
        \g3[11][42] , \g3[11][41] , \g3[11][40] , \g3[11][39] , \g3[11][38] , 
        \g3[11][37] , \g3[11][36] , \g3[11][35] , \g3[11][34] , \g3[11][33] , 
        \g3[11][32] , \g3[11][31] , \g3[11][30] , \g3[11][29] , \g3[11][28] , 
        \g3[11][27] , \g3[11][26] , \g3[11][25] , \g3[11][24] , \g3[11][23] , 
        \g3[11][22] , \g3[11][21] , \g3[11][20] , \g3[11][19] , \g3[11][18] , 
        \g3[11][17] , \g3[11][16] , \g3[11][15] , \g3[11][14] , \g3[11][13] , 
        \g3[11][12] , \g3[11][11] , \g3[11][10] , \g3[11][9] , \g3[11][8] , 
        \g3[11][7] , \g3[11][6] , \g3[11][5] , \g3[11][4] , \g3[11][3] , 
        \g3[11][2] , \g3[11][1] , SYNOPSYS_UNCONNECTED__37}) );
  FullAdder_24 \level3[3].x0  ( .a({\g2[9][63] , \g2[9][62] , \g2[9][61] , 
        \g2[9][60] , \g2[9][59] , \g2[9][58] , \g2[9][57] , \g2[9][56] , 
        \g2[9][55] , \g2[9][54] , \g2[9][53] , \g2[9][52] , \g2[9][51] , 
        \g2[9][50] , \g2[9][49] , \g2[9][48] , \g2[9][47] , \g2[9][46] , 
        \g2[9][45] , \g2[9][44] , \g2[9][43] , \g2[9][42] , \g2[9][41] , 
        \g2[9][40] , \g2[9][39] , \g2[9][38] , \g2[9][37] , \g2[9][36] , 
        \g2[9][35] , \g2[9][34] , \g2[9][33] , \g2[9][32] , \g2[9][31] , 
        \g2[9][30] , \g2[9][29] , \g2[9][28] , \g2[9][27] , \g2[9][26] , 
        \g2[9][25] , \g2[9][24] , \g2[9][23] , \g2[9][22] , \g2[9][21] , 
        \g2[9][20] , \g2[9][19] , \g2[9][18] , \g2[9][17] , \g2[9][16] , 
        \g2[9][15] , \g2[9][14] , \g2[9][13] , \g2[9][12] , \g2[9][11] , 
        \g2[9][10] , \g2[9][9] , \g2[9][8] , \g2[9][7] , \g2[9][6] , 
        \g2[9][5] , \g2[9][4] , \g2[9][3] , \g2[9][2] , \g2[9][1] , \g2[9][0] }), .b({\g2[10][63] , \g2[10][62] , \g2[10][61] , \g2[10][60] , \g2[10][59] , 
        \g2[10][58] , \g2[10][57] , \g2[10][56] , \g2[10][55] , \g2[10][54] , 
        \g2[10][53] , \g2[10][52] , \g2[10][51] , \g2[10][50] , \g2[10][49] , 
        \g2[10][48] , \g2[10][47] , \g2[10][46] , \g2[10][45] , \g2[10][44] , 
        \g2[10][43] , \g2[10][42] , \g2[10][41] , \g2[10][40] , \g2[10][39] , 
        \g2[10][38] , \g2[10][37] , \g2[10][36] , \g2[10][35] , \g2[10][34] , 
        \g2[10][33] , \g2[10][32] , \g2[10][31] , \g2[10][30] , \g2[10][29] , 
        \g2[10][28] , \g2[10][27] , \g2[10][26] , \g2[10][25] , \g2[10][24] , 
        \g2[10][23] , \g2[10][22] , \g2[10][21] , \g2[10][20] , \g2[10][19] , 
        \g2[10][18] , \g2[10][17] , \g2[10][16] , \g2[10][15] , \g2[10][14] , 
        \g2[10][13] , \g2[10][12] , \g2[10][11] , \g2[10][10] , \g2[10][9] , 
        \g2[10][8] , \g2[10][7] , \g2[10][6] , \g2[10][5] , \g2[10][4] , 
        \g2[10][3] , \g2[10][2] , \g2[10][1] , \g2[10][0] }), .cin({
        \g2[11][63] , \g2[11][62] , \g2[11][61] , \g2[11][60] , \g2[11][59] , 
        \g2[11][58] , \g2[11][57] , \g2[11][56] , \g2[11][55] , \g2[11][54] , 
        \g2[11][53] , \g2[11][52] , \g2[11][51] , \g2[11][50] , \g2[11][49] , 
        \g2[11][48] , \g2[11][47] , \g2[11][46] , \g2[11][45] , \g2[11][44] , 
        \g2[11][43] , \g2[11][42] , \g2[11][41] , \g2[11][40] , \g2[11][39] , 
        \g2[11][38] , \g2[11][37] , \g2[11][36] , \g2[11][35] , \g2[11][34] , 
        \g2[11][33] , \g2[11][32] , \g2[11][31] , \g2[11][30] , \g2[11][29] , 
        \g2[11][28] , \g2[11][27] , \g2[11][26] , \g2[11][25] , \g2[11][24] , 
        \g2[11][23] , \g2[11][22] , \g2[11][21] , \g2[11][20] , \g2[11][19] , 
        \g2[11][18] , \g2[11][17] , \g2[11][16] , \g2[11][15] , \g2[11][14] , 
        \g2[11][13] , \g2[11][12] , \g2[11][11] , \g2[11][10] , \g2[11][9] , 
        \g2[11][8] , \g2[11][7] , \g2[11][6] , \g2[11][5] , \g2[11][4] , 
        \g2[11][3] , \g2[11][2] , \g2[11][1] , \g2[11][0] }), .sum({
        \g3[3][63] , \g3[3][62] , \g3[3][61] , \g3[3][60] , \g3[3][59] , 
        \g3[3][58] , \g3[3][57] , \g3[3][56] , \g3[3][55] , \g3[3][54] , 
        \g3[3][53] , \g3[3][52] , \g3[3][51] , \g3[3][50] , \g3[3][49] , 
        \g3[3][48] , \g3[3][47] , \g3[3][46] , \g3[3][45] , \g3[3][44] , 
        \g3[3][43] , \g3[3][42] , \g3[3][41] , \g3[3][40] , \g3[3][39] , 
        \g3[3][38] , \g3[3][37] , \g3[3][36] , \g3[3][35] , \g3[3][34] , 
        \g3[3][33] , \g3[3][32] , \g3[3][31] , \g3[3][30] , \g3[3][29] , 
        \g3[3][28] , \g3[3][27] , \g3[3][26] , \g3[3][25] , \g3[3][24] , 
        \g3[3][23] , \g3[3][22] , \g3[3][21] , \g3[3][20] , \g3[3][19] , 
        \g3[3][18] , \g3[3][17] , \g3[3][16] , \g3[3][15] , \g3[3][14] , 
        \g3[3][13] , \g3[3][12] , \g3[3][11] , \g3[3][10] , \g3[3][9] , 
        \g3[3][8] , \g3[3][7] , \g3[3][6] , \g3[3][5] , \g3[3][4] , \g3[3][3] , 
        \g3[3][2] , \g3[3][1] , \g3[3][0] }), .cout({\g3[12][63] , 
        \g3[12][62] , \g3[12][61] , \g3[12][60] , \g3[12][59] , \g3[12][58] , 
        \g3[12][57] , \g3[12][56] , \g3[12][55] , \g3[12][54] , \g3[12][53] , 
        \g3[12][52] , \g3[12][51] , \g3[12][50] , \g3[12][49] , \g3[12][48] , 
        \g3[12][47] , \g3[12][46] , \g3[12][45] , \g3[12][44] , \g3[12][43] , 
        \g3[12][42] , \g3[12][41] , \g3[12][40] , \g3[12][39] , \g3[12][38] , 
        \g3[12][37] , \g3[12][36] , \g3[12][35] , \g3[12][34] , \g3[12][33] , 
        \g3[12][32] , \g3[12][31] , \g3[12][30] , \g3[12][29] , \g3[12][28] , 
        \g3[12][27] , \g3[12][26] , \g3[12][25] , \g3[12][24] , \g3[12][23] , 
        \g3[12][22] , \g3[12][21] , \g3[12][20] , \g3[12][19] , \g3[12][18] , 
        \g3[12][17] , \g3[12][16] , \g3[12][15] , \g3[12][14] , \g3[12][13] , 
        \g3[12][12] , \g3[12][11] , \g3[12][10] , \g3[12][9] , \g3[12][8] , 
        \g3[12][7] , \g3[12][6] , \g3[12][5] , \g3[12][4] , \g3[12][3] , 
        \g3[12][2] , \g3[12][1] , SYNOPSYS_UNCONNECTED__38}) );
  FullAdder_23 \level3[4].x0  ( .a({\g2[12][63] , \g2[12][62] , \g2[12][61] , 
        \g2[12][60] , \g2[12][59] , \g2[12][58] , \g2[12][57] , \g2[12][56] , 
        \g2[12][55] , \g2[12][54] , \g2[12][53] , \g2[12][52] , \g2[12][51] , 
        \g2[12][50] , \g2[12][49] , \g2[12][48] , \g2[12][47] , \g2[12][46] , 
        \g2[12][45] , \g2[12][44] , \g2[12][43] , \g2[12][42] , \g2[12][41] , 
        \g2[12][40] , \g2[12][39] , \g2[12][38] , \g2[12][37] , \g2[12][36] , 
        \g2[12][35] , \g2[12][34] , \g2[12][33] , \g2[12][32] , \g2[12][31] , 
        \g2[12][30] , \g2[12][29] , \g2[12][28] , \g2[12][27] , \g2[12][26] , 
        \g2[12][25] , \g2[12][24] , \g2[12][23] , \g2[12][22] , \g2[12][21] , 
        \g2[12][20] , \g2[12][19] , \g2[12][18] , \g2[12][17] , \g2[12][16] , 
        \g2[12][15] , \g2[12][14] , \g2[12][13] , \g2[12][12] , \g2[12][11] , 
        \g2[12][10] , \g2[12][9] , \g2[12][8] , \g2[12][7] , \g2[12][6] , 
        \g2[12][5] , \g2[12][4] , \g2[12][3] , \g2[12][2] , \g2[12][1] , 
        \g2[12][0] }), .b({\g2[13][63] , \g2[13][62] , \g2[13][61] , 
        \g2[13][60] , \g2[13][59] , \g2[13][58] , \g2[13][57] , \g2[13][56] , 
        \g2[13][55] , \g2[13][54] , \g2[13][53] , \g2[13][52] , \g2[13][51] , 
        \g2[13][50] , \g2[13][49] , \g2[13][48] , \g2[13][47] , \g2[13][46] , 
        \g2[13][45] , \g2[13][44] , \g2[13][43] , \g2[13][42] , \g2[13][41] , 
        \g2[13][40] , \g2[13][39] , \g2[13][38] , \g2[13][37] , \g2[13][36] , 
        \g2[13][35] , \g2[13][34] , \g2[13][33] , \g2[13][32] , \g2[13][31] , 
        \g2[13][30] , \g2[13][29] , \g2[13][28] , \g2[13][27] , \g2[13][26] , 
        \g2[13][25] , \g2[13][24] , \g2[13][23] , \g2[13][22] , \g2[13][21] , 
        \g2[13][20] , \g2[13][19] , \g2[13][18] , \g2[13][17] , \g2[13][16] , 
        \g2[13][15] , \g2[13][14] , \g2[13][13] , \g2[13][12] , \g2[13][11] , 
        \g2[13][10] , \g2[13][9] , \g2[13][8] , \g2[13][7] , \g2[13][6] , 
        \g2[13][5] , \g2[13][4] , \g2[13][3] , \g2[13][2] , \g2[13][1] , 
        \g2[13][0] }), .cin({\g2[14][63] , \g2[14][62] , \g2[14][61] , 
        \g2[14][60] , \g2[14][59] , \g2[14][58] , \g2[14][57] , \g2[14][56] , 
        \g2[14][55] , \g2[14][54] , \g2[14][53] , \g2[14][52] , \g2[14][51] , 
        \g2[14][50] , \g2[14][49] , \g2[14][48] , \g2[14][47] , \g2[14][46] , 
        \g2[14][45] , \g2[14][44] , \g2[14][43] , \g2[14][42] , \g2[14][41] , 
        \g2[14][40] , \g2[14][39] , \g2[14][38] , \g2[14][37] , \g2[14][36] , 
        \g2[14][35] , \g2[14][34] , \g2[14][33] , \g2[14][32] , \g2[14][31] , 
        \g2[14][30] , \g2[14][29] , \g2[14][28] , \g2[14][27] , \g2[14][26] , 
        \g2[14][25] , \g2[14][24] , \g2[14][23] , \g2[14][22] , \g2[14][21] , 
        \g2[14][20] , \g2[14][19] , \g2[14][18] , \g2[14][17] , \g2[14][16] , 
        \g2[14][15] , \g2[14][14] , \g2[14][13] , \g2[14][12] , \g2[14][11] , 
        \g2[14][10] , \g2[14][9] , \g2[14][8] , \g2[14][7] , \g2[14][6] , 
        \g2[14][5] , \g2[14][4] , \g2[14][3] , \g2[14][2] , \g2[14][1] , 1'b0}), .sum({\g3[4][63] , \g3[4][62] , \g3[4][61] , \g3[4][60] , \g3[4][59] , 
        \g3[4][58] , \g3[4][57] , \g3[4][56] , \g3[4][55] , \g3[4][54] , 
        \g3[4][53] , \g3[4][52] , \g3[4][51] , \g3[4][50] , \g3[4][49] , 
        \g3[4][48] , \g3[4][47] , \g3[4][46] , \g3[4][45] , \g3[4][44] , 
        \g3[4][43] , \g3[4][42] , \g3[4][41] , \g3[4][40] , \g3[4][39] , 
        \g3[4][38] , \g3[4][37] , \g3[4][36] , \g3[4][35] , \g3[4][34] , 
        \g3[4][33] , \g3[4][32] , \g3[4][31] , \g3[4][30] , \g3[4][29] , 
        \g3[4][28] , \g3[4][27] , \g3[4][26] , \g3[4][25] , \g3[4][24] , 
        \g3[4][23] , \g3[4][22] , \g3[4][21] , \g3[4][20] , \g3[4][19] , 
        \g3[4][18] , \g3[4][17] , \g3[4][16] , \g3[4][15] , \g3[4][14] , 
        \g3[4][13] , \g3[4][12] , \g3[4][11] , \g3[4][10] , \g3[4][9] , 
        \g3[4][8] , \g3[4][7] , \g3[4][6] , \g3[4][5] , \g3[4][4] , \g3[4][3] , 
        \g3[4][2] , \g3[4][1] , \g3[4][0] }), .cout({\g3[13][63] , 
        \g3[13][62] , \g3[13][61] , \g3[13][60] , \g3[13][59] , \g3[13][58] , 
        \g3[13][57] , \g3[13][56] , \g3[13][55] , \g3[13][54] , \g3[13][53] , 
        \g3[13][52] , \g3[13][51] , \g3[13][50] , \g3[13][49] , \g3[13][48] , 
        \g3[13][47] , \g3[13][46] , \g3[13][45] , \g3[13][44] , \g3[13][43] , 
        \g3[13][42] , \g3[13][41] , \g3[13][40] , \g3[13][39] , \g3[13][38] , 
        \g3[13][37] , \g3[13][36] , \g3[13][35] , \g3[13][34] , \g3[13][33] , 
        \g3[13][32] , \g3[13][31] , \g3[13][30] , \g3[13][29] , \g3[13][28] , 
        \g3[13][27] , \g3[13][26] , \g3[13][25] , \g3[13][24] , \g3[13][23] , 
        \g3[13][22] , \g3[13][21] , \g3[13][20] , \g3[13][19] , \g3[13][18] , 
        \g3[13][17] , \g3[13][16] , \g3[13][15] , \g3[13][14] , \g3[13][13] , 
        \g3[13][12] , \g3[13][11] , \g3[13][10] , \g3[13][9] , \g3[13][8] , 
        \g3[13][7] , \g3[13][6] , \g3[13][5] , \g3[13][4] , \g3[13][3] , 
        \g3[13][2] , \g3[13][1] , SYNOPSYS_UNCONNECTED__39}) );
  FullAdder_22 \level3[5].x0  ( .a({\g2[15][63] , \g2[15][62] , \g2[15][61] , 
        \g2[15][60] , \g2[15][59] , \g2[15][58] , \g2[15][57] , \g2[15][56] , 
        \g2[15][55] , \g2[15][54] , \g2[15][53] , \g2[15][52] , \g2[15][51] , 
        \g2[15][50] , \g2[15][49] , \g2[15][48] , \g2[15][47] , \g2[15][46] , 
        \g2[15][45] , \g2[15][44] , \g2[15][43] , \g2[15][42] , \g2[15][41] , 
        \g2[15][40] , \g2[15][39] , \g2[15][38] , \g2[15][37] , \g2[15][36] , 
        \g2[15][35] , \g2[15][34] , \g2[15][33] , \g2[15][32] , \g2[15][31] , 
        \g2[15][30] , \g2[15][29] , \g2[15][28] , \g2[15][27] , \g2[15][26] , 
        \g2[15][25] , \g2[15][24] , \g2[15][23] , \g2[15][22] , \g2[15][21] , 
        \g2[15][20] , \g2[15][19] , \g2[15][18] , \g2[15][17] , \g2[15][16] , 
        \g2[15][15] , \g2[15][14] , \g2[15][13] , \g2[15][12] , \g2[15][11] , 
        \g2[15][10] , \g2[15][9] , \g2[15][8] , \g2[15][7] , \g2[15][6] , 
        \g2[15][5] , \g2[15][4] , \g2[15][3] , \g2[15][2] , \g2[15][1] , 1'b0}), .b({\g2[16][63] , \g2[16][62] , \g2[16][61] , \g2[16][60] , \g2[16][59] , 
        \g2[16][58] , \g2[16][57] , \g2[16][56] , \g2[16][55] , \g2[16][54] , 
        \g2[16][53] , \g2[16][52] , \g2[16][51] , \g2[16][50] , \g2[16][49] , 
        \g2[16][48] , \g2[16][47] , \g2[16][46] , \g2[16][45] , \g2[16][44] , 
        \g2[16][43] , \g2[16][42] , \g2[16][41] , \g2[16][40] , \g2[16][39] , 
        \g2[16][38] , \g2[16][37] , \g2[16][36] , \g2[16][35] , \g2[16][34] , 
        \g2[16][33] , \g2[16][32] , \g2[16][31] , \g2[16][30] , \g2[16][29] , 
        \g2[16][28] , \g2[16][27] , \g2[16][26] , \g2[16][25] , \g2[16][24] , 
        \g2[16][23] , \g2[16][22] , \g2[16][21] , \g2[16][20] , \g2[16][19] , 
        \g2[16][18] , \g2[16][17] , \g2[16][16] , \g2[16][15] , \g2[16][14] , 
        \g2[16][13] , \g2[16][12] , \g2[16][11] , \g2[16][10] , \g2[16][9] , 
        \g2[16][8] , \g2[16][7] , \g2[16][6] , \g2[16][5] , \g2[16][4] , 
        \g2[16][3] , \g2[16][2] , \g2[16][1] , 1'b0}), .cin({\g2[17][63] , 
        \g2[17][62] , \g2[17][61] , \g2[17][60] , \g2[17][59] , \g2[17][58] , 
        \g2[17][57] , \g2[17][56] , \g2[17][55] , \g2[17][54] , \g2[17][53] , 
        \g2[17][52] , \g2[17][51] , \g2[17][50] , \g2[17][49] , \g2[17][48] , 
        \g2[17][47] , \g2[17][46] , \g2[17][45] , \g2[17][44] , \g2[17][43] , 
        \g2[17][42] , \g2[17][41] , \g2[17][40] , \g2[17][39] , \g2[17][38] , 
        \g2[17][37] , \g2[17][36] , \g2[17][35] , \g2[17][34] , \g2[17][33] , 
        \g2[17][32] , \g2[17][31] , \g2[17][30] , \g2[17][29] , \g2[17][28] , 
        \g2[17][27] , \g2[17][26] , \g2[17][25] , \g2[17][24] , \g2[17][23] , 
        \g2[17][22] , \g2[17][21] , \g2[17][20] , \g2[17][19] , \g2[17][18] , 
        \g2[17][17] , \g2[17][16] , \g2[17][15] , \g2[17][14] , \g2[17][13] , 
        \g2[17][12] , \g2[17][11] , \g2[17][10] , \g2[17][9] , \g2[17][8] , 
        \g2[17][7] , \g2[17][6] , \g2[17][5] , \g2[17][4] , \g2[17][3] , 
        \g2[17][2] , \g2[17][1] , 1'b0}), .sum({\g3[5][63] , \g3[5][62] , 
        \g3[5][61] , \g3[5][60] , \g3[5][59] , \g3[5][58] , \g3[5][57] , 
        \g3[5][56] , \g3[5][55] , \g3[5][54] , \g3[5][53] , \g3[5][52] , 
        \g3[5][51] , \g3[5][50] , \g3[5][49] , \g3[5][48] , \g3[5][47] , 
        \g3[5][46] , \g3[5][45] , \g3[5][44] , \g3[5][43] , \g3[5][42] , 
        \g3[5][41] , \g3[5][40] , \g3[5][39] , \g3[5][38] , \g3[5][37] , 
        \g3[5][36] , \g3[5][35] , \g3[5][34] , \g3[5][33] , \g3[5][32] , 
        \g3[5][31] , \g3[5][30] , \g3[5][29] , \g3[5][28] , \g3[5][27] , 
        \g3[5][26] , \g3[5][25] , \g3[5][24] , \g3[5][23] , \g3[5][22] , 
        \g3[5][21] , \g3[5][20] , \g3[5][19] , \g3[5][18] , \g3[5][17] , 
        \g3[5][16] , \g3[5][15] , \g3[5][14] , \g3[5][13] , \g3[5][12] , 
        \g3[5][11] , \g3[5][10] , \g3[5][9] , \g3[5][8] , \g3[5][7] , 
        \g3[5][6] , \g3[5][5] , \g3[5][4] , \g3[5][3] , \g3[5][2] , \g3[5][1] , 
        \g3[5][0] }), .cout({\g3[14][63] , \g3[14][62] , \g3[14][61] , 
        \g3[14][60] , \g3[14][59] , \g3[14][58] , \g3[14][57] , \g3[14][56] , 
        \g3[14][55] , \g3[14][54] , \g3[14][53] , \g3[14][52] , \g3[14][51] , 
        \g3[14][50] , \g3[14][49] , \g3[14][48] , \g3[14][47] , \g3[14][46] , 
        \g3[14][45] , \g3[14][44] , \g3[14][43] , \g3[14][42] , \g3[14][41] , 
        \g3[14][40] , \g3[14][39] , \g3[14][38] , \g3[14][37] , \g3[14][36] , 
        \g3[14][35] , \g3[14][34] , \g3[14][33] , \g3[14][32] , \g3[14][31] , 
        \g3[14][30] , \g3[14][29] , \g3[14][28] , \g3[14][27] , \g3[14][26] , 
        \g3[14][25] , \g3[14][24] , \g3[14][23] , \g3[14][22] , \g3[14][21] , 
        \g3[14][20] , \g3[14][19] , \g3[14][18] , \g3[14][17] , \g3[14][16] , 
        \g3[14][15] , \g3[14][14] , \g3[14][13] , \g3[14][12] , \g3[14][11] , 
        \g3[14][10] , \g3[14][9] , \g3[14][8] , \g3[14][7] , \g3[14][6] , 
        \g3[14][5] , \g3[14][4] , \g3[14][3] , \g3[14][2] , \g3[14][1] , 
        SYNOPSYS_UNCONNECTED__40}) );
  FullAdder_21 \level3[6].x0  ( .a({\g2[18][63] , \g2[18][62] , \g2[18][61] , 
        \g2[18][60] , \g2[18][59] , \g2[18][58] , \g2[18][57] , \g2[18][56] , 
        \g2[18][55] , \g2[18][54] , \g2[18][53] , \g2[18][52] , \g2[18][51] , 
        \g2[18][50] , \g2[18][49] , \g2[18][48] , \g2[18][47] , \g2[18][46] , 
        \g2[18][45] , \g2[18][44] , \g2[18][43] , \g2[18][42] , \g2[18][41] , 
        \g2[18][40] , \g2[18][39] , \g2[18][38] , \g2[18][37] , \g2[18][36] , 
        \g2[18][35] , \g2[18][34] , \g2[18][33] , \g2[18][32] , \g2[18][31] , 
        \g2[18][30] , \g2[18][29] , \g2[18][28] , \g2[18][27] , \g2[18][26] , 
        \g2[18][25] , \g2[18][24] , \g2[18][23] , \g2[18][22] , \g2[18][21] , 
        \g2[18][20] , \g2[18][19] , \g2[18][18] , \g2[18][17] , \g2[18][16] , 
        \g2[18][15] , \g2[18][14] , \g2[18][13] , \g2[18][12] , \g2[18][11] , 
        \g2[18][10] , \g2[18][9] , \g2[18][8] , \g2[18][7] , \g2[18][6] , 
        \g2[18][5] , \g2[18][4] , \g2[18][3] , \g2[18][2] , \g2[18][1] , 1'b0}), .b({\g2[19][63] , \g2[19][62] , \g2[19][61] , \g2[19][60] , \g2[19][59] , 
        \g2[19][58] , \g2[19][57] , \g2[19][56] , \g2[19][55] , \g2[19][54] , 
        \g2[19][53] , \g2[19][52] , \g2[19][51] , \g2[19][50] , \g2[19][49] , 
        \g2[19][48] , \g2[19][47] , \g2[19][46] , \g2[19][45] , \g2[19][44] , 
        \g2[19][43] , \g2[19][42] , \g2[19][41] , \g2[19][40] , \g2[19][39] , 
        \g2[19][38] , \g2[19][37] , \g2[19][36] , \g2[19][35] , \g2[19][34] , 
        \g2[19][33] , \g2[19][32] , \g2[19][31] , \g2[19][30] , \g2[19][29] , 
        \g2[19][28] , \g2[19][27] , \g2[19][26] , \g2[19][25] , \g2[19][24] , 
        \g2[19][23] , \g2[19][22] , \g2[19][21] , \g2[19][20] , \g2[19][19] , 
        \g2[19][18] , \g2[19][17] , \g2[19][16] , \g2[19][15] , \g2[19][14] , 
        \g2[19][13] , \g2[19][12] , \g2[19][11] , \g2[19][10] , \g2[19][9] , 
        \g2[19][8] , \g2[19][7] , \g2[19][6] , \g2[19][5] , \g2[19][4] , 
        \g2[19][3] , \g2[19][2] , \g2[19][1] , 1'b0}), .cin({\g2[20][63] , 
        \g2[20][62] , \g2[20][61] , \g2[20][60] , \g2[20][59] , \g2[20][58] , 
        \g2[20][57] , \g2[20][56] , \g2[20][55] , \g2[20][54] , \g2[20][53] , 
        \g2[20][52] , \g2[20][51] , \g2[20][50] , \g2[20][49] , \g2[20][48] , 
        \g2[20][47] , \g2[20][46] , \g2[20][45] , \g2[20][44] , \g2[20][43] , 
        \g2[20][42] , \g2[20][41] , \g2[20][40] , \g2[20][39] , \g2[20][38] , 
        \g2[20][37] , \g2[20][36] , \g2[20][35] , \g2[20][34] , \g2[20][33] , 
        \g2[20][32] , \g2[20][31] , \g2[20][30] , \g2[20][29] , \g2[20][28] , 
        \g2[20][27] , \g2[20][26] , \g2[20][25] , \g2[20][24] , \g2[20][23] , 
        \g2[20][22] , \g2[20][21] , \g2[20][20] , \g2[20][19] , \g2[20][18] , 
        \g2[20][17] , \g2[20][16] , \g2[20][15] , \g2[20][14] , \g2[20][13] , 
        \g2[20][12] , \g2[20][11] , \g2[20][10] , \g2[20][9] , \g2[20][8] , 
        \g2[20][7] , \g2[20][6] , \g2[20][5] , \g2[20][4] , \g2[20][3] , 
        \g2[20][2] , \g2[20][1] , 1'b0}), .sum({\g3[6][63] , \g3[6][62] , 
        \g3[6][61] , \g3[6][60] , \g3[6][59] , \g3[6][58] , \g3[6][57] , 
        \g3[6][56] , \g3[6][55] , \g3[6][54] , \g3[6][53] , \g3[6][52] , 
        \g3[6][51] , \g3[6][50] , \g3[6][49] , \g3[6][48] , \g3[6][47] , 
        \g3[6][46] , \g3[6][45] , \g3[6][44] , \g3[6][43] , \g3[6][42] , 
        \g3[6][41] , \g3[6][40] , \g3[6][39] , \g3[6][38] , \g3[6][37] , 
        \g3[6][36] , \g3[6][35] , \g3[6][34] , \g3[6][33] , \g3[6][32] , 
        \g3[6][31] , \g3[6][30] , \g3[6][29] , \g3[6][28] , \g3[6][27] , 
        \g3[6][26] , \g3[6][25] , \g3[6][24] , \g3[6][23] , \g3[6][22] , 
        \g3[6][21] , \g3[6][20] , \g3[6][19] , \g3[6][18] , \g3[6][17] , 
        \g3[6][16] , \g3[6][15] , \g3[6][14] , \g3[6][13] , \g3[6][12] , 
        \g3[6][11] , \g3[6][10] , \g3[6][9] , \g3[6][8] , \g3[6][7] , 
        \g3[6][6] , \g3[6][5] , \g3[6][4] , \g3[6][3] , \g3[6][2] , \g3[6][1] , 
        \g3[6][0] }), .cout({\g3[15][63] , \g3[15][62] , \g3[15][61] , 
        \g3[15][60] , \g3[15][59] , \g3[15][58] , \g3[15][57] , \g3[15][56] , 
        \g3[15][55] , \g3[15][54] , \g3[15][53] , \g3[15][52] , \g3[15][51] , 
        \g3[15][50] , \g3[15][49] , \g3[15][48] , \g3[15][47] , \g3[15][46] , 
        \g3[15][45] , \g3[15][44] , \g3[15][43] , \g3[15][42] , \g3[15][41] , 
        \g3[15][40] , \g3[15][39] , \g3[15][38] , \g3[15][37] , \g3[15][36] , 
        \g3[15][35] , \g3[15][34] , \g3[15][33] , \g3[15][32] , \g3[15][31] , 
        \g3[15][30] , \g3[15][29] , \g3[15][28] , \g3[15][27] , \g3[15][26] , 
        \g3[15][25] , \g3[15][24] , \g3[15][23] , \g3[15][22] , \g3[15][21] , 
        \g3[15][20] , \g3[15][19] , \g3[15][18] , \g3[15][17] , \g3[15][16] , 
        \g3[15][15] , \g3[15][14] , \g3[15][13] , \g3[15][12] , \g3[15][11] , 
        \g3[15][10] , \g3[15][9] , \g3[15][8] , \g3[15][7] , \g3[15][6] , 
        \g3[15][5] , \g3[15][4] , \g3[15][3] , \g3[15][2] , \g3[15][1] , 
        SYNOPSYS_UNCONNECTED__41}) );
  FullAdder_20 \level3[7].x0  ( .a({\g2[21][63] , \g2[21][62] , \g2[21][61] , 
        \g2[21][60] , \g2[21][59] , \g2[21][58] , \g2[21][57] , \g2[21][56] , 
        \g2[21][55] , \g2[21][54] , \g2[21][53] , \g2[21][52] , \g2[21][51] , 
        \g2[21][50] , \g2[21][49] , \g2[21][48] , \g2[21][47] , \g2[21][46] , 
        \g2[21][45] , \g2[21][44] , \g2[21][43] , \g2[21][42] , \g2[21][41] , 
        \g2[21][40] , \g2[21][39] , \g2[21][38] , \g2[21][37] , \g2[21][36] , 
        \g2[21][35] , \g2[21][34] , \g2[21][33] , \g2[21][32] , \g2[21][31] , 
        \g2[21][30] , \g2[21][29] , \g2[21][28] , \g2[21][27] , \g2[21][26] , 
        \g2[21][25] , \g2[21][24] , \g2[21][23] , \g2[21][22] , \g2[21][21] , 
        \g2[21][20] , \g2[21][19] , \g2[21][18] , \g2[21][17] , \g2[21][16] , 
        \g2[21][15] , \g2[21][14] , \g2[21][13] , \g2[21][12] , \g2[21][11] , 
        \g2[21][10] , \g2[21][9] , \g2[21][8] , \g2[21][7] , \g2[21][6] , 
        \g2[21][5] , \g2[21][4] , \g2[21][3] , \g2[21][2] , \g2[21][1] , 1'b0}), .b({\g2[22][63] , \g2[22][62] , \g2[22][61] , \g2[22][60] , \g2[22][59] , 
        \g2[22][58] , \g2[22][57] , \g2[22][56] , \g2[22][55] , \g2[22][54] , 
        \g2[22][53] , \g2[22][52] , \g2[22][51] , \g2[22][50] , \g2[22][49] , 
        \g2[22][48] , \g2[22][47] , \g2[22][46] , \g2[22][45] , \g2[22][44] , 
        \g2[22][43] , \g2[22][42] , \g2[22][41] , \g2[22][40] , \g2[22][39] , 
        \g2[22][38] , \g2[22][37] , \g2[22][36] , \g2[22][35] , \g2[22][34] , 
        \g2[22][33] , \g2[22][32] , \g2[22][31] , \g2[22][30] , \g2[22][29] , 
        \g2[22][28] , \g2[22][27] , \g2[22][26] , \g2[22][25] , \g2[22][24] , 
        \g2[22][23] , \g2[22][22] , \g2[22][21] , \g2[22][20] , \g2[22][19] , 
        \g2[22][18] , \g2[22][17] , \g2[22][16] , \g2[22][15] , \g2[22][14] , 
        \g2[22][13] , \g2[22][12] , \g2[22][11] , \g2[22][10] , \g2[22][9] , 
        \g2[22][8] , \g2[22][7] , \g2[22][6] , \g2[22][5] , \g2[22][4] , 
        \g2[22][3] , \g2[22][2] , \g2[22][1] , 1'b0}), .cin({\g2[23][63] , 
        \g2[23][62] , \g2[23][61] , \g2[23][60] , \g2[23][59] , \g2[23][58] , 
        \g2[23][57] , \g2[23][56] , \g2[23][55] , \g2[23][54] , \g2[23][53] , 
        \g2[23][52] , \g2[23][51] , \g2[23][50] , \g2[23][49] , \g2[23][48] , 
        \g2[23][47] , \g2[23][46] , \g2[23][45] , \g2[23][44] , \g2[23][43] , 
        \g2[23][42] , \g2[23][41] , \g2[23][40] , \g2[23][39] , \g2[23][38] , 
        \g2[23][37] , \g2[23][36] , \g2[23][35] , \g2[23][34] , \g2[23][33] , 
        \g2[23][32] , \g2[23][31] , \g2[23][30] , \g2[23][29] , \g2[23][28] , 
        \g2[23][27] , \g2[23][26] , \g2[23][25] , \g2[23][24] , \g2[23][23] , 
        \g2[23][22] , \g2[23][21] , \g2[23][20] , \g2[23][19] , \g2[23][18] , 
        \g2[23][17] , \g2[23][16] , \g2[23][15] , \g2[23][14] , \g2[23][13] , 
        \g2[23][12] , \g2[23][11] , \g2[23][10] , \g2[23][9] , \g2[23][8] , 
        \g2[23][7] , \g2[23][6] , \g2[23][5] , \g2[23][4] , \g2[23][3] , 
        \g2[23][2] , \g2[23][1] , 1'b0}), .sum({\g3[7][63] , \g3[7][62] , 
        \g3[7][61] , \g3[7][60] , \g3[7][59] , \g3[7][58] , \g3[7][57] , 
        \g3[7][56] , \g3[7][55] , \g3[7][54] , \g3[7][53] , \g3[7][52] , 
        \g3[7][51] , \g3[7][50] , \g3[7][49] , \g3[7][48] , \g3[7][47] , 
        \g3[7][46] , \g3[7][45] , \g3[7][44] , \g3[7][43] , \g3[7][42] , 
        \g3[7][41] , \g3[7][40] , \g3[7][39] , \g3[7][38] , \g3[7][37] , 
        \g3[7][36] , \g3[7][35] , \g3[7][34] , \g3[7][33] , \g3[7][32] , 
        \g3[7][31] , \g3[7][30] , \g3[7][29] , \g3[7][28] , \g3[7][27] , 
        \g3[7][26] , \g3[7][25] , \g3[7][24] , \g3[7][23] , \g3[7][22] , 
        \g3[7][21] , \g3[7][20] , \g3[7][19] , \g3[7][18] , \g3[7][17] , 
        \g3[7][16] , \g3[7][15] , \g3[7][14] , \g3[7][13] , \g3[7][12] , 
        \g3[7][11] , \g3[7][10] , \g3[7][9] , \g3[7][8] , \g3[7][7] , 
        \g3[7][6] , \g3[7][5] , \g3[7][4] , \g3[7][3] , \g3[7][2] , \g3[7][1] , 
        \g3[7][0] }), .cout({\g3[16][63] , \g3[16][62] , \g3[16][61] , 
        \g3[16][60] , \g3[16][59] , \g3[16][58] , \g3[16][57] , \g3[16][56] , 
        \g3[16][55] , \g3[16][54] , \g3[16][53] , \g3[16][52] , \g3[16][51] , 
        \g3[16][50] , \g3[16][49] , \g3[16][48] , \g3[16][47] , \g3[16][46] , 
        \g3[16][45] , \g3[16][44] , \g3[16][43] , \g3[16][42] , \g3[16][41] , 
        \g3[16][40] , \g3[16][39] , \g3[16][38] , \g3[16][37] , \g3[16][36] , 
        \g3[16][35] , \g3[16][34] , \g3[16][33] , \g3[16][32] , \g3[16][31] , 
        \g3[16][30] , \g3[16][29] , \g3[16][28] , \g3[16][27] , \g3[16][26] , 
        \g3[16][25] , \g3[16][24] , \g3[16][23] , \g3[16][22] , \g3[16][21] , 
        \g3[16][20] , \g3[16][19] , \g3[16][18] , \g3[16][17] , \g3[16][16] , 
        \g3[16][15] , \g3[16][14] , \g3[16][13] , \g3[16][12] , \g3[16][11] , 
        \g3[16][10] , \g3[16][9] , \g3[16][8] , \g3[16][7] , \g3[16][6] , 
        \g3[16][5] , \g3[16][4] , \g3[16][3] , \g3[16][2] , \g3[16][1] , 
        SYNOPSYS_UNCONNECTED__42}) );
  FullAdder_19 \level3[8].x0  ( .a({\g2[24][63] , \g2[24][62] , \g2[24][61] , 
        \g2[24][60] , \g2[24][59] , \g2[24][58] , \g2[24][57] , \g2[24][56] , 
        \g2[24][55] , \g2[24][54] , \g2[24][53] , \g2[24][52] , \g2[24][51] , 
        \g2[24][50] , \g2[24][49] , \g2[24][48] , \g2[24][47] , \g2[24][46] , 
        \g2[24][45] , \g2[24][44] , \g2[24][43] , \g2[24][42] , \g2[24][41] , 
        \g2[24][40] , \g2[24][39] , \g2[24][38] , \g2[24][37] , \g2[24][36] , 
        \g2[24][35] , \g2[24][34] , \g2[24][33] , \g2[24][32] , \g2[24][31] , 
        \g2[24][30] , \g2[24][29] , \g2[24][28] , \g2[24][27] , \g2[24][26] , 
        \g2[24][25] , \g2[24][24] , \g2[24][23] , \g2[24][22] , \g2[24][21] , 
        \g2[24][20] , \g2[24][19] , \g2[24][18] , \g2[24][17] , \g2[24][16] , 
        \g2[24][15] , \g2[24][14] , \g2[24][13] , \g2[24][12] , \g2[24][11] , 
        \g2[24][10] , \g2[24][9] , \g2[24][8] , \g2[24][7] , \g2[24][6] , 
        \g2[24][5] , \g2[24][4] , \g2[24][3] , \g2[24][2] , \g2[24][1] , 1'b0}), .b({\g2[25][63] , \g2[25][62] , \g2[25][61] , \g2[25][60] , \g2[25][59] , 
        \g2[25][58] , \g2[25][57] , \g2[25][56] , \g2[25][55] , \g2[25][54] , 
        \g2[25][53] , \g2[25][52] , \g2[25][51] , \g2[25][50] , \g2[25][49] , 
        \g2[25][48] , \g2[25][47] , \g2[25][46] , \g2[25][45] , \g2[25][44] , 
        \g2[25][43] , \g2[25][42] , \g2[25][41] , \g2[25][40] , \g2[25][39] , 
        \g2[25][38] , \g2[25][37] , \g2[25][36] , \g2[25][35] , \g2[25][34] , 
        \g2[25][33] , \g2[25][32] , \g2[25][31] , \g2[25][30] , \g2[25][29] , 
        \g2[25][28] , \g2[25][27] , \g2[25][26] , \g2[25][25] , \g2[25][24] , 
        \g2[25][23] , \g2[25][22] , \g2[25][21] , \g2[25][20] , \g2[25][19] , 
        \g2[25][18] , \g2[25][17] , \g2[25][16] , \g2[25][15] , \g2[25][14] , 
        \g2[25][13] , \g2[25][12] , \g2[25][11] , \g2[25][10] , \g2[25][9] , 
        \g2[25][8] , \g2[25][7] , \g2[25][6] , \g2[25][5] , \g2[25][4] , 
        \g2[25][3] , \g2[25][2] , \g2[25][1] , 1'b0}), .cin({\g2[26][63] , 
        \g2[26][62] , \g2[26][61] , \g2[26][60] , \g2[26][59] , \g2[26][58] , 
        \g2[26][57] , \g2[26][56] , \g2[26][55] , \g2[26][54] , \g2[26][53] , 
        \g2[26][52] , \g2[26][51] , \g2[26][50] , \g2[26][49] , \g2[26][48] , 
        \g2[26][47] , \g2[26][46] , \g2[26][45] , \g2[26][44] , \g2[26][43] , 
        \g2[26][42] , \g2[26][41] , \g2[26][40] , \g2[26][39] , \g2[26][38] , 
        \g2[26][37] , \g2[26][36] , \g2[26][35] , \g2[26][34] , \g2[26][33] , 
        \g2[26][32] , \g2[26][31] , \g2[26][30] , \g2[26][29] , \g2[26][28] , 
        \g2[26][27] , \g2[26][26] , \g2[26][25] , \g2[26][24] , \g2[26][23] , 
        \g2[26][22] , \g2[26][21] , \g2[26][20] , \g2[26][19] , \g2[26][18] , 
        \g2[26][17] , \g2[26][16] , \g2[26][15] , \g2[26][14] , \g2[26][13] , 
        \g2[26][12] , \g2[26][11] , \g2[26][10] , \g2[26][9] , \g2[26][8] , 
        \g2[26][7] , \g2[26][6] , \g2[26][5] , \g2[26][4] , \g2[26][3] , 
        \g2[26][2] , \g2[26][1] , 1'b0}), .sum({\g3[8][63] , \g3[8][62] , 
        \g3[8][61] , \g3[8][60] , \g3[8][59] , \g3[8][58] , \g3[8][57] , 
        \g3[8][56] , \g3[8][55] , \g3[8][54] , \g3[8][53] , \g3[8][52] , 
        \g3[8][51] , \g3[8][50] , \g3[8][49] , \g3[8][48] , \g3[8][47] , 
        \g3[8][46] , \g3[8][45] , \g3[8][44] , \g3[8][43] , \g3[8][42] , 
        \g3[8][41] , \g3[8][40] , \g3[8][39] , \g3[8][38] , \g3[8][37] , 
        \g3[8][36] , \g3[8][35] , \g3[8][34] , \g3[8][33] , \g3[8][32] , 
        \g3[8][31] , \g3[8][30] , \g3[8][29] , \g3[8][28] , \g3[8][27] , 
        \g3[8][26] , \g3[8][25] , \g3[8][24] , \g3[8][23] , \g3[8][22] , 
        \g3[8][21] , \g3[8][20] , \g3[8][19] , \g3[8][18] , \g3[8][17] , 
        \g3[8][16] , \g3[8][15] , \g3[8][14] , \g3[8][13] , \g3[8][12] , 
        \g3[8][11] , \g3[8][10] , \g3[8][9] , \g3[8][8] , \g3[8][7] , 
        \g3[8][6] , \g3[8][5] , \g3[8][4] , \g3[8][3] , \g3[8][2] , \g3[8][1] , 
        \g3[8][0] }), .cout({\g3[17][63] , \g3[17][62] , \g3[17][61] , 
        \g3[17][60] , \g3[17][59] , \g3[17][58] , \g3[17][57] , \g3[17][56] , 
        \g3[17][55] , \g3[17][54] , \g3[17][53] , \g3[17][52] , \g3[17][51] , 
        \g3[17][50] , \g3[17][49] , \g3[17][48] , \g3[17][47] , \g3[17][46] , 
        \g3[17][45] , \g3[17][44] , \g3[17][43] , \g3[17][42] , \g3[17][41] , 
        \g3[17][40] , \g3[17][39] , \g3[17][38] , \g3[17][37] , \g3[17][36] , 
        \g3[17][35] , \g3[17][34] , \g3[17][33] , \g3[17][32] , \g3[17][31] , 
        \g3[17][30] , \g3[17][29] , \g3[17][28] , \g3[17][27] , \g3[17][26] , 
        \g3[17][25] , \g3[17][24] , \g3[17][23] , \g3[17][22] , \g3[17][21] , 
        \g3[17][20] , \g3[17][19] , \g3[17][18] , \g3[17][17] , \g3[17][16] , 
        \g3[17][15] , \g3[17][14] , \g3[17][13] , \g3[17][12] , \g3[17][11] , 
        \g3[17][10] , \g3[17][9] , \g3[17][8] , \g3[17][7] , \g3[17][6] , 
        \g3[17][5] , \g3[17][4] , \g3[17][3] , \g3[17][2] , \g3[17][1] , 
        SYNOPSYS_UNCONNECTED__43}) );
  FullAdder_18 \level4[0].x1  ( .a({\g3[0][63] , \g3[0][62] , \g3[0][61] , 
        \g3[0][60] , \g3[0][59] , \g3[0][58] , \g3[0][57] , \g3[0][56] , 
        \g3[0][55] , \g3[0][54] , \g3[0][53] , \g3[0][52] , \g3[0][51] , 
        \g3[0][50] , \g3[0][49] , \g3[0][48] , \g3[0][47] , \g3[0][46] , 
        \g3[0][45] , \g3[0][44] , \g3[0][43] , \g3[0][42] , \g3[0][41] , 
        \g3[0][40] , \g3[0][39] , \g3[0][38] , \g3[0][37] , \g3[0][36] , 
        \g3[0][35] , \g3[0][34] , \g3[0][33] , \g3[0][32] , \g3[0][31] , 
        \g3[0][30] , \g3[0][29] , \g3[0][28] , \g3[0][27] , \g3[0][26] , 
        \g3[0][25] , \g3[0][24] , \g3[0][23] , \g3[0][22] , \g3[0][21] , 
        \g3[0][20] , \g3[0][19] , \g3[0][18] , \g3[0][17] , \g3[0][16] , 
        \g3[0][15] , \g3[0][14] , \g3[0][13] , \g3[0][12] , \g3[0][11] , 
        \g3[0][10] , \g3[0][9] , \g3[0][8] , \g3[0][7] , \g3[0][6] , 
        \g3[0][5] , \g3[0][4] , \g3[0][3] , \g3[0][2] , \g3[0][1] , \g3[0][0] }), .b({\g3[1][63] , \g3[1][62] , \g3[1][61] , \g3[1][60] , \g3[1][59] , 
        \g3[1][58] , \g3[1][57] , \g3[1][56] , \g3[1][55] , \g3[1][54] , 
        \g3[1][53] , \g3[1][52] , \g3[1][51] , \g3[1][50] , \g3[1][49] , 
        \g3[1][48] , \g3[1][47] , \g3[1][46] , \g3[1][45] , \g3[1][44] , 
        \g3[1][43] , \g3[1][42] , \g3[1][41] , \g3[1][40] , \g3[1][39] , 
        \g3[1][38] , \g3[1][37] , \g3[1][36] , \g3[1][35] , \g3[1][34] , 
        \g3[1][33] , \g3[1][32] , \g3[1][31] , \g3[1][30] , \g3[1][29] , 
        \g3[1][28] , \g3[1][27] , \g3[1][26] , \g3[1][25] , \g3[1][24] , 
        \g3[1][23] , \g3[1][22] , \g3[1][21] , \g3[1][20] , \g3[1][19] , 
        \g3[1][18] , \g3[1][17] , \g3[1][16] , \g3[1][15] , \g3[1][14] , 
        \g3[1][13] , \g3[1][12] , \g3[1][11] , \g3[1][10] , \g3[1][9] , 
        \g3[1][8] , \g3[1][7] , \g3[1][6] , \g3[1][5] , \g3[1][4] , \g3[1][3] , 
        \g3[1][2] , \g3[1][1] , \g3[1][0] }), .cin({\g3[2][63] , \g3[2][62] , 
        \g3[2][61] , \g3[2][60] , \g3[2][59] , \g3[2][58] , \g3[2][57] , 
        \g3[2][56] , \g3[2][55] , \g3[2][54] , \g3[2][53] , \g3[2][52] , 
        \g3[2][51] , \g3[2][50] , \g3[2][49] , \g3[2][48] , \g3[2][47] , 
        \g3[2][46] , \g3[2][45] , \g3[2][44] , \g3[2][43] , \g3[2][42] , 
        \g3[2][41] , \g3[2][40] , \g3[2][39] , \g3[2][38] , \g3[2][37] , 
        \g3[2][36] , \g3[2][35] , \g3[2][34] , \g3[2][33] , \g3[2][32] , 
        \g3[2][31] , \g3[2][30] , \g3[2][29] , \g3[2][28] , \g3[2][27] , 
        \g3[2][26] , \g3[2][25] , \g3[2][24] , \g3[2][23] , \g3[2][22] , 
        \g3[2][21] , \g3[2][20] , \g3[2][19] , \g3[2][18] , \g3[2][17] , 
        \g3[2][16] , \g3[2][15] , \g3[2][14] , \g3[2][13] , \g3[2][12] , 
        \g3[2][11] , \g3[2][10] , \g3[2][9] , \g3[2][8] , \g3[2][7] , 
        \g3[2][6] , \g3[2][5] , \g3[2][4] , \g3[2][3] , \g3[2][2] , \g3[2][1] , 
        \g3[2][0] }), .sum({\g4[0][63] , \g4[0][62] , \g4[0][61] , \g4[0][60] , 
        \g4[0][59] , \g4[0][58] , \g4[0][57] , \g4[0][56] , \g4[0][55] , 
        \g4[0][54] , \g4[0][53] , \g4[0][52] , \g4[0][51] , \g4[0][50] , 
        \g4[0][49] , \g4[0][48] , \g4[0][47] , \g4[0][46] , \g4[0][45] , 
        \g4[0][44] , \g4[0][43] , \g4[0][42] , \g4[0][41] , \g4[0][40] , 
        \g4[0][39] , \g4[0][38] , \g4[0][37] , \g4[0][36] , \g4[0][35] , 
        \g4[0][34] , \g4[0][33] , \g4[0][32] , \g4[0][31] , \g4[0][30] , 
        \g4[0][29] , \g4[0][28] , \g4[0][27] , \g4[0][26] , \g4[0][25] , 
        \g4[0][24] , \g4[0][23] , \g4[0][22] , \g4[0][21] , \g4[0][20] , 
        \g4[0][19] , \g4[0][18] , \g4[0][17] , \g4[0][16] , \g4[0][15] , 
        \g4[0][14] , \g4[0][13] , \g4[0][12] , \g4[0][11] , \g4[0][10] , 
        \g4[0][9] , \g4[0][8] , \g4[0][7] , \g4[0][6] , \g4[0][5] , \g4[0][4] , 
        \g4[0][3] , \g4[0][2] , \g4[0][1] , \g4[0][0] }), .cout({\g4[6][63] , 
        \g4[6][62] , \g4[6][61] , \g4[6][60] , \g4[6][59] , \g4[6][58] , 
        \g4[6][57] , \g4[6][56] , \g4[6][55] , \g4[6][54] , \g4[6][53] , 
        \g4[6][52] , \g4[6][51] , \g4[6][50] , \g4[6][49] , \g4[6][48] , 
        \g4[6][47] , \g4[6][46] , \g4[6][45] , \g4[6][44] , \g4[6][43] , 
        \g4[6][42] , \g4[6][41] , \g4[6][40] , \g4[6][39] , \g4[6][38] , 
        \g4[6][37] , \g4[6][36] , \g4[6][35] , \g4[6][34] , \g4[6][33] , 
        \g4[6][32] , \g4[6][31] , \g4[6][30] , \g4[6][29] , \g4[6][28] , 
        \g4[6][27] , \g4[6][26] , \g4[6][25] , \g4[6][24] , \g4[6][23] , 
        \g4[6][22] , \g4[6][21] , \g4[6][20] , \g4[6][19] , \g4[6][18] , 
        \g4[6][17] , \g4[6][16] , \g4[6][15] , \g4[6][14] , \g4[6][13] , 
        \g4[6][12] , \g4[6][11] , \g4[6][10] , \g4[6][9] , \g4[6][8] , 
        \g4[6][7] , \g4[6][6] , \g4[6][5] , \g4[6][4] , \g4[6][3] , \g4[6][2] , 
        \g4[6][1] , SYNOPSYS_UNCONNECTED__44}) );
  FullAdder_17 \level4[1].x1  ( .a({\g3[3][63] , \g3[3][62] , \g3[3][61] , 
        \g3[3][60] , \g3[3][59] , \g3[3][58] , \g3[3][57] , \g3[3][56] , 
        \g3[3][55] , \g3[3][54] , \g3[3][53] , \g3[3][52] , \g3[3][51] , 
        \g3[3][50] , \g3[3][49] , \g3[3][48] , \g3[3][47] , \g3[3][46] , 
        \g3[3][45] , \g3[3][44] , \g3[3][43] , \g3[3][42] , \g3[3][41] , 
        \g3[3][40] , \g3[3][39] , \g3[3][38] , \g3[3][37] , \g3[3][36] , 
        \g3[3][35] , \g3[3][34] , \g3[3][33] , \g3[3][32] , \g3[3][31] , 
        \g3[3][30] , \g3[3][29] , \g3[3][28] , \g3[3][27] , \g3[3][26] , 
        \g3[3][25] , \g3[3][24] , \g3[3][23] , \g3[3][22] , \g3[3][21] , 
        \g3[3][20] , \g3[3][19] , \g3[3][18] , \g3[3][17] , \g3[3][16] , 
        \g3[3][15] , \g3[3][14] , \g3[3][13] , \g3[3][12] , \g3[3][11] , 
        \g3[3][10] , \g3[3][9] , \g3[3][8] , \g3[3][7] , \g3[3][6] , 
        \g3[3][5] , \g3[3][4] , \g3[3][3] , \g3[3][2] , \g3[3][1] , \g3[3][0] }), .b({\g3[4][63] , \g3[4][62] , \g3[4][61] , \g3[4][60] , \g3[4][59] , 
        \g3[4][58] , \g3[4][57] , \g3[4][56] , \g3[4][55] , \g3[4][54] , 
        \g3[4][53] , \g3[4][52] , \g3[4][51] , \g3[4][50] , \g3[4][49] , 
        \g3[4][48] , \g3[4][47] , \g3[4][46] , \g3[4][45] , \g3[4][44] , 
        \g3[4][43] , \g3[4][42] , \g3[4][41] , \g3[4][40] , \g3[4][39] , 
        \g3[4][38] , \g3[4][37] , \g3[4][36] , \g3[4][35] , \g3[4][34] , 
        \g3[4][33] , \g3[4][32] , \g3[4][31] , \g3[4][30] , \g3[4][29] , 
        \g3[4][28] , \g3[4][27] , \g3[4][26] , \g3[4][25] , \g3[4][24] , 
        \g3[4][23] , \g3[4][22] , \g3[4][21] , \g3[4][20] , \g3[4][19] , 
        \g3[4][18] , \g3[4][17] , \g3[4][16] , \g3[4][15] , \g3[4][14] , 
        \g3[4][13] , \g3[4][12] , \g3[4][11] , \g3[4][10] , \g3[4][9] , 
        \g3[4][8] , \g3[4][7] , \g3[4][6] , \g3[4][5] , \g3[4][4] , \g3[4][3] , 
        \g3[4][2] , \g3[4][1] , \g3[4][0] }), .cin({\g3[5][63] , \g3[5][62] , 
        \g3[5][61] , \g3[5][60] , \g3[5][59] , \g3[5][58] , \g3[5][57] , 
        \g3[5][56] , \g3[5][55] , \g3[5][54] , \g3[5][53] , \g3[5][52] , 
        \g3[5][51] , \g3[5][50] , \g3[5][49] , \g3[5][48] , \g3[5][47] , 
        \g3[5][46] , \g3[5][45] , \g3[5][44] , \g3[5][43] , \g3[5][42] , 
        \g3[5][41] , \g3[5][40] , \g3[5][39] , \g3[5][38] , \g3[5][37] , 
        \g3[5][36] , \g3[5][35] , \g3[5][34] , \g3[5][33] , \g3[5][32] , 
        \g3[5][31] , \g3[5][30] , \g3[5][29] , \g3[5][28] , \g3[5][27] , 
        \g3[5][26] , \g3[5][25] , \g3[5][24] , \g3[5][23] , \g3[5][22] , 
        \g3[5][21] , \g3[5][20] , \g3[5][19] , \g3[5][18] , \g3[5][17] , 
        \g3[5][16] , \g3[5][15] , \g3[5][14] , \g3[5][13] , \g3[5][12] , 
        \g3[5][11] , \g3[5][10] , \g3[5][9] , \g3[5][8] , \g3[5][7] , 
        \g3[5][6] , \g3[5][5] , \g3[5][4] , \g3[5][3] , \g3[5][2] , \g3[5][1] , 
        \g3[5][0] }), .sum({\g4[1][63] , \g4[1][62] , \g4[1][61] , \g4[1][60] , 
        \g4[1][59] , \g4[1][58] , \g4[1][57] , \g4[1][56] , \g4[1][55] , 
        \g4[1][54] , \g4[1][53] , \g4[1][52] , \g4[1][51] , \g4[1][50] , 
        \g4[1][49] , \g4[1][48] , \g4[1][47] , \g4[1][46] , \g4[1][45] , 
        \g4[1][44] , \g4[1][43] , \g4[1][42] , \g4[1][41] , \g4[1][40] , 
        \g4[1][39] , \g4[1][38] , \g4[1][37] , \g4[1][36] , \g4[1][35] , 
        \g4[1][34] , \g4[1][33] , \g4[1][32] , \g4[1][31] , \g4[1][30] , 
        \g4[1][29] , \g4[1][28] , \g4[1][27] , \g4[1][26] , \g4[1][25] , 
        \g4[1][24] , \g4[1][23] , \g4[1][22] , \g4[1][21] , \g4[1][20] , 
        \g4[1][19] , \g4[1][18] , \g4[1][17] , \g4[1][16] , \g4[1][15] , 
        \g4[1][14] , \g4[1][13] , \g4[1][12] , \g4[1][11] , \g4[1][10] , 
        \g4[1][9] , \g4[1][8] , \g4[1][7] , \g4[1][6] , \g4[1][5] , \g4[1][4] , 
        \g4[1][3] , \g4[1][2] , \g4[1][1] , \g4[1][0] }), .cout({\g4[7][63] , 
        \g4[7][62] , \g4[7][61] , \g4[7][60] , \g4[7][59] , \g4[7][58] , 
        \g4[7][57] , \g4[7][56] , \g4[7][55] , \g4[7][54] , \g4[7][53] , 
        \g4[7][52] , \g4[7][51] , \g4[7][50] , \g4[7][49] , \g4[7][48] , 
        \g4[7][47] , \g4[7][46] , \g4[7][45] , \g4[7][44] , \g4[7][43] , 
        \g4[7][42] , \g4[7][41] , \g4[7][40] , \g4[7][39] , \g4[7][38] , 
        \g4[7][37] , \g4[7][36] , \g4[7][35] , \g4[7][34] , \g4[7][33] , 
        \g4[7][32] , \g4[7][31] , \g4[7][30] , \g4[7][29] , \g4[7][28] , 
        \g4[7][27] , \g4[7][26] , \g4[7][25] , \g4[7][24] , \g4[7][23] , 
        \g4[7][22] , \g4[7][21] , \g4[7][20] , \g4[7][19] , \g4[7][18] , 
        \g4[7][17] , \g4[7][16] , \g4[7][15] , \g4[7][14] , \g4[7][13] , 
        \g4[7][12] , \g4[7][11] , \g4[7][10] , \g4[7][9] , \g4[7][8] , 
        \g4[7][7] , \g4[7][6] , \g4[7][5] , \g4[7][4] , \g4[7][3] , \g4[7][2] , 
        \g4[7][1] , SYNOPSYS_UNCONNECTED__45}) );
  FullAdder_16 \level4[2].x1  ( .a({\g3[6][63] , \g3[6][62] , \g3[6][61] , 
        \g3[6][60] , \g3[6][59] , \g3[6][58] , \g3[6][57] , \g3[6][56] , 
        \g3[6][55] , \g3[6][54] , \g3[6][53] , \g3[6][52] , \g3[6][51] , 
        \g3[6][50] , \g3[6][49] , \g3[6][48] , \g3[6][47] , \g3[6][46] , 
        \g3[6][45] , \g3[6][44] , \g3[6][43] , \g3[6][42] , \g3[6][41] , 
        \g3[6][40] , \g3[6][39] , \g3[6][38] , \g3[6][37] , \g3[6][36] , 
        \g3[6][35] , \g3[6][34] , \g3[6][33] , \g3[6][32] , \g3[6][31] , 
        \g3[6][30] , \g3[6][29] , \g3[6][28] , \g3[6][27] , \g3[6][26] , 
        \g3[6][25] , \g3[6][24] , \g3[6][23] , \g3[6][22] , \g3[6][21] , 
        \g3[6][20] , \g3[6][19] , \g3[6][18] , \g3[6][17] , \g3[6][16] , 
        \g3[6][15] , \g3[6][14] , \g3[6][13] , \g3[6][12] , \g3[6][11] , 
        \g3[6][10] , \g3[6][9] , \g3[6][8] , \g3[6][7] , \g3[6][6] , 
        \g3[6][5] , \g3[6][4] , \g3[6][3] , \g3[6][2] , \g3[6][1] , \g3[6][0] }), .b({\g3[7][63] , \g3[7][62] , \g3[7][61] , \g3[7][60] , \g3[7][59] , 
        \g3[7][58] , \g3[7][57] , \g3[7][56] , \g3[7][55] , \g3[7][54] , 
        \g3[7][53] , \g3[7][52] , \g3[7][51] , \g3[7][50] , \g3[7][49] , 
        \g3[7][48] , \g3[7][47] , \g3[7][46] , \g3[7][45] , \g3[7][44] , 
        \g3[7][43] , \g3[7][42] , \g3[7][41] , \g3[7][40] , \g3[7][39] , 
        \g3[7][38] , \g3[7][37] , \g3[7][36] , \g3[7][35] , \g3[7][34] , 
        \g3[7][33] , \g3[7][32] , \g3[7][31] , \g3[7][30] , \g3[7][29] , 
        \g3[7][28] , \g3[7][27] , \g3[7][26] , \g3[7][25] , \g3[7][24] , 
        \g3[7][23] , \g3[7][22] , \g3[7][21] , \g3[7][20] , \g3[7][19] , 
        \g3[7][18] , \g3[7][17] , \g3[7][16] , \g3[7][15] , \g3[7][14] , 
        \g3[7][13] , \g3[7][12] , \g3[7][11] , \g3[7][10] , \g3[7][9] , 
        \g3[7][8] , \g3[7][7] , \g3[7][6] , \g3[7][5] , \g3[7][4] , \g3[7][3] , 
        \g3[7][2] , \g3[7][1] , \g3[7][0] }), .cin({\g3[8][63] , \g3[8][62] , 
        \g3[8][61] , \g3[8][60] , \g3[8][59] , \g3[8][58] , \g3[8][57] , 
        \g3[8][56] , \g3[8][55] , \g3[8][54] , \g3[8][53] , \g3[8][52] , 
        \g3[8][51] , \g3[8][50] , \g3[8][49] , \g3[8][48] , \g3[8][47] , 
        \g3[8][46] , \g3[8][45] , \g3[8][44] , \g3[8][43] , \g3[8][42] , 
        \g3[8][41] , \g3[8][40] , \g3[8][39] , \g3[8][38] , \g3[8][37] , 
        \g3[8][36] , \g3[8][35] , \g3[8][34] , \g3[8][33] , \g3[8][32] , 
        \g3[8][31] , \g3[8][30] , \g3[8][29] , \g3[8][28] , \g3[8][27] , 
        \g3[8][26] , \g3[8][25] , \g3[8][24] , \g3[8][23] , \g3[8][22] , 
        \g3[8][21] , \g3[8][20] , \g3[8][19] , \g3[8][18] , \g3[8][17] , 
        \g3[8][16] , \g3[8][15] , \g3[8][14] , \g3[8][13] , \g3[8][12] , 
        \g3[8][11] , \g3[8][10] , \g3[8][9] , \g3[8][8] , \g3[8][7] , 
        \g3[8][6] , \g3[8][5] , \g3[8][4] , \g3[8][3] , \g3[8][2] , \g3[8][1] , 
        \g3[8][0] }), .sum({\g4[2][63] , \g4[2][62] , \g4[2][61] , \g4[2][60] , 
        \g4[2][59] , \g4[2][58] , \g4[2][57] , \g4[2][56] , \g4[2][55] , 
        \g4[2][54] , \g4[2][53] , \g4[2][52] , \g4[2][51] , \g4[2][50] , 
        \g4[2][49] , \g4[2][48] , \g4[2][47] , \g4[2][46] , \g4[2][45] , 
        \g4[2][44] , \g4[2][43] , \g4[2][42] , \g4[2][41] , \g4[2][40] , 
        \g4[2][39] , \g4[2][38] , \g4[2][37] , \g4[2][36] , \g4[2][35] , 
        \g4[2][34] , \g4[2][33] , \g4[2][32] , \g4[2][31] , \g4[2][30] , 
        \g4[2][29] , \g4[2][28] , \g4[2][27] , \g4[2][26] , \g4[2][25] , 
        \g4[2][24] , \g4[2][23] , \g4[2][22] , \g4[2][21] , \g4[2][20] , 
        \g4[2][19] , \g4[2][18] , \g4[2][17] , \g4[2][16] , \g4[2][15] , 
        \g4[2][14] , \g4[2][13] , \g4[2][12] , \g4[2][11] , \g4[2][10] , 
        \g4[2][9] , \g4[2][8] , \g4[2][7] , \g4[2][6] , \g4[2][5] , \g4[2][4] , 
        \g4[2][3] , \g4[2][2] , \g4[2][1] , \g4[2][0] }), .cout({\g4[8][63] , 
        \g4[8][62] , \g4[8][61] , \g4[8][60] , \g4[8][59] , \g4[8][58] , 
        \g4[8][57] , \g4[8][56] , \g4[8][55] , \g4[8][54] , \g4[8][53] , 
        \g4[8][52] , \g4[8][51] , \g4[8][50] , \g4[8][49] , \g4[8][48] , 
        \g4[8][47] , \g4[8][46] , \g4[8][45] , \g4[8][44] , \g4[8][43] , 
        \g4[8][42] , \g4[8][41] , \g4[8][40] , \g4[8][39] , \g4[8][38] , 
        \g4[8][37] , \g4[8][36] , \g4[8][35] , \g4[8][34] , \g4[8][33] , 
        \g4[8][32] , \g4[8][31] , \g4[8][30] , \g4[8][29] , \g4[8][28] , 
        \g4[8][27] , \g4[8][26] , \g4[8][25] , \g4[8][24] , \g4[8][23] , 
        \g4[8][22] , \g4[8][21] , \g4[8][20] , \g4[8][19] , \g4[8][18] , 
        \g4[8][17] , \g4[8][16] , \g4[8][15] , \g4[8][14] , \g4[8][13] , 
        \g4[8][12] , \g4[8][11] , \g4[8][10] , \g4[8][9] , \g4[8][8] , 
        \g4[8][7] , \g4[8][6] , \g4[8][5] , \g4[8][4] , \g4[8][3] , \g4[8][2] , 
        \g4[8][1] , SYNOPSYS_UNCONNECTED__46}) );
  FullAdder_15 \level4[3].x1  ( .a({\g3[9][63] , \g3[9][62] , \g3[9][61] , 
        \g3[9][60] , \g3[9][59] , \g3[9][58] , \g3[9][57] , \g3[9][56] , 
        \g3[9][55] , \g3[9][54] , \g3[9][53] , \g3[9][52] , \g3[9][51] , 
        \g3[9][50] , \g3[9][49] , \g3[9][48] , \g3[9][47] , \g3[9][46] , 
        \g3[9][45] , \g3[9][44] , \g3[9][43] , \g3[9][42] , \g3[9][41] , 
        \g3[9][40] , \g3[9][39] , \g3[9][38] , \g3[9][37] , \g3[9][36] , 
        \g3[9][35] , \g3[9][34] , \g3[9][33] , \g3[9][32] , \g3[9][31] , 
        \g3[9][30] , \g3[9][29] , \g3[9][28] , \g3[9][27] , \g3[9][26] , 
        \g3[9][25] , \g3[9][24] , \g3[9][23] , \g3[9][22] , \g3[9][21] , 
        \g3[9][20] , \g3[9][19] , \g3[9][18] , \g3[9][17] , \g3[9][16] , 
        \g3[9][15] , \g3[9][14] , \g3[9][13] , \g3[9][12] , \g3[9][11] , 
        \g3[9][10] , \g3[9][9] , \g3[9][8] , \g3[9][7] , \g3[9][6] , 
        \g3[9][5] , \g3[9][4] , \g3[9][3] , \g3[9][2] , \g3[9][1] , 1'b0}), 
        .b({\g3[10][63] , \g3[10][62] , \g3[10][61] , \g3[10][60] , 
        \g3[10][59] , \g3[10][58] , \g3[10][57] , \g3[10][56] , \g3[10][55] , 
        \g3[10][54] , \g3[10][53] , \g3[10][52] , \g3[10][51] , \g3[10][50] , 
        \g3[10][49] , \g3[10][48] , \g3[10][47] , \g3[10][46] , \g3[10][45] , 
        \g3[10][44] , \g3[10][43] , \g3[10][42] , \g3[10][41] , \g3[10][40] , 
        \g3[10][39] , \g3[10][38] , \g3[10][37] , \g3[10][36] , \g3[10][35] , 
        \g3[10][34] , \g3[10][33] , \g3[10][32] , \g3[10][31] , \g3[10][30] , 
        \g3[10][29] , \g3[10][28] , \g3[10][27] , \g3[10][26] , \g3[10][25] , 
        \g3[10][24] , \g3[10][23] , \g3[10][22] , \g3[10][21] , \g3[10][20] , 
        \g3[10][19] , \g3[10][18] , \g3[10][17] , \g3[10][16] , \g3[10][15] , 
        \g3[10][14] , \g3[10][13] , \g3[10][12] , \g3[10][11] , \g3[10][10] , 
        \g3[10][9] , \g3[10][8] , \g3[10][7] , \g3[10][6] , \g3[10][5] , 
        \g3[10][4] , \g3[10][3] , \g3[10][2] , \g3[10][1] , 1'b0}), .cin({
        \g3[11][63] , \g3[11][62] , \g3[11][61] , \g3[11][60] , \g3[11][59] , 
        \g3[11][58] , \g3[11][57] , \g3[11][56] , \g3[11][55] , \g3[11][54] , 
        \g3[11][53] , \g3[11][52] , \g3[11][51] , \g3[11][50] , \g3[11][49] , 
        \g3[11][48] , \g3[11][47] , \g3[11][46] , \g3[11][45] , \g3[11][44] , 
        \g3[11][43] , \g3[11][42] , \g3[11][41] , \g3[11][40] , \g3[11][39] , 
        \g3[11][38] , \g3[11][37] , \g3[11][36] , \g3[11][35] , \g3[11][34] , 
        \g3[11][33] , \g3[11][32] , \g3[11][31] , \g3[11][30] , \g3[11][29] , 
        \g3[11][28] , \g3[11][27] , \g3[11][26] , \g3[11][25] , \g3[11][24] , 
        \g3[11][23] , \g3[11][22] , \g3[11][21] , \g3[11][20] , \g3[11][19] , 
        \g3[11][18] , \g3[11][17] , \g3[11][16] , \g3[11][15] , \g3[11][14] , 
        \g3[11][13] , \g3[11][12] , \g3[11][11] , \g3[11][10] , \g3[11][9] , 
        \g3[11][8] , \g3[11][7] , \g3[11][6] , \g3[11][5] , \g3[11][4] , 
        \g3[11][3] , \g3[11][2] , \g3[11][1] , 1'b0}), .sum({\g4[3][63] , 
        \g4[3][62] , \g4[3][61] , \g4[3][60] , \g4[3][59] , \g4[3][58] , 
        \g4[3][57] , \g4[3][56] , \g4[3][55] , \g4[3][54] , \g4[3][53] , 
        \g4[3][52] , \g4[3][51] , \g4[3][50] , \g4[3][49] , \g4[3][48] , 
        \g4[3][47] , \g4[3][46] , \g4[3][45] , \g4[3][44] , \g4[3][43] , 
        \g4[3][42] , \g4[3][41] , \g4[3][40] , \g4[3][39] , \g4[3][38] , 
        \g4[3][37] , \g4[3][36] , \g4[3][35] , \g4[3][34] , \g4[3][33] , 
        \g4[3][32] , \g4[3][31] , \g4[3][30] , \g4[3][29] , \g4[3][28] , 
        \g4[3][27] , \g4[3][26] , \g4[3][25] , \g4[3][24] , \g4[3][23] , 
        \g4[3][22] , \g4[3][21] , \g4[3][20] , \g4[3][19] , \g4[3][18] , 
        \g4[3][17] , \g4[3][16] , \g4[3][15] , \g4[3][14] , \g4[3][13] , 
        \g4[3][12] , \g4[3][11] , \g4[3][10] , \g4[3][9] , \g4[3][8] , 
        \g4[3][7] , \g4[3][6] , \g4[3][5] , \g4[3][4] , \g4[3][3] , \g4[3][2] , 
        \g4[3][1] , \g4[3][0] }), .cout({\g4[9][63] , \g4[9][62] , \g4[9][61] , 
        \g4[9][60] , \g4[9][59] , \g4[9][58] , \g4[9][57] , \g4[9][56] , 
        \g4[9][55] , \g4[9][54] , \g4[9][53] , \g4[9][52] , \g4[9][51] , 
        \g4[9][50] , \g4[9][49] , \g4[9][48] , \g4[9][47] , \g4[9][46] , 
        \g4[9][45] , \g4[9][44] , \g4[9][43] , \g4[9][42] , \g4[9][41] , 
        \g4[9][40] , \g4[9][39] , \g4[9][38] , \g4[9][37] , \g4[9][36] , 
        \g4[9][35] , \g4[9][34] , \g4[9][33] , \g4[9][32] , \g4[9][31] , 
        \g4[9][30] , \g4[9][29] , \g4[9][28] , \g4[9][27] , \g4[9][26] , 
        \g4[9][25] , \g4[9][24] , \g4[9][23] , \g4[9][22] , \g4[9][21] , 
        \g4[9][20] , \g4[9][19] , \g4[9][18] , \g4[9][17] , \g4[9][16] , 
        \g4[9][15] , \g4[9][14] , \g4[9][13] , \g4[9][12] , \g4[9][11] , 
        \g4[9][10] , \g4[9][9] , \g4[9][8] , \g4[9][7] , \g4[9][6] , 
        \g4[9][5] , \g4[9][4] , \g4[9][3] , \g4[9][2] , \g4[9][1] , 
        SYNOPSYS_UNCONNECTED__47}) );
  FullAdder_14 \level4[4].x1  ( .a({\g3[12][63] , \g3[12][62] , \g3[12][61] , 
        \g3[12][60] , \g3[12][59] , \g3[12][58] , \g3[12][57] , \g3[12][56] , 
        \g3[12][55] , \g3[12][54] , \g3[12][53] , \g3[12][52] , \g3[12][51] , 
        \g3[12][50] , \g3[12][49] , \g3[12][48] , \g3[12][47] , \g3[12][46] , 
        \g3[12][45] , \g3[12][44] , \g3[12][43] , \g3[12][42] , \g3[12][41] , 
        \g3[12][40] , \g3[12][39] , \g3[12][38] , \g3[12][37] , \g3[12][36] , 
        \g3[12][35] , \g3[12][34] , \g3[12][33] , \g3[12][32] , \g3[12][31] , 
        \g3[12][30] , \g3[12][29] , \g3[12][28] , \g3[12][27] , \g3[12][26] , 
        \g3[12][25] , \g3[12][24] , \g3[12][23] , \g3[12][22] , \g3[12][21] , 
        \g3[12][20] , \g3[12][19] , \g3[12][18] , \g3[12][17] , \g3[12][16] , 
        \g3[12][15] , \g3[12][14] , \g3[12][13] , \g3[12][12] , \g3[12][11] , 
        \g3[12][10] , \g3[12][9] , \g3[12][8] , \g3[12][7] , \g3[12][6] , 
        \g3[12][5] , \g3[12][4] , \g3[12][3] , \g3[12][2] , \g3[12][1] , 1'b0}), .b({\g3[13][63] , \g3[13][62] , \g3[13][61] , \g3[13][60] , \g3[13][59] , 
        \g3[13][58] , \g3[13][57] , \g3[13][56] , \g3[13][55] , \g3[13][54] , 
        \g3[13][53] , \g3[13][52] , \g3[13][51] , \g3[13][50] , \g3[13][49] , 
        \g3[13][48] , \g3[13][47] , \g3[13][46] , \g3[13][45] , \g3[13][44] , 
        \g3[13][43] , \g3[13][42] , \g3[13][41] , \g3[13][40] , \g3[13][39] , 
        \g3[13][38] , \g3[13][37] , \g3[13][36] , \g3[13][35] , \g3[13][34] , 
        \g3[13][33] , \g3[13][32] , \g3[13][31] , \g3[13][30] , \g3[13][29] , 
        \g3[13][28] , \g3[13][27] , \g3[13][26] , \g3[13][25] , \g3[13][24] , 
        \g3[13][23] , \g3[13][22] , \g3[13][21] , \g3[13][20] , \g3[13][19] , 
        \g3[13][18] , \g3[13][17] , \g3[13][16] , \g3[13][15] , \g3[13][14] , 
        \g3[13][13] , \g3[13][12] , \g3[13][11] , \g3[13][10] , \g3[13][9] , 
        \g3[13][8] , \g3[13][7] , \g3[13][6] , \g3[13][5] , \g3[13][4] , 
        \g3[13][3] , \g3[13][2] , \g3[13][1] , 1'b0}), .cin({\g3[14][63] , 
        \g3[14][62] , \g3[14][61] , \g3[14][60] , \g3[14][59] , \g3[14][58] , 
        \g3[14][57] , \g3[14][56] , \g3[14][55] , \g3[14][54] , \g3[14][53] , 
        \g3[14][52] , \g3[14][51] , \g3[14][50] , \g3[14][49] , \g3[14][48] , 
        \g3[14][47] , \g3[14][46] , \g3[14][45] , \g3[14][44] , \g3[14][43] , 
        \g3[14][42] , \g3[14][41] , \g3[14][40] , \g3[14][39] , \g3[14][38] , 
        \g3[14][37] , \g3[14][36] , \g3[14][35] , \g3[14][34] , \g3[14][33] , 
        \g3[14][32] , \g3[14][31] , \g3[14][30] , \g3[14][29] , \g3[14][28] , 
        \g3[14][27] , \g3[14][26] , \g3[14][25] , \g3[14][24] , \g3[14][23] , 
        \g3[14][22] , \g3[14][21] , \g3[14][20] , \g3[14][19] , \g3[14][18] , 
        \g3[14][17] , \g3[14][16] , \g3[14][15] , \g3[14][14] , \g3[14][13] , 
        \g3[14][12] , \g3[14][11] , \g3[14][10] , \g3[14][9] , \g3[14][8] , 
        \g3[14][7] , \g3[14][6] , \g3[14][5] , \g3[14][4] , \g3[14][3] , 
        \g3[14][2] , \g3[14][1] , 1'b0}), .sum({\g4[4][63] , \g4[4][62] , 
        \g4[4][61] , \g4[4][60] , \g4[4][59] , \g4[4][58] , \g4[4][57] , 
        \g4[4][56] , \g4[4][55] , \g4[4][54] , \g4[4][53] , \g4[4][52] , 
        \g4[4][51] , \g4[4][50] , \g4[4][49] , \g4[4][48] , \g4[4][47] , 
        \g4[4][46] , \g4[4][45] , \g4[4][44] , \g4[4][43] , \g4[4][42] , 
        \g4[4][41] , \g4[4][40] , \g4[4][39] , \g4[4][38] , \g4[4][37] , 
        \g4[4][36] , \g4[4][35] , \g4[4][34] , \g4[4][33] , \g4[4][32] , 
        \g4[4][31] , \g4[4][30] , \g4[4][29] , \g4[4][28] , \g4[4][27] , 
        \g4[4][26] , \g4[4][25] , \g4[4][24] , \g4[4][23] , \g4[4][22] , 
        \g4[4][21] , \g4[4][20] , \g4[4][19] , \g4[4][18] , \g4[4][17] , 
        \g4[4][16] , \g4[4][15] , \g4[4][14] , \g4[4][13] , \g4[4][12] , 
        \g4[4][11] , \g4[4][10] , \g4[4][9] , \g4[4][8] , \g4[4][7] , 
        \g4[4][6] , \g4[4][5] , \g4[4][4] , \g4[4][3] , \g4[4][2] , \g4[4][1] , 
        \g4[4][0] }), .cout({\g4[10][63] , \g4[10][62] , \g4[10][61] , 
        \g4[10][60] , \g4[10][59] , \g4[10][58] , \g4[10][57] , \g4[10][56] , 
        \g4[10][55] , \g4[10][54] , \g4[10][53] , \g4[10][52] , \g4[10][51] , 
        \g4[10][50] , \g4[10][49] , \g4[10][48] , \g4[10][47] , \g4[10][46] , 
        \g4[10][45] , \g4[10][44] , \g4[10][43] , \g4[10][42] , \g4[10][41] , 
        \g4[10][40] , \g4[10][39] , \g4[10][38] , \g4[10][37] , \g4[10][36] , 
        \g4[10][35] , \g4[10][34] , \g4[10][33] , \g4[10][32] , \g4[10][31] , 
        \g4[10][30] , \g4[10][29] , \g4[10][28] , \g4[10][27] , \g4[10][26] , 
        \g4[10][25] , \g4[10][24] , \g4[10][23] , \g4[10][22] , \g4[10][21] , 
        \g4[10][20] , \g4[10][19] , \g4[10][18] , \g4[10][17] , \g4[10][16] , 
        \g4[10][15] , \g4[10][14] , \g4[10][13] , \g4[10][12] , \g4[10][11] , 
        \g4[10][10] , \g4[10][9] , \g4[10][8] , \g4[10][7] , \g4[10][6] , 
        \g4[10][5] , \g4[10][4] , \g4[10][3] , \g4[10][2] , \g4[10][1] , 
        SYNOPSYS_UNCONNECTED__48}) );
  FullAdder_13 \level4[5].x1  ( .a({\g3[15][63] , \g3[15][62] , \g3[15][61] , 
        \g3[15][60] , \g3[15][59] , \g3[15][58] , \g3[15][57] , \g3[15][56] , 
        \g3[15][55] , \g3[15][54] , \g3[15][53] , \g3[15][52] , \g3[15][51] , 
        \g3[15][50] , \g3[15][49] , \g3[15][48] , \g3[15][47] , \g3[15][46] , 
        \g3[15][45] , \g3[15][44] , \g3[15][43] , \g3[15][42] , \g3[15][41] , 
        \g3[15][40] , \g3[15][39] , \g3[15][38] , \g3[15][37] , \g3[15][36] , 
        \g3[15][35] , \g3[15][34] , \g3[15][33] , \g3[15][32] , \g3[15][31] , 
        \g3[15][30] , \g3[15][29] , \g3[15][28] , \g3[15][27] , \g3[15][26] , 
        \g3[15][25] , \g3[15][24] , \g3[15][23] , \g3[15][22] , \g3[15][21] , 
        \g3[15][20] , \g3[15][19] , \g3[15][18] , \g3[15][17] , \g3[15][16] , 
        \g3[15][15] , \g3[15][14] , \g3[15][13] , \g3[15][12] , \g3[15][11] , 
        \g3[15][10] , \g3[15][9] , \g3[15][8] , \g3[15][7] , \g3[15][6] , 
        \g3[15][5] , \g3[15][4] , \g3[15][3] , \g3[15][2] , \g3[15][1] , 1'b0}), .b({\g3[16][63] , \g3[16][62] , \g3[16][61] , \g3[16][60] , \g3[16][59] , 
        \g3[16][58] , \g3[16][57] , \g3[16][56] , \g3[16][55] , \g3[16][54] , 
        \g3[16][53] , \g3[16][52] , \g3[16][51] , \g3[16][50] , \g3[16][49] , 
        \g3[16][48] , \g3[16][47] , \g3[16][46] , \g3[16][45] , \g3[16][44] , 
        \g3[16][43] , \g3[16][42] , \g3[16][41] , \g3[16][40] , \g3[16][39] , 
        \g3[16][38] , \g3[16][37] , \g3[16][36] , \g3[16][35] , \g3[16][34] , 
        \g3[16][33] , \g3[16][32] , \g3[16][31] , \g3[16][30] , \g3[16][29] , 
        \g3[16][28] , \g3[16][27] , \g3[16][26] , \g3[16][25] , \g3[16][24] , 
        \g3[16][23] , \g3[16][22] , \g3[16][21] , \g3[16][20] , \g3[16][19] , 
        \g3[16][18] , \g3[16][17] , \g3[16][16] , \g3[16][15] , \g3[16][14] , 
        \g3[16][13] , \g3[16][12] , \g3[16][11] , \g3[16][10] , \g3[16][9] , 
        \g3[16][8] , \g3[16][7] , \g3[16][6] , \g3[16][5] , \g3[16][4] , 
        \g3[16][3] , \g3[16][2] , \g3[16][1] , 1'b0}), .cin({\g3[17][63] , 
        \g3[17][62] , \g3[17][61] , \g3[17][60] , \g3[17][59] , \g3[17][58] , 
        \g3[17][57] , \g3[17][56] , \g3[17][55] , \g3[17][54] , \g3[17][53] , 
        \g3[17][52] , \g3[17][51] , \g3[17][50] , \g3[17][49] , \g3[17][48] , 
        \g3[17][47] , \g3[17][46] , \g3[17][45] , \g3[17][44] , \g3[17][43] , 
        \g3[17][42] , \g3[17][41] , \g3[17][40] , \g3[17][39] , \g3[17][38] , 
        \g3[17][37] , \g3[17][36] , \g3[17][35] , \g3[17][34] , \g3[17][33] , 
        \g3[17][32] , \g3[17][31] , \g3[17][30] , \g3[17][29] , \g3[17][28] , 
        \g3[17][27] , \g3[17][26] , \g3[17][25] , \g3[17][24] , \g3[17][23] , 
        \g3[17][22] , \g3[17][21] , \g3[17][20] , \g3[17][19] , \g3[17][18] , 
        \g3[17][17] , \g3[17][16] , \g3[17][15] , \g3[17][14] , \g3[17][13] , 
        \g3[17][12] , \g3[17][11] , \g3[17][10] , \g3[17][9] , \g3[17][8] , 
        \g3[17][7] , \g3[17][6] , \g3[17][5] , \g3[17][4] , \g3[17][3] , 
        \g3[17][2] , \g3[17][1] , 1'b0}), .sum({\g4[5][63] , \g4[5][62] , 
        \g4[5][61] , \g4[5][60] , \g4[5][59] , \g4[5][58] , \g4[5][57] , 
        \g4[5][56] , \g4[5][55] , \g4[5][54] , \g4[5][53] , \g4[5][52] , 
        \g4[5][51] , \g4[5][50] , \g4[5][49] , \g4[5][48] , \g4[5][47] , 
        \g4[5][46] , \g4[5][45] , \g4[5][44] , \g4[5][43] , \g4[5][42] , 
        \g4[5][41] , \g4[5][40] , \g4[5][39] , \g4[5][38] , \g4[5][37] , 
        \g4[5][36] , \g4[5][35] , \g4[5][34] , \g4[5][33] , \g4[5][32] , 
        \g4[5][31] , \g4[5][30] , \g4[5][29] , \g4[5][28] , \g4[5][27] , 
        \g4[5][26] , \g4[5][25] , \g4[5][24] , \g4[5][23] , \g4[5][22] , 
        \g4[5][21] , \g4[5][20] , \g4[5][19] , \g4[5][18] , \g4[5][17] , 
        \g4[5][16] , \g4[5][15] , \g4[5][14] , \g4[5][13] , \g4[5][12] , 
        \g4[5][11] , \g4[5][10] , \g4[5][9] , \g4[5][8] , \g4[5][7] , 
        \g4[5][6] , \g4[5][5] , \g4[5][4] , \g4[5][3] , \g4[5][2] , \g4[5][1] , 
        \g4[5][0] }), .cout({\g4[11][63] , \g4[11][62] , \g4[11][61] , 
        \g4[11][60] , \g4[11][59] , \g4[11][58] , \g4[11][57] , \g4[11][56] , 
        \g4[11][55] , \g4[11][54] , \g4[11][53] , \g4[11][52] , \g4[11][51] , 
        \g4[11][50] , \g4[11][49] , \g4[11][48] , \g4[11][47] , \g4[11][46] , 
        \g4[11][45] , \g4[11][44] , \g4[11][43] , \g4[11][42] , \g4[11][41] , 
        \g4[11][40] , \g4[11][39] , \g4[11][38] , \g4[11][37] , \g4[11][36] , 
        \g4[11][35] , \g4[11][34] , \g4[11][33] , \g4[11][32] , \g4[11][31] , 
        \g4[11][30] , \g4[11][29] , \g4[11][28] , \g4[11][27] , \g4[11][26] , 
        \g4[11][25] , \g4[11][24] , \g4[11][23] , \g4[11][22] , \g4[11][21] , 
        \g4[11][20] , \g4[11][19] , \g4[11][18] , \g4[11][17] , \g4[11][16] , 
        \g4[11][15] , \g4[11][14] , \g4[11][13] , \g4[11][12] , \g4[11][11] , 
        \g4[11][10] , \g4[11][9] , \g4[11][8] , \g4[11][7] , \g4[11][6] , 
        \g4[11][5] , \g4[11][4] , \g4[11][3] , \g4[11][2] , \g4[11][1] , 
        SYNOPSYS_UNCONNECTED__49}) );
  FullAdder_12 \level5[0].x2  ( .a({\g4[0][63] , \g4[0][62] , \g4[0][61] , 
        \g4[0][60] , \g4[0][59] , \g4[0][58] , \g4[0][57] , \g4[0][56] , 
        \g4[0][55] , \g4[0][54] , \g4[0][53] , \g4[0][52] , \g4[0][51] , 
        \g4[0][50] , \g4[0][49] , \g4[0][48] , \g4[0][47] , \g4[0][46] , 
        \g4[0][45] , \g4[0][44] , \g4[0][43] , \g4[0][42] , \g4[0][41] , 
        \g4[0][40] , \g4[0][39] , \g4[0][38] , \g4[0][37] , \g4[0][36] , 
        \g4[0][35] , \g4[0][34] , \g4[0][33] , \g4[0][32] , \g4[0][31] , 
        \g4[0][30] , \g4[0][29] , \g4[0][28] , \g4[0][27] , \g4[0][26] , 
        \g4[0][25] , \g4[0][24] , \g4[0][23] , \g4[0][22] , \g4[0][21] , 
        \g4[0][20] , \g4[0][19] , \g4[0][18] , \g4[0][17] , \g4[0][16] , 
        \g4[0][15] , \g4[0][14] , \g4[0][13] , \g4[0][12] , \g4[0][11] , 
        \g4[0][10] , \g4[0][9] , \g4[0][8] , \g4[0][7] , \g4[0][6] , 
        \g4[0][5] , \g4[0][4] , \g4[0][3] , \g4[0][2] , \g4[0][1] , \g4[0][0] }), .b({\g4[1][63] , \g4[1][62] , \g4[1][61] , \g4[1][60] , \g4[1][59] , 
        \g4[1][58] , \g4[1][57] , \g4[1][56] , \g4[1][55] , \g4[1][54] , 
        \g4[1][53] , \g4[1][52] , \g4[1][51] , \g4[1][50] , \g4[1][49] , 
        \g4[1][48] , \g4[1][47] , \g4[1][46] , \g4[1][45] , \g4[1][44] , 
        \g4[1][43] , \g4[1][42] , \g4[1][41] , \g4[1][40] , \g4[1][39] , 
        \g4[1][38] , \g4[1][37] , \g4[1][36] , \g4[1][35] , \g4[1][34] , 
        \g4[1][33] , \g4[1][32] , \g4[1][31] , \g4[1][30] , \g4[1][29] , 
        \g4[1][28] , \g4[1][27] , \g4[1][26] , \g4[1][25] , \g4[1][24] , 
        \g4[1][23] , \g4[1][22] , \g4[1][21] , \g4[1][20] , \g4[1][19] , 
        \g4[1][18] , \g4[1][17] , \g4[1][16] , \g4[1][15] , \g4[1][14] , 
        \g4[1][13] , \g4[1][12] , \g4[1][11] , \g4[1][10] , \g4[1][9] , 
        \g4[1][8] , \g4[1][7] , \g4[1][6] , \g4[1][5] , \g4[1][4] , \g4[1][3] , 
        \g4[1][2] , \g4[1][1] , \g4[1][0] }), .cin({\g4[2][63] , \g4[2][62] , 
        \g4[2][61] , \g4[2][60] , \g4[2][59] , \g4[2][58] , \g4[2][57] , 
        \g4[2][56] , \g4[2][55] , \g4[2][54] , \g4[2][53] , \g4[2][52] , 
        \g4[2][51] , \g4[2][50] , \g4[2][49] , \g4[2][48] , \g4[2][47] , 
        \g4[2][46] , \g4[2][45] , \g4[2][44] , \g4[2][43] , \g4[2][42] , 
        \g4[2][41] , \g4[2][40] , \g4[2][39] , \g4[2][38] , \g4[2][37] , 
        \g4[2][36] , \g4[2][35] , \g4[2][34] , \g4[2][33] , \g4[2][32] , 
        \g4[2][31] , \g4[2][30] , \g4[2][29] , \g4[2][28] , \g4[2][27] , 
        \g4[2][26] , \g4[2][25] , \g4[2][24] , \g4[2][23] , \g4[2][22] , 
        \g4[2][21] , \g4[2][20] , \g4[2][19] , \g4[2][18] , \g4[2][17] , 
        \g4[2][16] , \g4[2][15] , \g4[2][14] , \g4[2][13] , \g4[2][12] , 
        \g4[2][11] , \g4[2][10] , \g4[2][9] , \g4[2][8] , \g4[2][7] , 
        \g4[2][6] , \g4[2][5] , \g4[2][4] , \g4[2][3] , \g4[2][2] , \g4[2][1] , 
        \g4[2][0] }), .sum({\g5[0][63] , \g5[0][62] , \g5[0][61] , \g5[0][60] , 
        \g5[0][59] , \g5[0][58] , \g5[0][57] , \g5[0][56] , \g5[0][55] , 
        \g5[0][54] , \g5[0][53] , \g5[0][52] , \g5[0][51] , \g5[0][50] , 
        \g5[0][49] , \g5[0][48] , \g5[0][47] , \g5[0][46] , \g5[0][45] , 
        \g5[0][44] , \g5[0][43] , \g5[0][42] , \g5[0][41] , \g5[0][40] , 
        \g5[0][39] , \g5[0][38] , \g5[0][37] , \g5[0][36] , \g5[0][35] , 
        \g5[0][34] , \g5[0][33] , \g5[0][32] , \g5[0][31] , \g5[0][30] , 
        \g5[0][29] , \g5[0][28] , \g5[0][27] , \g5[0][26] , \g5[0][25] , 
        \g5[0][24] , \g5[0][23] , \g5[0][22] , \g5[0][21] , \g5[0][20] , 
        \g5[0][19] , \g5[0][18] , \g5[0][17] , \g5[0][16] , \g5[0][15] , 
        \g5[0][14] , \g5[0][13] , \g5[0][12] , \g5[0][11] , \g5[0][10] , 
        \g5[0][9] , \g5[0][8] , \g5[0][7] , \g5[0][6] , \g5[0][5] , \g5[0][4] , 
        \g5[0][3] , \g5[0][2] , \g5[0][1] , \g5[0][0] }), .cout({\g5[4][63] , 
        \g5[4][62] , \g5[4][61] , \g5[4][60] , \g5[4][59] , \g5[4][58] , 
        \g5[4][57] , \g5[4][56] , \g5[4][55] , \g5[4][54] , \g5[4][53] , 
        \g5[4][52] , \g5[4][51] , \g5[4][50] , \g5[4][49] , \g5[4][48] , 
        \g5[4][47] , \g5[4][46] , \g5[4][45] , \g5[4][44] , \g5[4][43] , 
        \g5[4][42] , \g5[4][41] , \g5[4][40] , \g5[4][39] , \g5[4][38] , 
        \g5[4][37] , \g5[4][36] , \g5[4][35] , \g5[4][34] , \g5[4][33] , 
        \g5[4][32] , \g5[4][31] , \g5[4][30] , \g5[4][29] , \g5[4][28] , 
        \g5[4][27] , \g5[4][26] , \g5[4][25] , \g5[4][24] , \g5[4][23] , 
        \g5[4][22] , \g5[4][21] , \g5[4][20] , \g5[4][19] , \g5[4][18] , 
        \g5[4][17] , \g5[4][16] , \g5[4][15] , \g5[4][14] , \g5[4][13] , 
        \g5[4][12] , \g5[4][11] , \g5[4][10] , \g5[4][9] , \g5[4][8] , 
        \g5[4][7] , \g5[4][6] , \g5[4][5] , \g5[4][4] , \g5[4][3] , \g5[4][2] , 
        \g5[4][1] , SYNOPSYS_UNCONNECTED__50}) );
  FullAdder_11 \level5[1].x2  ( .a({\g4[3][63] , \g4[3][62] , \g4[3][61] , 
        \g4[3][60] , \g4[3][59] , \g4[3][58] , \g4[3][57] , \g4[3][56] , 
        \g4[3][55] , \g4[3][54] , \g4[3][53] , \g4[3][52] , \g4[3][51] , 
        \g4[3][50] , \g4[3][49] , \g4[3][48] , \g4[3][47] , \g4[3][46] , 
        \g4[3][45] , \g4[3][44] , \g4[3][43] , \g4[3][42] , \g4[3][41] , 
        \g4[3][40] , \g4[3][39] , \g4[3][38] , \g4[3][37] , \g4[3][36] , 
        \g4[3][35] , \g4[3][34] , \g4[3][33] , \g4[3][32] , \g4[3][31] , 
        \g4[3][30] , \g4[3][29] , \g4[3][28] , \g4[3][27] , \g4[3][26] , 
        \g4[3][25] , \g4[3][24] , \g4[3][23] , \g4[3][22] , \g4[3][21] , 
        \g4[3][20] , \g4[3][19] , \g4[3][18] , \g4[3][17] , \g4[3][16] , 
        \g4[3][15] , \g4[3][14] , \g4[3][13] , \g4[3][12] , \g4[3][11] , 
        \g4[3][10] , \g4[3][9] , \g4[3][8] , \g4[3][7] , \g4[3][6] , 
        \g4[3][5] , \g4[3][4] , \g4[3][3] , \g4[3][2] , \g4[3][1] , \g4[3][0] }), .b({\g4[4][63] , \g4[4][62] , \g4[4][61] , \g4[4][60] , \g4[4][59] , 
        \g4[4][58] , \g4[4][57] , \g4[4][56] , \g4[4][55] , \g4[4][54] , 
        \g4[4][53] , \g4[4][52] , \g4[4][51] , \g4[4][50] , \g4[4][49] , 
        \g4[4][48] , \g4[4][47] , \g4[4][46] , \g4[4][45] , \g4[4][44] , 
        \g4[4][43] , \g4[4][42] , \g4[4][41] , \g4[4][40] , \g4[4][39] , 
        \g4[4][38] , \g4[4][37] , \g4[4][36] , \g4[4][35] , \g4[4][34] , 
        \g4[4][33] , \g4[4][32] , \g4[4][31] , \g4[4][30] , \g4[4][29] , 
        \g4[4][28] , \g4[4][27] , \g4[4][26] , \g4[4][25] , \g4[4][24] , 
        \g4[4][23] , \g4[4][22] , \g4[4][21] , \g4[4][20] , \g4[4][19] , 
        \g4[4][18] , \g4[4][17] , \g4[4][16] , \g4[4][15] , \g4[4][14] , 
        \g4[4][13] , \g4[4][12] , \g4[4][11] , \g4[4][10] , \g4[4][9] , 
        \g4[4][8] , \g4[4][7] , \g4[4][6] , \g4[4][5] , \g4[4][4] , \g4[4][3] , 
        \g4[4][2] , \g4[4][1] , \g4[4][0] }), .cin({\g4[5][63] , \g4[5][62] , 
        \g4[5][61] , \g4[5][60] , \g4[5][59] , \g4[5][58] , \g4[5][57] , 
        \g4[5][56] , \g4[5][55] , \g4[5][54] , \g4[5][53] , \g4[5][52] , 
        \g4[5][51] , \g4[5][50] , \g4[5][49] , \g4[5][48] , \g4[5][47] , 
        \g4[5][46] , \g4[5][45] , \g4[5][44] , \g4[5][43] , \g4[5][42] , 
        \g4[5][41] , \g4[5][40] , \g4[5][39] , \g4[5][38] , \g4[5][37] , 
        \g4[5][36] , \g4[5][35] , \g4[5][34] , \g4[5][33] , \g4[5][32] , 
        \g4[5][31] , \g4[5][30] , \g4[5][29] , \g4[5][28] , \g4[5][27] , 
        \g4[5][26] , \g4[5][25] , \g4[5][24] , \g4[5][23] , \g4[5][22] , 
        \g4[5][21] , \g4[5][20] , \g4[5][19] , \g4[5][18] , \g4[5][17] , 
        \g4[5][16] , \g4[5][15] , \g4[5][14] , \g4[5][13] , \g4[5][12] , 
        \g4[5][11] , \g4[5][10] , \g4[5][9] , \g4[5][8] , \g4[5][7] , 
        \g4[5][6] , \g4[5][5] , \g4[5][4] , \g4[5][3] , \g4[5][2] , \g4[5][1] , 
        \g4[5][0] }), .sum({\g5[1][63] , \g5[1][62] , \g5[1][61] , \g5[1][60] , 
        \g5[1][59] , \g5[1][58] , \g5[1][57] , \g5[1][56] , \g5[1][55] , 
        \g5[1][54] , \g5[1][53] , \g5[1][52] , \g5[1][51] , \g5[1][50] , 
        \g5[1][49] , \g5[1][48] , \g5[1][47] , \g5[1][46] , \g5[1][45] , 
        \g5[1][44] , \g5[1][43] , \g5[1][42] , \g5[1][41] , \g5[1][40] , 
        \g5[1][39] , \g5[1][38] , \g5[1][37] , \g5[1][36] , \g5[1][35] , 
        \g5[1][34] , \g5[1][33] , \g5[1][32] , \g5[1][31] , \g5[1][30] , 
        \g5[1][29] , \g5[1][28] , \g5[1][27] , \g5[1][26] , \g5[1][25] , 
        \g5[1][24] , \g5[1][23] , \g5[1][22] , \g5[1][21] , \g5[1][20] , 
        \g5[1][19] , \g5[1][18] , \g5[1][17] , \g5[1][16] , \g5[1][15] , 
        \g5[1][14] , \g5[1][13] , \g5[1][12] , \g5[1][11] , \g5[1][10] , 
        \g5[1][9] , \g5[1][8] , \g5[1][7] , \g5[1][6] , \g5[1][5] , \g5[1][4] , 
        \g5[1][3] , \g5[1][2] , \g5[1][1] , \g5[1][0] }), .cout({\g5[5][63] , 
        \g5[5][62] , \g5[5][61] , \g5[5][60] , \g5[5][59] , \g5[5][58] , 
        \g5[5][57] , \g5[5][56] , \g5[5][55] , \g5[5][54] , \g5[5][53] , 
        \g5[5][52] , \g5[5][51] , \g5[5][50] , \g5[5][49] , \g5[5][48] , 
        \g5[5][47] , \g5[5][46] , \g5[5][45] , \g5[5][44] , \g5[5][43] , 
        \g5[5][42] , \g5[5][41] , \g5[5][40] , \g5[5][39] , \g5[5][38] , 
        \g5[5][37] , \g5[5][36] , \g5[5][35] , \g5[5][34] , \g5[5][33] , 
        \g5[5][32] , \g5[5][31] , \g5[5][30] , \g5[5][29] , \g5[5][28] , 
        \g5[5][27] , \g5[5][26] , \g5[5][25] , \g5[5][24] , \g5[5][23] , 
        \g5[5][22] , \g5[5][21] , \g5[5][20] , \g5[5][19] , \g5[5][18] , 
        \g5[5][17] , \g5[5][16] , \g5[5][15] , \g5[5][14] , \g5[5][13] , 
        \g5[5][12] , \g5[5][11] , \g5[5][10] , \g5[5][9] , \g5[5][8] , 
        \g5[5][7] , \g5[5][6] , \g5[5][5] , \g5[5][4] , \g5[5][3] , \g5[5][2] , 
        \g5[5][1] , SYNOPSYS_UNCONNECTED__51}) );
  FullAdder_10 \level5[2].x2  ( .a({\g4[6][63] , \g4[6][62] , \g4[6][61] , 
        \g4[6][60] , \g4[6][59] , \g4[6][58] , \g4[6][57] , \g4[6][56] , 
        \g4[6][55] , \g4[6][54] , \g4[6][53] , \g4[6][52] , \g4[6][51] , 
        \g4[6][50] , \g4[6][49] , \g4[6][48] , \g4[6][47] , \g4[6][46] , 
        \g4[6][45] , \g4[6][44] , \g4[6][43] , \g4[6][42] , \g4[6][41] , 
        \g4[6][40] , \g4[6][39] , \g4[6][38] , \g4[6][37] , \g4[6][36] , 
        \g4[6][35] , \g4[6][34] , \g4[6][33] , \g4[6][32] , \g4[6][31] , 
        \g4[6][30] , \g4[6][29] , \g4[6][28] , \g4[6][27] , \g4[6][26] , 
        \g4[6][25] , \g4[6][24] , \g4[6][23] , \g4[6][22] , \g4[6][21] , 
        \g4[6][20] , \g4[6][19] , \g4[6][18] , \g4[6][17] , \g4[6][16] , 
        \g4[6][15] , \g4[6][14] , \g4[6][13] , \g4[6][12] , \g4[6][11] , 
        \g4[6][10] , \g4[6][9] , \g4[6][8] , \g4[6][7] , \g4[6][6] , 
        \g4[6][5] , \g4[6][4] , \g4[6][3] , \g4[6][2] , \g4[6][1] , 1'b0}), 
        .b({\g4[7][63] , \g4[7][62] , \g4[7][61] , \g4[7][60] , \g4[7][59] , 
        \g4[7][58] , \g4[7][57] , \g4[7][56] , \g4[7][55] , \g4[7][54] , 
        \g4[7][53] , \g4[7][52] , \g4[7][51] , \g4[7][50] , \g4[7][49] , 
        \g4[7][48] , \g4[7][47] , \g4[7][46] , \g4[7][45] , \g4[7][44] , 
        \g4[7][43] , \g4[7][42] , \g4[7][41] , \g4[7][40] , \g4[7][39] , 
        \g4[7][38] , \g4[7][37] , \g4[7][36] , \g4[7][35] , \g4[7][34] , 
        \g4[7][33] , \g4[7][32] , \g4[7][31] , \g4[7][30] , \g4[7][29] , 
        \g4[7][28] , \g4[7][27] , \g4[7][26] , \g4[7][25] , \g4[7][24] , 
        \g4[7][23] , \g4[7][22] , \g4[7][21] , \g4[7][20] , \g4[7][19] , 
        \g4[7][18] , \g4[7][17] , \g4[7][16] , \g4[7][15] , \g4[7][14] , 
        \g4[7][13] , \g4[7][12] , \g4[7][11] , \g4[7][10] , \g4[7][9] , 
        \g4[7][8] , \g4[7][7] , \g4[7][6] , \g4[7][5] , \g4[7][4] , \g4[7][3] , 
        \g4[7][2] , \g4[7][1] , 1'b0}), .cin({\g4[8][63] , \g4[8][62] , 
        \g4[8][61] , \g4[8][60] , \g4[8][59] , \g4[8][58] , \g4[8][57] , 
        \g4[8][56] , \g4[8][55] , \g4[8][54] , \g4[8][53] , \g4[8][52] , 
        \g4[8][51] , \g4[8][50] , \g4[8][49] , \g4[8][48] , \g4[8][47] , 
        \g4[8][46] , \g4[8][45] , \g4[8][44] , \g4[8][43] , \g4[8][42] , 
        \g4[8][41] , \g4[8][40] , \g4[8][39] , \g4[8][38] , \g4[8][37] , 
        \g4[8][36] , \g4[8][35] , \g4[8][34] , \g4[8][33] , \g4[8][32] , 
        \g4[8][31] , \g4[8][30] , \g4[8][29] , \g4[8][28] , \g4[8][27] , 
        \g4[8][26] , \g4[8][25] , \g4[8][24] , \g4[8][23] , \g4[8][22] , 
        \g4[8][21] , \g4[8][20] , \g4[8][19] , \g4[8][18] , \g4[8][17] , 
        \g4[8][16] , \g4[8][15] , \g4[8][14] , \g4[8][13] , \g4[8][12] , 
        \g4[8][11] , \g4[8][10] , \g4[8][9] , \g4[8][8] , \g4[8][7] , 
        \g4[8][6] , \g4[8][5] , \g4[8][4] , \g4[8][3] , \g4[8][2] , \g4[8][1] , 
        1'b0}), .sum({\g5[2][63] , \g5[2][62] , \g5[2][61] , \g5[2][60] , 
        \g5[2][59] , \g5[2][58] , \g5[2][57] , \g5[2][56] , \g5[2][55] , 
        \g5[2][54] , \g5[2][53] , \g5[2][52] , \g5[2][51] , \g5[2][50] , 
        \g5[2][49] , \g5[2][48] , \g5[2][47] , \g5[2][46] , \g5[2][45] , 
        \g5[2][44] , \g5[2][43] , \g5[2][42] , \g5[2][41] , \g5[2][40] , 
        \g5[2][39] , \g5[2][38] , \g5[2][37] , \g5[2][36] , \g5[2][35] , 
        \g5[2][34] , \g5[2][33] , \g5[2][32] , \g5[2][31] , \g5[2][30] , 
        \g5[2][29] , \g5[2][28] , \g5[2][27] , \g5[2][26] , \g5[2][25] , 
        \g5[2][24] , \g5[2][23] , \g5[2][22] , \g5[2][21] , \g5[2][20] , 
        \g5[2][19] , \g5[2][18] , \g5[2][17] , \g5[2][16] , \g5[2][15] , 
        \g5[2][14] , \g5[2][13] , \g5[2][12] , \g5[2][11] , \g5[2][10] , 
        \g5[2][9] , \g5[2][8] , \g5[2][7] , \g5[2][6] , \g5[2][5] , \g5[2][4] , 
        \g5[2][3] , \g5[2][2] , \g5[2][1] , \g5[2][0] }), .cout({\g5[6][63] , 
        \g5[6][62] , \g5[6][61] , \g5[6][60] , \g5[6][59] , \g5[6][58] , 
        \g5[6][57] , \g5[6][56] , \g5[6][55] , \g5[6][54] , \g5[6][53] , 
        \g5[6][52] , \g5[6][51] , \g5[6][50] , \g5[6][49] , \g5[6][48] , 
        \g5[6][47] , \g5[6][46] , \g5[6][45] , \g5[6][44] , \g5[6][43] , 
        \g5[6][42] , \g5[6][41] , \g5[6][40] , \g5[6][39] , \g5[6][38] , 
        \g5[6][37] , \g5[6][36] , \g5[6][35] , \g5[6][34] , \g5[6][33] , 
        \g5[6][32] , \g5[6][31] , \g5[6][30] , \g5[6][29] , \g5[6][28] , 
        \g5[6][27] , \g5[6][26] , \g5[6][25] , \g5[6][24] , \g5[6][23] , 
        \g5[6][22] , \g5[6][21] , \g5[6][20] , \g5[6][19] , \g5[6][18] , 
        \g5[6][17] , \g5[6][16] , \g5[6][15] , \g5[6][14] , \g5[6][13] , 
        \g5[6][12] , \g5[6][11] , \g5[6][10] , \g5[6][9] , \g5[6][8] , 
        \g5[6][7] , \g5[6][6] , \g5[6][5] , \g5[6][4] , \g5[6][3] , \g5[6][2] , 
        \g5[6][1] , SYNOPSYS_UNCONNECTED__52}) );
  FullAdder_9 \level5[3].x2  ( .a({\g4[9][63] , \g4[9][62] , \g4[9][61] , 
        \g4[9][60] , \g4[9][59] , \g4[9][58] , \g4[9][57] , \g4[9][56] , 
        \g4[9][55] , \g4[9][54] , \g4[9][53] , \g4[9][52] , \g4[9][51] , 
        \g4[9][50] , \g4[9][49] , \g4[9][48] , \g4[9][47] , \g4[9][46] , 
        \g4[9][45] , \g4[9][44] , \g4[9][43] , \g4[9][42] , \g4[9][41] , 
        \g4[9][40] , \g4[9][39] , \g4[9][38] , \g4[9][37] , \g4[9][36] , 
        \g4[9][35] , \g4[9][34] , \g4[9][33] , \g4[9][32] , \g4[9][31] , 
        \g4[9][30] , \g4[9][29] , \g4[9][28] , \g4[9][27] , \g4[9][26] , 
        \g4[9][25] , \g4[9][24] , \g4[9][23] , \g4[9][22] , \g4[9][21] , 
        \g4[9][20] , \g4[9][19] , \g4[9][18] , \g4[9][17] , \g4[9][16] , 
        \g4[9][15] , \g4[9][14] , \g4[9][13] , \g4[9][12] , \g4[9][11] , 
        \g4[9][10] , \g4[9][9] , \g4[9][8] , \g4[9][7] , \g4[9][6] , 
        \g4[9][5] , \g4[9][4] , \g4[9][3] , \g4[9][2] , \g4[9][1] , 1'b0}), 
        .b({\g4[10][63] , \g4[10][62] , \g4[10][61] , \g4[10][60] , 
        \g4[10][59] , \g4[10][58] , \g4[10][57] , \g4[10][56] , \g4[10][55] , 
        \g4[10][54] , \g4[10][53] , \g4[10][52] , \g4[10][51] , \g4[10][50] , 
        \g4[10][49] , \g4[10][48] , \g4[10][47] , \g4[10][46] , \g4[10][45] , 
        \g4[10][44] , \g4[10][43] , \g4[10][42] , \g4[10][41] , \g4[10][40] , 
        \g4[10][39] , \g4[10][38] , \g4[10][37] , \g4[10][36] , \g4[10][35] , 
        \g4[10][34] , \g4[10][33] , \g4[10][32] , \g4[10][31] , \g4[10][30] , 
        \g4[10][29] , \g4[10][28] , \g4[10][27] , \g4[10][26] , \g4[10][25] , 
        \g4[10][24] , \g4[10][23] , \g4[10][22] , \g4[10][21] , \g4[10][20] , 
        \g4[10][19] , \g4[10][18] , \g4[10][17] , \g4[10][16] , \g4[10][15] , 
        \g4[10][14] , \g4[10][13] , \g4[10][12] , \g4[10][11] , \g4[10][10] , 
        \g4[10][9] , \g4[10][8] , \g4[10][7] , \g4[10][6] , \g4[10][5] , 
        \g4[10][4] , \g4[10][3] , \g4[10][2] , \g4[10][1] , 1'b0}), .cin({
        \g4[11][63] , \g4[11][62] , \g4[11][61] , \g4[11][60] , \g4[11][59] , 
        \g4[11][58] , \g4[11][57] , \g4[11][56] , \g4[11][55] , \g4[11][54] , 
        \g4[11][53] , \g4[11][52] , \g4[11][51] , \g4[11][50] , \g4[11][49] , 
        \g4[11][48] , \g4[11][47] , \g4[11][46] , \g4[11][45] , \g4[11][44] , 
        \g4[11][43] , \g4[11][42] , \g4[11][41] , \g4[11][40] , \g4[11][39] , 
        \g4[11][38] , \g4[11][37] , \g4[11][36] , \g4[11][35] , \g4[11][34] , 
        \g4[11][33] , \g4[11][32] , \g4[11][31] , \g4[11][30] , \g4[11][29] , 
        \g4[11][28] , \g4[11][27] , \g4[11][26] , \g4[11][25] , \g4[11][24] , 
        \g4[11][23] , \g4[11][22] , \g4[11][21] , \g4[11][20] , \g4[11][19] , 
        \g4[11][18] , \g4[11][17] , \g4[11][16] , \g4[11][15] , \g4[11][14] , 
        \g4[11][13] , \g4[11][12] , \g4[11][11] , \g4[11][10] , \g4[11][9] , 
        \g4[11][8] , \g4[11][7] , \g4[11][6] , \g4[11][5] , \g4[11][4] , 
        \g4[11][3] , \g4[11][2] , \g4[11][1] , 1'b0}), .sum({\g5[3][63] , 
        \g5[3][62] , \g5[3][61] , \g5[3][60] , \g5[3][59] , \g5[3][58] , 
        \g5[3][57] , \g5[3][56] , \g5[3][55] , \g5[3][54] , \g5[3][53] , 
        \g5[3][52] , \g5[3][51] , \g5[3][50] , \g5[3][49] , \g5[3][48] , 
        \g5[3][47] , \g5[3][46] , \g5[3][45] , \g5[3][44] , \g5[3][43] , 
        \g5[3][42] , \g5[3][41] , \g5[3][40] , \g5[3][39] , \g5[3][38] , 
        \g5[3][37] , \g5[3][36] , \g5[3][35] , \g5[3][34] , \g5[3][33] , 
        \g5[3][32] , \g5[3][31] , \g5[3][30] , \g5[3][29] , \g5[3][28] , 
        \g5[3][27] , \g5[3][26] , \g5[3][25] , \g5[3][24] , \g5[3][23] , 
        \g5[3][22] , \g5[3][21] , \g5[3][20] , \g5[3][19] , \g5[3][18] , 
        \g5[3][17] , \g5[3][16] , \g5[3][15] , \g5[3][14] , \g5[3][13] , 
        \g5[3][12] , \g5[3][11] , \g5[3][10] , \g5[3][9] , \g5[3][8] , 
        \g5[3][7] , \g5[3][6] , \g5[3][5] , \g5[3][4] , \g5[3][3] , \g5[3][2] , 
        \g5[3][1] , \g5[3][0] }), .cout({\g5[7][63] , \g5[7][62] , \g5[7][61] , 
        \g5[7][60] , \g5[7][59] , \g5[7][58] , \g5[7][57] , \g5[7][56] , 
        \g5[7][55] , \g5[7][54] , \g5[7][53] , \g5[7][52] , \g5[7][51] , 
        \g5[7][50] , \g5[7][49] , \g5[7][48] , \g5[7][47] , \g5[7][46] , 
        \g5[7][45] , \g5[7][44] , \g5[7][43] , \g5[7][42] , \g5[7][41] , 
        \g5[7][40] , \g5[7][39] , \g5[7][38] , \g5[7][37] , \g5[7][36] , 
        \g5[7][35] , \g5[7][34] , \g5[7][33] , \g5[7][32] , \g5[7][31] , 
        \g5[7][30] , \g5[7][29] , \g5[7][28] , \g5[7][27] , \g5[7][26] , 
        \g5[7][25] , \g5[7][24] , \g5[7][23] , \g5[7][22] , \g5[7][21] , 
        \g5[7][20] , \g5[7][19] , \g5[7][18] , \g5[7][17] , \g5[7][16] , 
        \g5[7][15] , \g5[7][14] , \g5[7][13] , \g5[7][12] , \g5[7][11] , 
        \g5[7][10] , \g5[7][9] , \g5[7][8] , \g5[7][7] , \g5[7][6] , 
        \g5[7][5] , \g5[7][4] , \g5[7][3] , \g5[7][2] , \g5[7][1] , 
        SYNOPSYS_UNCONNECTED__53}) );
  FullAdder_8 F0 ( .a({\g5[0][63] , \g5[0][62] , \g5[0][61] , \g5[0][60] , 
        \g5[0][59] , \g5[0][58] , \g5[0][57] , \g5[0][56] , \g5[0][55] , 
        \g5[0][54] , \g5[0][53] , \g5[0][52] , \g5[0][51] , \g5[0][50] , 
        \g5[0][49] , \g5[0][48] , \g5[0][47] , \g5[0][46] , \g5[0][45] , 
        \g5[0][44] , \g5[0][43] , \g5[0][42] , \g5[0][41] , \g5[0][40] , 
        \g5[0][39] , \g5[0][38] , \g5[0][37] , \g5[0][36] , \g5[0][35] , 
        \g5[0][34] , \g5[0][33] , \g5[0][32] , \g5[0][31] , \g5[0][30] , 
        \g5[0][29] , \g5[0][28] , \g5[0][27] , \g5[0][26] , \g5[0][25] , 
        \g5[0][24] , \g5[0][23] , \g5[0][22] , \g5[0][21] , \g5[0][20] , 
        \g5[0][19] , \g5[0][18] , \g5[0][17] , \g5[0][16] , \g5[0][15] , 
        \g5[0][14] , \g5[0][13] , \g5[0][12] , \g5[0][11] , \g5[0][10] , 
        \g5[0][9] , \g5[0][8] , \g5[0][7] , \g5[0][6] , \g5[0][5] , \g5[0][4] , 
        \g5[0][3] , \g5[0][2] , \g5[0][1] , \g5[0][0] }), .b({\g5[1][63] , 
        \g5[1][62] , \g5[1][61] , \g5[1][60] , \g5[1][59] , \g5[1][58] , 
        \g5[1][57] , \g5[1][56] , \g5[1][55] , \g5[1][54] , \g5[1][53] , 
        \g5[1][52] , \g5[1][51] , \g5[1][50] , \g5[1][49] , \g5[1][48] , 
        \g5[1][47] , \g5[1][46] , \g5[1][45] , \g5[1][44] , \g5[1][43] , 
        \g5[1][42] , \g5[1][41] , \g5[1][40] , \g5[1][39] , \g5[1][38] , 
        \g5[1][37] , \g5[1][36] , \g5[1][35] , \g5[1][34] , \g5[1][33] , 
        \g5[1][32] , \g5[1][31] , \g5[1][30] , \g5[1][29] , \g5[1][28] , 
        \g5[1][27] , \g5[1][26] , \g5[1][25] , \g5[1][24] , \g5[1][23] , 
        \g5[1][22] , \g5[1][21] , \g5[1][20] , \g5[1][19] , \g5[1][18] , 
        \g5[1][17] , \g5[1][16] , \g5[1][15] , \g5[1][14] , \g5[1][13] , 
        \g5[1][12] , \g5[1][11] , \g5[1][10] , \g5[1][9] , \g5[1][8] , 
        \g5[1][7] , \g5[1][6] , \g5[1][5] , \g5[1][4] , \g5[1][3] , \g5[1][2] , 
        \g5[1][1] , \g5[1][0] }), .cin({\g5[2][63] , \g5[2][62] , \g5[2][61] , 
        \g5[2][60] , \g5[2][59] , \g5[2][58] , \g5[2][57] , \g5[2][56] , 
        \g5[2][55] , \g5[2][54] , \g5[2][53] , \g5[2][52] , \g5[2][51] , 
        \g5[2][50] , \g5[2][49] , \g5[2][48] , \g5[2][47] , \g5[2][46] , 
        \g5[2][45] , \g5[2][44] , \g5[2][43] , \g5[2][42] , \g5[2][41] , 
        \g5[2][40] , \g5[2][39] , \g5[2][38] , \g5[2][37] , \g5[2][36] , 
        \g5[2][35] , \g5[2][34] , \g5[2][33] , \g5[2][32] , \g5[2][31] , 
        \g5[2][30] , \g5[2][29] , \g5[2][28] , \g5[2][27] , \g5[2][26] , 
        \g5[2][25] , \g5[2][24] , \g5[2][23] , \g5[2][22] , \g5[2][21] , 
        \g5[2][20] , \g5[2][19] , \g5[2][18] , \g5[2][17] , \g5[2][16] , 
        \g5[2][15] , \g5[2][14] , \g5[2][13] , \g5[2][12] , \g5[2][11] , 
        \g5[2][10] , \g5[2][9] , \g5[2][8] , \g5[2][7] , \g5[2][6] , 
        \g5[2][5] , \g5[2][4] , \g5[2][3] , \g5[2][2] , \g5[2][1] , \g5[2][0] }), .sum({\g6[0][63] , \g6[0][62] , \g6[0][61] , \g6[0][60] , \g6[0][59] , 
        \g6[0][58] , \g6[0][57] , \g6[0][56] , \g6[0][55] , \g6[0][54] , 
        \g6[0][53] , \g6[0][52] , \g6[0][51] , \g6[0][50] , \g6[0][49] , 
        \g6[0][48] , \g6[0][47] , \g6[0][46] , \g6[0][45] , \g6[0][44] , 
        \g6[0][43] , \g6[0][42] , \g6[0][41] , \g6[0][40] , \g6[0][39] , 
        \g6[0][38] , \g6[0][37] , \g6[0][36] , \g6[0][35] , \g6[0][34] , 
        \g6[0][33] , \g6[0][32] , \g6[0][31] , \g6[0][30] , \g6[0][29] , 
        \g6[0][28] , \g6[0][27] , \g6[0][26] , \g6[0][25] , \g6[0][24] , 
        \g6[0][23] , \g6[0][22] , \g6[0][21] , \g6[0][20] , \g6[0][19] , 
        \g6[0][18] , \g6[0][17] , \g6[0][16] , \g6[0][15] , \g6[0][14] , 
        \g6[0][13] , \g6[0][12] , \g6[0][11] , \g6[0][10] , \g6[0][9] , 
        \g6[0][8] , \g6[0][7] , \g6[0][6] , \g6[0][5] , \g6[0][4] , \g6[0][3] , 
        \g6[0][2] , \g6[0][1] , \g6[0][0] }), .cout({\g6[1][63] , \g6[1][62] , 
        \g6[1][61] , \g6[1][60] , \g6[1][59] , \g6[1][58] , \g6[1][57] , 
        \g6[1][56] , \g6[1][55] , \g6[1][54] , \g6[1][53] , \g6[1][52] , 
        \g6[1][51] , \g6[1][50] , \g6[1][49] , \g6[1][48] , \g6[1][47] , 
        \g6[1][46] , \g6[1][45] , \g6[1][44] , \g6[1][43] , \g6[1][42] , 
        \g6[1][41] , \g6[1][40] , \g6[1][39] , \g6[1][38] , \g6[1][37] , 
        \g6[1][36] , \g6[1][35] , \g6[1][34] , \g6[1][33] , \g6[1][32] , 
        \g6[1][31] , \g6[1][30] , \g6[1][29] , \g6[1][28] , \g6[1][27] , 
        \g6[1][26] , \g6[1][25] , \g6[1][24] , \g6[1][23] , \g6[1][22] , 
        \g6[1][21] , \g6[1][20] , \g6[1][19] , \g6[1][18] , \g6[1][17] , 
        \g6[1][16] , \g6[1][15] , \g6[1][14] , \g6[1][13] , \g6[1][12] , 
        \g6[1][11] , \g6[1][10] , \g6[1][9] , \g6[1][8] , \g6[1][7] , 
        \g6[1][6] , \g6[1][5] , \g6[1][4] , \g6[1][3] , \g6[1][2] , \g6[1][1] , 
        SYNOPSYS_UNCONNECTED__54}) );
  FullAdder_7 F1 ( .a({\g5[3][63] , \g5[3][62] , \g5[3][61] , \g5[3][60] , 
        \g5[3][59] , \g5[3][58] , \g5[3][57] , \g5[3][56] , \g5[3][55] , 
        \g5[3][54] , \g5[3][53] , \g5[3][52] , \g5[3][51] , \g5[3][50] , 
        \g5[3][49] , \g5[3][48] , \g5[3][47] , \g5[3][46] , \g5[3][45] , 
        \g5[3][44] , \g5[3][43] , \g5[3][42] , \g5[3][41] , \g5[3][40] , 
        \g5[3][39] , \g5[3][38] , \g5[3][37] , \g5[3][36] , \g5[3][35] , 
        \g5[3][34] , \g5[3][33] , \g5[3][32] , \g5[3][31] , \g5[3][30] , 
        \g5[3][29] , \g5[3][28] , \g5[3][27] , \g5[3][26] , \g5[3][25] , 
        \g5[3][24] , \g5[3][23] , \g5[3][22] , \g5[3][21] , \g5[3][20] , 
        \g5[3][19] , \g5[3][18] , \g5[3][17] , \g5[3][16] , \g5[3][15] , 
        \g5[3][14] , \g5[3][13] , \g5[3][12] , \g5[3][11] , \g5[3][10] , 
        \g5[3][9] , \g5[3][8] , \g5[3][7] , \g5[3][6] , \g5[3][5] , \g5[3][4] , 
        \g5[3][3] , \g5[3][2] , \g5[3][1] , \g5[3][0] }), .b({\g5[4][63] , 
        \g5[4][62] , \g5[4][61] , \g5[4][60] , \g5[4][59] , \g5[4][58] , 
        \g5[4][57] , \g5[4][56] , \g5[4][55] , \g5[4][54] , \g5[4][53] , 
        \g5[4][52] , \g5[4][51] , \g5[4][50] , \g5[4][49] , \g5[4][48] , 
        \g5[4][47] , \g5[4][46] , \g5[4][45] , \g5[4][44] , \g5[4][43] , 
        \g5[4][42] , \g5[4][41] , \g5[4][40] , \g5[4][39] , \g5[4][38] , 
        \g5[4][37] , \g5[4][36] , \g5[4][35] , \g5[4][34] , \g5[4][33] , 
        \g5[4][32] , \g5[4][31] , \g5[4][30] , \g5[4][29] , \g5[4][28] , 
        \g5[4][27] , \g5[4][26] , \g5[4][25] , \g5[4][24] , \g5[4][23] , 
        \g5[4][22] , \g5[4][21] , \g5[4][20] , \g5[4][19] , \g5[4][18] , 
        \g5[4][17] , \g5[4][16] , \g5[4][15] , \g5[4][14] , \g5[4][13] , 
        \g5[4][12] , \g5[4][11] , \g5[4][10] , \g5[4][9] , \g5[4][8] , 
        \g5[4][7] , \g5[4][6] , \g5[4][5] , \g5[4][4] , \g5[4][3] , \g5[4][2] , 
        \g5[4][1] , 1'b0}), .cin({\g5[5][63] , \g5[5][62] , \g5[5][61] , 
        \g5[5][60] , \g5[5][59] , \g5[5][58] , \g5[5][57] , \g5[5][56] , 
        \g5[5][55] , \g5[5][54] , \g5[5][53] , \g5[5][52] , \g5[5][51] , 
        \g5[5][50] , \g5[5][49] , \g5[5][48] , \g5[5][47] , \g5[5][46] , 
        \g5[5][45] , \g5[5][44] , \g5[5][43] , \g5[5][42] , \g5[5][41] , 
        \g5[5][40] , \g5[5][39] , \g5[5][38] , \g5[5][37] , \g5[5][36] , 
        \g5[5][35] , \g5[5][34] , \g5[5][33] , \g5[5][32] , \g5[5][31] , 
        \g5[5][30] , \g5[5][29] , \g5[5][28] , \g5[5][27] , \g5[5][26] , 
        \g5[5][25] , \g5[5][24] , \g5[5][23] , \g5[5][22] , \g5[5][21] , 
        \g5[5][20] , \g5[5][19] , \g5[5][18] , \g5[5][17] , \g5[5][16] , 
        \g5[5][15] , \g5[5][14] , \g5[5][13] , \g5[5][12] , \g5[5][11] , 
        \g5[5][10] , \g5[5][9] , \g5[5][8] , \g5[5][7] , \g5[5][6] , 
        \g5[5][5] , \g5[5][4] , \g5[5][3] , \g5[5][2] , \g5[5][1] , 1'b0}), 
        .sum({\g6[2][63] , \g6[2][62] , \g6[2][61] , \g6[2][60] , \g6[2][59] , 
        \g6[2][58] , \g6[2][57] , \g6[2][56] , \g6[2][55] , \g6[2][54] , 
        \g6[2][53] , \g6[2][52] , \g6[2][51] , \g6[2][50] , \g6[2][49] , 
        \g6[2][48] , \g6[2][47] , \g6[2][46] , \g6[2][45] , \g6[2][44] , 
        \g6[2][43] , \g6[2][42] , \g6[2][41] , \g6[2][40] , \g6[2][39] , 
        \g6[2][38] , \g6[2][37] , \g6[2][36] , \g6[2][35] , \g6[2][34] , 
        \g6[2][33] , \g6[2][32] , \g6[2][31] , \g6[2][30] , \g6[2][29] , 
        \g6[2][28] , \g6[2][27] , \g6[2][26] , \g6[2][25] , \g6[2][24] , 
        \g6[2][23] , \g6[2][22] , \g6[2][21] , \g6[2][20] , \g6[2][19] , 
        \g6[2][18] , \g6[2][17] , \g6[2][16] , \g6[2][15] , \g6[2][14] , 
        \g6[2][13] , \g6[2][12] , \g6[2][11] , \g6[2][10] , \g6[2][9] , 
        \g6[2][8] , \g6[2][7] , \g6[2][6] , \g6[2][5] , \g6[2][4] , \g6[2][3] , 
        \g6[2][2] , \g6[2][1] , \g6[2][0] }), .cout({\g6[3][63] , \g6[3][62] , 
        \g6[3][61] , \g6[3][60] , \g6[3][59] , \g6[3][58] , \g6[3][57] , 
        \g6[3][56] , \g6[3][55] , \g6[3][54] , \g6[3][53] , \g6[3][52] , 
        \g6[3][51] , \g6[3][50] , \g6[3][49] , \g6[3][48] , \g6[3][47] , 
        \g6[3][46] , \g6[3][45] , \g6[3][44] , \g6[3][43] , \g6[3][42] , 
        \g6[3][41] , \g6[3][40] , \g6[3][39] , \g6[3][38] , \g6[3][37] , 
        \g6[3][36] , \g6[3][35] , \g6[3][34] , \g6[3][33] , \g6[3][32] , 
        \g6[3][31] , \g6[3][30] , \g6[3][29] , \g6[3][28] , \g6[3][27] , 
        \g6[3][26] , \g6[3][25] , \g6[3][24] , \g6[3][23] , \g6[3][22] , 
        \g6[3][21] , \g6[3][20] , \g6[3][19] , \g6[3][18] , \g6[3][17] , 
        \g6[3][16] , \g6[3][15] , \g6[3][14] , \g6[3][13] , \g6[3][12] , 
        \g6[3][11] , \g6[3][10] , \g6[3][9] , \g6[3][8] , \g6[3][7] , 
        \g6[3][6] , \g6[3][5] , \g6[3][4] , \g6[3][3] , \g6[3][2] , \g6[3][1] , 
        SYNOPSYS_UNCONNECTED__55}) );
  FullAdder_6 F2 ( .a({\g5[6][63] , \g5[6][62] , \g5[6][61] , \g5[6][60] , 
        \g5[6][59] , \g5[6][58] , \g5[6][57] , \g5[6][56] , \g5[6][55] , 
        \g5[6][54] , \g5[6][53] , \g5[6][52] , \g5[6][51] , \g5[6][50] , 
        \g5[6][49] , \g5[6][48] , \g5[6][47] , \g5[6][46] , \g5[6][45] , 
        \g5[6][44] , \g5[6][43] , \g5[6][42] , \g5[6][41] , \g5[6][40] , 
        \g5[6][39] , \g5[6][38] , \g5[6][37] , \g5[6][36] , \g5[6][35] , 
        \g5[6][34] , \g5[6][33] , \g5[6][32] , \g5[6][31] , \g5[6][30] , 
        \g5[6][29] , \g5[6][28] , \g5[6][27] , \g5[6][26] , \g5[6][25] , 
        \g5[6][24] , \g5[6][23] , \g5[6][22] , \g5[6][21] , \g5[6][20] , 
        \g5[6][19] , \g5[6][18] , \g5[6][17] , \g5[6][16] , \g5[6][15] , 
        \g5[6][14] , \g5[6][13] , \g5[6][12] , \g5[6][11] , \g5[6][10] , 
        \g5[6][9] , \g5[6][8] , \g5[6][7] , \g5[6][6] , \g5[6][5] , \g5[6][4] , 
        \g5[6][3] , \g5[6][2] , \g5[6][1] , 1'b0}), .b({\g5[7][63] , 
        \g5[7][62] , \g5[7][61] , \g5[7][60] , \g5[7][59] , \g5[7][58] , 
        \g5[7][57] , \g5[7][56] , \g5[7][55] , \g5[7][54] , \g5[7][53] , 
        \g5[7][52] , \g5[7][51] , \g5[7][50] , \g5[7][49] , \g5[7][48] , 
        \g5[7][47] , \g5[7][46] , \g5[7][45] , \g5[7][44] , \g5[7][43] , 
        \g5[7][42] , \g5[7][41] , \g5[7][40] , \g5[7][39] , \g5[7][38] , 
        \g5[7][37] , \g5[7][36] , \g5[7][35] , \g5[7][34] , \g5[7][33] , 
        \g5[7][32] , \g5[7][31] , \g5[7][30] , \g5[7][29] , \g5[7][28] , 
        \g5[7][27] , \g5[7][26] , \g5[7][25] , \g5[7][24] , \g5[7][23] , 
        \g5[7][22] , \g5[7][21] , \g5[7][20] , \g5[7][19] , \g5[7][18] , 
        \g5[7][17] , \g5[7][16] , \g5[7][15] , \g5[7][14] , \g5[7][13] , 
        \g5[7][12] , \g5[7][11] , \g5[7][10] , \g5[7][9] , \g5[7][8] , 
        \g5[7][7] , \g5[7][6] , \g5[7][5] , \g5[7][4] , \g5[7][3] , \g5[7][2] , 
        \g5[7][1] , 1'b0}), .cin({\g2[27][63] , \g2[27][62] , \g2[27][61] , 
        \g2[27][60] , \g2[27][59] , \g2[27][58] , \g2[27][57] , \g2[27][56] , 
        \g2[27][55] , \g2[27][54] , \g2[27][53] , \g2[27][52] , \g2[27][51] , 
        \g2[27][50] , \g2[27][49] , \g2[27][48] , \g2[27][47] , \g2[27][46] , 
        \g2[27][45] , \g2[27][44] , \g2[27][43] , \g2[27][42] , \g2[27][41] , 
        \g2[27][40] , \g2[27][39] , \g2[27][38] , \g2[27][37] , \g2[27][36] , 
        \g2[27][35] , \g2[27][34] , \g2[27][33] , \g2[27][32] , \g2[27][31] , 
        \g2[27][30] , \g2[27][29] , \g2[27][28] , \g2[27][27] , \g2[27][26] , 
        \g2[27][25] , \g2[27][24] , \g2[27][23] , \g2[27][22] , \g2[27][21] , 
        \g2[27][20] , \g2[27][19] , \g2[27][18] , \g2[27][17] , \g2[27][16] , 
        \g2[27][15] , \g2[27][14] , \g2[27][13] , \g2[27][12] , \g2[27][11] , 
        \g2[27][10] , \g2[27][9] , \g2[27][8] , \g2[27][7] , \g2[27][6] , 
        \g2[27][5] , \g2[27][4] , \g2[27][3] , \g2[27][2] , \g2[27][1] , 1'b0}), .sum({\g6[4][63] , \g6[4][62] , \g6[4][61] , \g6[4][60] , \g6[4][59] , 
        \g6[4][58] , \g6[4][57] , \g6[4][56] , \g6[4][55] , \g6[4][54] , 
        \g6[4][53] , \g6[4][52] , \g6[4][51] , \g6[4][50] , \g6[4][49] , 
        \g6[4][48] , \g6[4][47] , \g6[4][46] , \g6[4][45] , \g6[4][44] , 
        \g6[4][43] , \g6[4][42] , \g6[4][41] , \g6[4][40] , \g6[4][39] , 
        \g6[4][38] , \g6[4][37] , \g6[4][36] , \g6[4][35] , \g6[4][34] , 
        \g6[4][33] , \g6[4][32] , \g6[4][31] , \g6[4][30] , \g6[4][29] , 
        \g6[4][28] , \g6[4][27] , \g6[4][26] , \g6[4][25] , \g6[4][24] , 
        \g6[4][23] , \g6[4][22] , \g6[4][21] , \g6[4][20] , \g6[4][19] , 
        \g6[4][18] , \g6[4][17] , \g6[4][16] , \g6[4][15] , \g6[4][14] , 
        \g6[4][13] , \g6[4][12] , \g6[4][11] , \g6[4][10] , \g6[4][9] , 
        \g6[4][8] , \g6[4][7] , \g6[4][6] , \g6[4][5] , \g6[4][4] , \g6[4][3] , 
        \g6[4][2] , \g6[4][1] , \g6[4][0] }), .cout({\g6[5][63] , \g6[5][62] , 
        \g6[5][61] , \g6[5][60] , \g6[5][59] , \g6[5][58] , \g6[5][57] , 
        \g6[5][56] , \g6[5][55] , \g6[5][54] , \g6[5][53] , \g6[5][52] , 
        \g6[5][51] , \g6[5][50] , \g6[5][49] , \g6[5][48] , \g6[5][47] , 
        \g6[5][46] , \g6[5][45] , \g6[5][44] , \g6[5][43] , \g6[5][42] , 
        \g6[5][41] , \g6[5][40] , \g6[5][39] , \g6[5][38] , \g6[5][37] , 
        \g6[5][36] , \g6[5][35] , \g6[5][34] , \g6[5][33] , \g6[5][32] , 
        \g6[5][31] , \g6[5][30] , \g6[5][29] , \g6[5][28] , \g6[5][27] , 
        \g6[5][26] , \g6[5][25] , \g6[5][24] , \g6[5][23] , \g6[5][22] , 
        \g6[5][21] , \g6[5][20] , \g6[5][19] , \g6[5][18] , \g6[5][17] , 
        \g6[5][16] , \g6[5][15] , \g6[5][14] , \g6[5][13] , \g6[5][12] , 
        \g6[5][11] , \g6[5][10] , \g6[5][9] , \g6[5][8] , \g6[5][7] , 
        \g6[5][6] , \g6[5][5] , \g6[5][4] , \g6[5][3] , \g6[5][2] , \g6[5][1] , 
        SYNOPSYS_UNCONNECTED__56}) );
  FullAdder_5 F3 ( .a({\g6[0][63] , \g6[0][62] , \g6[0][61] , \g6[0][60] , 
        \g6[0][59] , \g6[0][58] , \g6[0][57] , \g6[0][56] , \g6[0][55] , 
        \g6[0][54] , \g6[0][53] , \g6[0][52] , \g6[0][51] , \g6[0][50] , 
        \g6[0][49] , \g6[0][48] , \g6[0][47] , \g6[0][46] , \g6[0][45] , 
        \g6[0][44] , \g6[0][43] , \g6[0][42] , \g6[0][41] , \g6[0][40] , 
        \g6[0][39] , \g6[0][38] , \g6[0][37] , \g6[0][36] , \g6[0][35] , 
        \g6[0][34] , \g6[0][33] , \g6[0][32] , \g6[0][31] , \g6[0][30] , 
        \g6[0][29] , \g6[0][28] , \g6[0][27] , \g6[0][26] , \g6[0][25] , 
        \g6[0][24] , \g6[0][23] , \g6[0][22] , \g6[0][21] , \g6[0][20] , 
        \g6[0][19] , \g6[0][18] , \g6[0][17] , \g6[0][16] , \g6[0][15] , 
        \g6[0][14] , \g6[0][13] , \g6[0][12] , \g6[0][11] , \g6[0][10] , 
        \g6[0][9] , \g6[0][8] , \g6[0][7] , \g6[0][6] , \g6[0][5] , \g6[0][4] , 
        \g6[0][3] , \g6[0][2] , \g6[0][1] , \g6[0][0] }), .b({\g6[1][63] , 
        \g6[1][62] , \g6[1][61] , \g6[1][60] , \g6[1][59] , \g6[1][58] , 
        \g6[1][57] , \g6[1][56] , \g6[1][55] , \g6[1][54] , \g6[1][53] , 
        \g6[1][52] , \g6[1][51] , \g6[1][50] , \g6[1][49] , \g6[1][48] , 
        \g6[1][47] , \g6[1][46] , \g6[1][45] , \g6[1][44] , \g6[1][43] , 
        \g6[1][42] , \g6[1][41] , \g6[1][40] , \g6[1][39] , \g6[1][38] , 
        \g6[1][37] , \g6[1][36] , \g6[1][35] , \g6[1][34] , \g6[1][33] , 
        \g6[1][32] , \g6[1][31] , \g6[1][30] , \g6[1][29] , \g6[1][28] , 
        \g6[1][27] , \g6[1][26] , \g6[1][25] , \g6[1][24] , \g6[1][23] , 
        \g6[1][22] , \g6[1][21] , \g6[1][20] , \g6[1][19] , \g6[1][18] , 
        \g6[1][17] , \g6[1][16] , \g6[1][15] , \g6[1][14] , \g6[1][13] , 
        \g6[1][12] , \g6[1][11] , \g6[1][10] , \g6[1][9] , \g6[1][8] , 
        \g6[1][7] , \g6[1][6] , \g6[1][5] , \g6[1][4] , \g6[1][3] , \g6[1][2] , 
        \g6[1][1] , 1'b0}), .cin({\g6[2][63] , \g6[2][62] , \g6[2][61] , 
        \g6[2][60] , \g6[2][59] , \g6[2][58] , \g6[2][57] , \g6[2][56] , 
        \g6[2][55] , \g6[2][54] , \g6[2][53] , \g6[2][52] , \g6[2][51] , 
        \g6[2][50] , \g6[2][49] , \g6[2][48] , \g6[2][47] , \g6[2][46] , 
        \g6[2][45] , \g6[2][44] , \g6[2][43] , \g6[2][42] , \g6[2][41] , 
        \g6[2][40] , \g6[2][39] , \g6[2][38] , \g6[2][37] , \g6[2][36] , 
        \g6[2][35] , \g6[2][34] , \g6[2][33] , \g6[2][32] , \g6[2][31] , 
        \g6[2][30] , \g6[2][29] , \g6[2][28] , \g6[2][27] , \g6[2][26] , 
        \g6[2][25] , \g6[2][24] , \g6[2][23] , \g6[2][22] , \g6[2][21] , 
        \g6[2][20] , \g6[2][19] , \g6[2][18] , \g6[2][17] , \g6[2][16] , 
        \g6[2][15] , \g6[2][14] , \g6[2][13] , \g6[2][12] , \g6[2][11] , 
        \g6[2][10] , \g6[2][9] , \g6[2][8] , \g6[2][7] , \g6[2][6] , 
        \g6[2][5] , \g6[2][4] , \g6[2][3] , \g6[2][2] , \g6[2][1] , \g6[2][0] }), .sum({\g7[0][63] , \g7[0][62] , \g7[0][61] , \g7[0][60] , \g7[0][59] , 
        \g7[0][58] , \g7[0][57] , \g7[0][56] , \g7[0][55] , \g7[0][54] , 
        \g7[0][53] , \g7[0][52] , \g7[0][51] , \g7[0][50] , \g7[0][49] , 
        \g7[0][48] , \g7[0][47] , \g7[0][46] , \g7[0][45] , \g7[0][44] , 
        \g7[0][43] , \g7[0][42] , \g7[0][41] , \g7[0][40] , \g7[0][39] , 
        \g7[0][38] , \g7[0][37] , \g7[0][36] , \g7[0][35] , \g7[0][34] , 
        \g7[0][33] , \g7[0][32] , \g7[0][31] , \g7[0][30] , \g7[0][29] , 
        \g7[0][28] , \g7[0][27] , \g7[0][26] , \g7[0][25] , \g7[0][24] , 
        \g7[0][23] , \g7[0][22] , \g7[0][21] , \g7[0][20] , \g7[0][19] , 
        \g7[0][18] , \g7[0][17] , \g7[0][16] , \g7[0][15] , \g7[0][14] , 
        \g7[0][13] , \g7[0][12] , \g7[0][11] , \g7[0][10] , \g7[0][9] , 
        \g7[0][8] , \g7[0][7] , \g7[0][6] , \g7[0][5] , \g7[0][4] , \g7[0][3] , 
        \g7[0][2] , \g7[0][1] , \g7[0][0] }), .cout({\g7[1][63] , \g7[1][62] , 
        \g7[1][61] , \g7[1][60] , \g7[1][59] , \g7[1][58] , \g7[1][57] , 
        \g7[1][56] , \g7[1][55] , \g7[1][54] , \g7[1][53] , \g7[1][52] , 
        \g7[1][51] , \g7[1][50] , \g7[1][49] , \g7[1][48] , \g7[1][47] , 
        \g7[1][46] , \g7[1][45] , \g7[1][44] , \g7[1][43] , \g7[1][42] , 
        \g7[1][41] , \g7[1][40] , \g7[1][39] , \g7[1][38] , \g7[1][37] , 
        \g7[1][36] , \g7[1][35] , \g7[1][34] , \g7[1][33] , \g7[1][32] , 
        \g7[1][31] , \g7[1][30] , \g7[1][29] , \g7[1][28] , \g7[1][27] , 
        \g7[1][26] , \g7[1][25] , \g7[1][24] , \g7[1][23] , \g7[1][22] , 
        \g7[1][21] , \g7[1][20] , \g7[1][19] , \g7[1][18] , \g7[1][17] , 
        \g7[1][16] , \g7[1][15] , \g7[1][14] , \g7[1][13] , \g7[1][12] , 
        \g7[1][11] , \g7[1][10] , \g7[1][9] , \g7[1][8] , \g7[1][7] , 
        \g7[1][6] , \g7[1][5] , \g7[1][4] , \g7[1][3] , \g7[1][2] , \g7[1][1] , 
        SYNOPSYS_UNCONNECTED__57}) );
  FullAdder_4 F4 ( .a({\g6[3][63] , \g6[3][62] , \g6[3][61] , \g6[3][60] , 
        \g6[3][59] , \g6[3][58] , \g6[3][57] , \g6[3][56] , \g6[3][55] , 
        \g6[3][54] , \g6[3][53] , \g6[3][52] , \g6[3][51] , \g6[3][50] , 
        \g6[3][49] , \g6[3][48] , \g6[3][47] , \g6[3][46] , \g6[3][45] , 
        \g6[3][44] , \g6[3][43] , \g6[3][42] , \g6[3][41] , \g6[3][40] , 
        \g6[3][39] , \g6[3][38] , \g6[3][37] , \g6[3][36] , \g6[3][35] , 
        \g6[3][34] , \g6[3][33] , \g6[3][32] , \g6[3][31] , \g6[3][30] , 
        \g6[3][29] , \g6[3][28] , \g6[3][27] , \g6[3][26] , \g6[3][25] , 
        \g6[3][24] , \g6[3][23] , \g6[3][22] , \g6[3][21] , \g6[3][20] , 
        \g6[3][19] , \g6[3][18] , \g6[3][17] , \g6[3][16] , \g6[3][15] , 
        \g6[3][14] , \g6[3][13] , \g6[3][12] , \g6[3][11] , \g6[3][10] , 
        \g6[3][9] , \g6[3][8] , \g6[3][7] , \g6[3][6] , \g6[3][5] , \g6[3][4] , 
        \g6[3][3] , \g6[3][2] , \g6[3][1] , 1'b0}), .b({\g6[4][63] , 
        \g6[4][62] , \g6[4][61] , \g6[4][60] , \g6[4][59] , \g6[4][58] , 
        \g6[4][57] , \g6[4][56] , \g6[4][55] , \g6[4][54] , \g6[4][53] , 
        \g6[4][52] , \g6[4][51] , \g6[4][50] , \g6[4][49] , \g6[4][48] , 
        \g6[4][47] , \g6[4][46] , \g6[4][45] , \g6[4][44] , \g6[4][43] , 
        \g6[4][42] , \g6[4][41] , \g6[4][40] , \g6[4][39] , \g6[4][38] , 
        \g6[4][37] , \g6[4][36] , \g6[4][35] , \g6[4][34] , \g6[4][33] , 
        \g6[4][32] , \g6[4][31] , \g6[4][30] , \g6[4][29] , \g6[4][28] , 
        \g6[4][27] , \g6[4][26] , \g6[4][25] , \g6[4][24] , \g6[4][23] , 
        \g6[4][22] , \g6[4][21] , \g6[4][20] , \g6[4][19] , \g6[4][18] , 
        \g6[4][17] , \g6[4][16] , \g6[4][15] , \g6[4][14] , \g6[4][13] , 
        \g6[4][12] , \g6[4][11] , \g6[4][10] , \g6[4][9] , \g6[4][8] , 
        \g6[4][7] , \g6[4][6] , \g6[4][5] , \g6[4][4] , \g6[4][3] , \g6[4][2] , 
        \g6[4][1] , \g6[4][0] }), .cin({\g6[5][63] , \g6[5][62] , \g6[5][61] , 
        \g6[5][60] , \g6[5][59] , \g6[5][58] , \g6[5][57] , \g6[5][56] , 
        \g6[5][55] , \g6[5][54] , \g6[5][53] , \g6[5][52] , \g6[5][51] , 
        \g6[5][50] , \g6[5][49] , \g6[5][48] , \g6[5][47] , \g6[5][46] , 
        \g6[5][45] , \g6[5][44] , \g6[5][43] , \g6[5][42] , \g6[5][41] , 
        \g6[5][40] , \g6[5][39] , \g6[5][38] , \g6[5][37] , \g6[5][36] , 
        \g6[5][35] , \g6[5][34] , \g6[5][33] , \g6[5][32] , \g6[5][31] , 
        \g6[5][30] , \g6[5][29] , \g6[5][28] , \g6[5][27] , \g6[5][26] , 
        \g6[5][25] , \g6[5][24] , \g6[5][23] , \g6[5][22] , \g6[5][21] , 
        \g6[5][20] , \g6[5][19] , \g6[5][18] , \g6[5][17] , \g6[5][16] , 
        \g6[5][15] , \g6[5][14] , \g6[5][13] , \g6[5][12] , \g6[5][11] , 
        \g6[5][10] , \g6[5][9] , \g6[5][8] , \g6[5][7] , \g6[5][6] , 
        \g6[5][5] , \g6[5][4] , \g6[5][3] , \g6[5][2] , \g6[5][1] , 1'b0}), 
        .sum({\g7[2][63] , \g7[2][62] , \g7[2][61] , \g7[2][60] , \g7[2][59] , 
        \g7[2][58] , \g7[2][57] , \g7[2][56] , \g7[2][55] , \g7[2][54] , 
        \g7[2][53] , \g7[2][52] , \g7[2][51] , \g7[2][50] , \g7[2][49] , 
        \g7[2][48] , \g7[2][47] , \g7[2][46] , \g7[2][45] , \g7[2][44] , 
        \g7[2][43] , \g7[2][42] , \g7[2][41] , \g7[2][40] , \g7[2][39] , 
        \g7[2][38] , \g7[2][37] , \g7[2][36] , \g7[2][35] , \g7[2][34] , 
        \g7[2][33] , \g7[2][32] , \g7[2][31] , \g7[2][30] , \g7[2][29] , 
        \g7[2][28] , \g7[2][27] , \g7[2][26] , \g7[2][25] , \g7[2][24] , 
        \g7[2][23] , \g7[2][22] , \g7[2][21] , \g7[2][20] , \g7[2][19] , 
        \g7[2][18] , \g7[2][17] , \g7[2][16] , \g7[2][15] , \g7[2][14] , 
        \g7[2][13] , \g7[2][12] , \g7[2][11] , \g7[2][10] , \g7[2][9] , 
        \g7[2][8] , \g7[2][7] , \g7[2][6] , \g7[2][5] , \g7[2][4] , \g7[2][3] , 
        \g7[2][2] , \g7[2][1] , \g7[2][0] }), .cout({\g7[3][63] , \g7[3][62] , 
        \g7[3][61] , \g7[3][60] , \g7[3][59] , \g7[3][58] , \g7[3][57] , 
        \g7[3][56] , \g7[3][55] , \g7[3][54] , \g7[3][53] , \g7[3][52] , 
        \g7[3][51] , \g7[3][50] , \g7[3][49] , \g7[3][48] , \g7[3][47] , 
        \g7[3][46] , \g7[3][45] , \g7[3][44] , \g7[3][43] , \g7[3][42] , 
        \g7[3][41] , \g7[3][40] , \g7[3][39] , \g7[3][38] , \g7[3][37] , 
        \g7[3][36] , \g7[3][35] , \g7[3][34] , \g7[3][33] , \g7[3][32] , 
        \g7[3][31] , \g7[3][30] , \g7[3][29] , \g7[3][28] , \g7[3][27] , 
        \g7[3][26] , \g7[3][25] , \g7[3][24] , \g7[3][23] , \g7[3][22] , 
        \g7[3][21] , \g7[3][20] , \g7[3][19] , \g7[3][18] , \g7[3][17] , 
        \g7[3][16] , \g7[3][15] , \g7[3][14] , \g7[3][13] , \g7[3][12] , 
        \g7[3][11] , \g7[3][10] , \g7[3][9] , \g7[3][8] , \g7[3][7] , 
        \g7[3][6] , \g7[3][5] , \g7[3][4] , \g7[3][3] , \g7[3][2] , \g7[3][1] , 
        SYNOPSYS_UNCONNECTED__58}) );
  FullAdder_3 F5 ( .a({\g7[0][63] , \g7[0][62] , \g7[0][61] , \g7[0][60] , 
        \g7[0][59] , \g7[0][58] , \g7[0][57] , \g7[0][56] , \g7[0][55] , 
        \g7[0][54] , \g7[0][53] , \g7[0][52] , \g7[0][51] , \g7[0][50] , 
        \g7[0][49] , \g7[0][48] , \g7[0][47] , \g7[0][46] , \g7[0][45] , 
        \g7[0][44] , \g7[0][43] , \g7[0][42] , \g7[0][41] , \g7[0][40] , 
        \g7[0][39] , \g7[0][38] , \g7[0][37] , \g7[0][36] , \g7[0][35] , 
        \g7[0][34] , \g7[0][33] , \g7[0][32] , \g7[0][31] , \g7[0][30] , 
        \g7[0][29] , \g7[0][28] , \g7[0][27] , \g7[0][26] , \g7[0][25] , 
        \g7[0][24] , \g7[0][23] , \g7[0][22] , \g7[0][21] , \g7[0][20] , 
        \g7[0][19] , \g7[0][18] , \g7[0][17] , \g7[0][16] , \g7[0][15] , 
        \g7[0][14] , \g7[0][13] , \g7[0][12] , \g7[0][11] , \g7[0][10] , 
        \g7[0][9] , \g7[0][8] , \g7[0][7] , \g7[0][6] , \g7[0][5] , \g7[0][4] , 
        \g7[0][3] , \g7[0][2] , \g7[0][1] , \g7[0][0] }), .b({\g7[1][63] , 
        \g7[1][62] , \g7[1][61] , \g7[1][60] , \g7[1][59] , \g7[1][58] , 
        \g7[1][57] , \g7[1][56] , \g7[1][55] , \g7[1][54] , \g7[1][53] , 
        \g7[1][52] , \g7[1][51] , \g7[1][50] , \g7[1][49] , \g7[1][48] , 
        \g7[1][47] , \g7[1][46] , \g7[1][45] , \g7[1][44] , \g7[1][43] , 
        \g7[1][42] , \g7[1][41] , \g7[1][40] , \g7[1][39] , \g7[1][38] , 
        \g7[1][37] , \g7[1][36] , \g7[1][35] , \g7[1][34] , \g7[1][33] , 
        \g7[1][32] , \g7[1][31] , \g7[1][30] , \g7[1][29] , \g7[1][28] , 
        \g7[1][27] , \g7[1][26] , \g7[1][25] , \g7[1][24] , \g7[1][23] , 
        \g7[1][22] , \g7[1][21] , \g7[1][20] , \g7[1][19] , \g7[1][18] , 
        \g7[1][17] , \g7[1][16] , \g7[1][15] , \g7[1][14] , \g7[1][13] , 
        \g7[1][12] , \g7[1][11] , \g7[1][10] , \g7[1][9] , \g7[1][8] , 
        \g7[1][7] , \g7[1][6] , \g7[1][5] , \g7[1][4] , \g7[1][3] , \g7[1][2] , 
        \g7[1][1] , 1'b0}), .cin({\g7[2][63] , \g7[2][62] , \g7[2][61] , 
        \g7[2][60] , \g7[2][59] , \g7[2][58] , \g7[2][57] , \g7[2][56] , 
        \g7[2][55] , \g7[2][54] , \g7[2][53] , \g7[2][52] , \g7[2][51] , 
        \g7[2][50] , \g7[2][49] , \g7[2][48] , \g7[2][47] , \g7[2][46] , 
        \g7[2][45] , \g7[2][44] , \g7[2][43] , \g7[2][42] , \g7[2][41] , 
        \g7[2][40] , \g7[2][39] , \g7[2][38] , \g7[2][37] , \g7[2][36] , 
        \g7[2][35] , \g7[2][34] , \g7[2][33] , \g7[2][32] , \g7[2][31] , 
        \g7[2][30] , \g7[2][29] , \g7[2][28] , \g7[2][27] , \g7[2][26] , 
        \g7[2][25] , \g7[2][24] , \g7[2][23] , \g7[2][22] , \g7[2][21] , 
        \g7[2][20] , \g7[2][19] , \g7[2][18] , \g7[2][17] , \g7[2][16] , 
        \g7[2][15] , \g7[2][14] , \g7[2][13] , \g7[2][12] , \g7[2][11] , 
        \g7[2][10] , \g7[2][9] , \g7[2][8] , \g7[2][7] , \g7[2][6] , 
        \g7[2][5] , \g7[2][4] , \g7[2][3] , \g7[2][2] , \g7[2][1] , \g7[2][0] }), .sum({\g8[0][63] , \g8[0][62] , \g8[0][61] , \g8[0][60] , \g8[0][59] , 
        \g8[0][58] , \g8[0][57] , \g8[0][56] , \g8[0][55] , \g8[0][54] , 
        \g8[0][53] , \g8[0][52] , \g8[0][51] , \g8[0][50] , \g8[0][49] , 
        \g8[0][48] , \g8[0][47] , \g8[0][46] , \g8[0][45] , \g8[0][44] , 
        \g8[0][43] , \g8[0][42] , \g8[0][41] , \g8[0][40] , \g8[0][39] , 
        \g8[0][38] , \g8[0][37] , \g8[0][36] , \g8[0][35] , \g8[0][34] , 
        \g8[0][33] , \g8[0][32] , \g8[0][31] , \g8[0][30] , \g8[0][29] , 
        \g8[0][28] , \g8[0][27] , \g8[0][26] , \g8[0][25] , \g8[0][24] , 
        \g8[0][23] , \g8[0][22] , \g8[0][21] , \g8[0][20] , \g8[0][19] , 
        \g8[0][18] , \g8[0][17] , \g8[0][16] , \g8[0][15] , \g8[0][14] , 
        \g8[0][13] , \g8[0][12] , \g8[0][11] , \g8[0][10] , \g8[0][9] , 
        \g8[0][8] , \g8[0][7] , \g8[0][6] , \g8[0][5] , \g8[0][4] , \g8[0][3] , 
        \g8[0][2] , \g8[0][1] , \g8[0][0] }), .cout({\g8[1][63] , \g8[1][62] , 
        \g8[1][61] , \g8[1][60] , \g8[1][59] , \g8[1][58] , \g8[1][57] , 
        \g8[1][56] , \g8[1][55] , \g8[1][54] , \g8[1][53] , \g8[1][52] , 
        \g8[1][51] , \g8[1][50] , \g8[1][49] , \g8[1][48] , \g8[1][47] , 
        \g8[1][46] , \g8[1][45] , \g8[1][44] , \g8[1][43] , \g8[1][42] , 
        \g8[1][41] , \g8[1][40] , \g8[1][39] , \g8[1][38] , \g8[1][37] , 
        \g8[1][36] , \g8[1][35] , \g8[1][34] , \g8[1][33] , \g8[1][32] , 
        \g8[1][31] , \g8[1][30] , \g8[1][29] , \g8[1][28] , \g8[1][27] , 
        \g8[1][26] , \g8[1][25] , \g8[1][24] , \g8[1][23] , \g8[1][22] , 
        \g8[1][21] , \g8[1][20] , \g8[1][19] , \g8[1][18] , \g8[1][17] , 
        \g8[1][16] , \g8[1][15] , \g8[1][14] , \g8[1][13] , \g8[1][12] , 
        \g8[1][11] , \g8[1][10] , \g8[1][9] , \g8[1][8] , \g8[1][7] , 
        \g8[1][6] , \g8[1][5] , \g8[1][4] , \g8[1][3] , \g8[1][2] , \g8[1][1] , 
        SYNOPSYS_UNCONNECTED__59}) );
  FullAdder_2 F6 ( .a({\g8[0][63] , \g8[0][62] , \g8[0][61] , \g8[0][60] , 
        \g8[0][59] , \g8[0][58] , \g8[0][57] , \g8[0][56] , \g8[0][55] , 
        \g8[0][54] , \g8[0][53] , \g8[0][52] , \g8[0][51] , \g8[0][50] , 
        \g8[0][49] , \g8[0][48] , \g8[0][47] , \g8[0][46] , \g8[0][45] , 
        \g8[0][44] , \g8[0][43] , \g8[0][42] , \g8[0][41] , \g8[0][40] , 
        \g8[0][39] , \g8[0][38] , \g8[0][37] , \g8[0][36] , \g8[0][35] , 
        \g8[0][34] , \g8[0][33] , \g8[0][32] , \g8[0][31] , \g8[0][30] , 
        \g8[0][29] , \g8[0][28] , \g8[0][27] , \g8[0][26] , \g8[0][25] , 
        \g8[0][24] , \g8[0][23] , \g8[0][22] , \g8[0][21] , \g8[0][20] , 
        \g8[0][19] , \g8[0][18] , \g8[0][17] , \g8[0][16] , \g8[0][15] , 
        \g8[0][14] , \g8[0][13] , \g8[0][12] , \g8[0][11] , \g8[0][10] , 
        \g8[0][9] , \g8[0][8] , \g8[0][7] , \g8[0][6] , \g8[0][5] , \g8[0][4] , 
        \g8[0][3] , \g8[0][2] , \g8[0][1] , \g8[0][0] }), .b({\g8[1][63] , 
        \g8[1][62] , \g8[1][61] , \g8[1][60] , \g8[1][59] , \g8[1][58] , 
        \g8[1][57] , \g8[1][56] , \g8[1][55] , \g8[1][54] , \g8[1][53] , 
        \g8[1][52] , \g8[1][51] , \g8[1][50] , \g8[1][49] , \g8[1][48] , 
        \g8[1][47] , \g8[1][46] , \g8[1][45] , \g8[1][44] , \g8[1][43] , 
        \g8[1][42] , \g8[1][41] , \g8[1][40] , \g8[1][39] , \g8[1][38] , 
        \g8[1][37] , \g8[1][36] , \g8[1][35] , \g8[1][34] , \g8[1][33] , 
        \g8[1][32] , \g8[1][31] , \g8[1][30] , \g8[1][29] , \g8[1][28] , 
        \g8[1][27] , \g8[1][26] , \g8[1][25] , \g8[1][24] , \g8[1][23] , 
        \g8[1][22] , \g8[1][21] , \g8[1][20] , \g8[1][19] , \g8[1][18] , 
        \g8[1][17] , \g8[1][16] , \g8[1][15] , \g8[1][14] , \g8[1][13] , 
        \g8[1][12] , \g8[1][11] , \g8[1][10] , \g8[1][9] , \g8[1][8] , 
        \g8[1][7] , \g8[1][6] , \g8[1][5] , \g8[1][4] , \g8[1][3] , \g8[1][2] , 
        \g8[1][1] , 1'b0}), .cin({\g7[3][63] , \g7[3][62] , \g7[3][61] , 
        \g7[3][60] , \g7[3][59] , \g7[3][58] , \g7[3][57] , \g7[3][56] , 
        \g7[3][55] , \g7[3][54] , \g7[3][53] , \g7[3][52] , \g7[3][51] , 
        \g7[3][50] , \g7[3][49] , \g7[3][48] , \g7[3][47] , \g7[3][46] , 
        \g7[3][45] , \g7[3][44] , \g7[3][43] , \g7[3][42] , \g7[3][41] , 
        \g7[3][40] , \g7[3][39] , \g7[3][38] , \g7[3][37] , \g7[3][36] , 
        \g7[3][35] , \g7[3][34] , \g7[3][33] , \g7[3][32] , \g7[3][31] , 
        \g7[3][30] , \g7[3][29] , \g7[3][28] , \g7[3][27] , \g7[3][26] , 
        \g7[3][25] , \g7[3][24] , \g7[3][23] , \g7[3][22] , \g7[3][21] , 
        \g7[3][20] , \g7[3][19] , \g7[3][18] , \g7[3][17] , \g7[3][16] , 
        \g7[3][15] , \g7[3][14] , \g7[3][13] , \g7[3][12] , \g7[3][11] , 
        \g7[3][10] , \g7[3][9] , \g7[3][8] , \g7[3][7] , \g7[3][6] , 
        \g7[3][5] , \g7[3][4] , \g7[3][3] , \g7[3][2] , \g7[3][1] , 1'b0}), 
        .sum({\g9[0][63] , \g9[0][62] , \g9[0][61] , \g9[0][60] , \g9[0][59] , 
        \g9[0][58] , \g9[0][57] , \g9[0][56] , \g9[0][55] , \g9[0][54] , 
        \g9[0][53] , \g9[0][52] , \g9[0][51] , \g9[0][50] , \g9[0][49] , 
        \g9[0][48] , \g9[0][47] , \g9[0][46] , \g9[0][45] , \g9[0][44] , 
        \g9[0][43] , \g9[0][42] , \g9[0][41] , \g9[0][40] , \g9[0][39] , 
        \g9[0][38] , \g9[0][37] , \g9[0][36] , \g9[0][35] , \g9[0][34] , 
        \g9[0][33] , \g9[0][32] , \g9[0][31] , \g9[0][30] , \g9[0][29] , 
        \g9[0][28] , \g9[0][27] , \g9[0][26] , \g9[0][25] , \g9[0][24] , 
        \g9[0][23] , \g9[0][22] , \g9[0][21] , \g9[0][20] , \g9[0][19] , 
        \g9[0][18] , \g9[0][17] , \g9[0][16] , \g9[0][15] , \g9[0][14] , 
        \g9[0][13] , \g9[0][12] , \g9[0][11] , \g9[0][10] , \g9[0][9] , 
        \g9[0][8] , \g9[0][7] , \g9[0][6] , \g9[0][5] , \g9[0][4] , \g9[0][3] , 
        \g9[0][2] , \g9[0][1] , \g9[0][0] }), .cout({\g9[1][63] , \g9[1][62] , 
        \g9[1][61] , \g9[1][60] , \g9[1][59] , \g9[1][58] , \g9[1][57] , 
        \g9[1][56] , \g9[1][55] , \g9[1][54] , \g9[1][53] , \g9[1][52] , 
        \g9[1][51] , \g9[1][50] , \g9[1][49] , \g9[1][48] , \g9[1][47] , 
        \g9[1][46] , \g9[1][45] , \g9[1][44] , \g9[1][43] , \g9[1][42] , 
        \g9[1][41] , \g9[1][40] , \g9[1][39] , \g9[1][38] , \g9[1][37] , 
        \g9[1][36] , \g9[1][35] , \g9[1][34] , \g9[1][33] , \g9[1][32] , 
        \g9[1][31] , \g9[1][30] , \g9[1][29] , \g9[1][28] , \g9[1][27] , 
        \g9[1][26] , \g9[1][25] , \g9[1][24] , \g9[1][23] , \g9[1][22] , 
        \g9[1][21] , \g9[1][20] , \g9[1][19] , \g9[1][18] , \g9[1][17] , 
        \g9[1][16] , \g9[1][15] , \g9[1][14] , \g9[1][13] , \g9[1][12] , 
        \g9[1][11] , \g9[1][10] , \g9[1][9] , \g9[1][8] , \g9[1][7] , 
        \g9[1][6] , \g9[1][5] , \g9[1][4] , \g9[1][3] , \g9[1][2] , \g9[1][1] , 
        SYNOPSYS_UNCONNECTED__60}) );
  FullAdder_1 F7 ( .a({\g9[0][63] , \g9[0][62] , \g9[0][61] , \g9[0][60] , 
        \g9[0][59] , \g9[0][58] , \g9[0][57] , \g9[0][56] , \g9[0][55] , 
        \g9[0][54] , \g9[0][53] , \g9[0][52] , \g9[0][51] , \g9[0][50] , 
        \g9[0][49] , \g9[0][48] , \g9[0][47] , \g9[0][46] , \g9[0][45] , 
        \g9[0][44] , \g9[0][43] , \g9[0][42] , \g9[0][41] , \g9[0][40] , 
        \g9[0][39] , \g9[0][38] , \g9[0][37] , \g9[0][36] , \g9[0][35] , 
        \g9[0][34] , \g9[0][33] , \g9[0][32] , \g9[0][31] , \g9[0][30] , 
        \g9[0][29] , \g9[0][28] , \g9[0][27] , \g9[0][26] , \g9[0][25] , 
        \g9[0][24] , \g9[0][23] , \g9[0][22] , \g9[0][21] , \g9[0][20] , 
        \g9[0][19] , \g9[0][18] , \g9[0][17] , \g9[0][16] , \g9[0][15] , 
        \g9[0][14] , \g9[0][13] , \g9[0][12] , \g9[0][11] , \g9[0][10] , 
        \g9[0][9] , \g9[0][8] , \g9[0][7] , \g9[0][6] , \g9[0][5] , \g9[0][4] , 
        \g9[0][3] , \g9[0][2] , \g9[0][1] , \g9[0][0] }), .b({\g9[1][63] , 
        \g9[1][62] , \g9[1][61] , \g9[1][60] , \g9[1][59] , \g9[1][58] , 
        \g9[1][57] , \g9[1][56] , \g9[1][55] , \g9[1][54] , \g9[1][53] , 
        \g9[1][52] , \g9[1][51] , \g9[1][50] , \g9[1][49] , \g9[1][48] , 
        \g9[1][47] , \g9[1][46] , \g9[1][45] , \g9[1][44] , \g9[1][43] , 
        \g9[1][42] , \g9[1][41] , \g9[1][40] , \g9[1][39] , \g9[1][38] , 
        \g9[1][37] , \g9[1][36] , \g9[1][35] , \g9[1][34] , \g9[1][33] , 
        \g9[1][32] , \g9[1][31] , \g9[1][30] , \g9[1][29] , \g9[1][28] , 
        \g9[1][27] , \g9[1][26] , \g9[1][25] , \g9[1][24] , \g9[1][23] , 
        \g9[1][22] , \g9[1][21] , \g9[1][20] , \g9[1][19] , \g9[1][18] , 
        \g9[1][17] , \g9[1][16] , \g9[1][15] , \g9[1][14] , \g9[1][13] , 
        \g9[1][12] , \g9[1][11] , \g9[1][10] , \g9[1][9] , \g9[1][8] , 
        \g9[1][7] , \g9[1][6] , \g9[1][5] , \g9[1][4] , \g9[1][3] , \g9[1][2] , 
        \g9[1][1] , 1'b0}), .cin({n499, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sum({
        \g10[0][63] , \g10[0][62] , \g10[0][61] , \g10[0][60] , \g10[0][59] , 
        \g10[0][58] , \g10[0][57] , \g10[0][56] , \g10[0][55] , \g10[0][54] , 
        \g10[0][53] , \g10[0][52] , \g10[0][51] , \g10[0][50] , \g10[0][49] , 
        \g10[0][48] , \g10[0][47] , \g10[0][46] , \g10[0][45] , \g10[0][44] , 
        \g10[0][43] , \g10[0][42] , \g10[0][41] , \g10[0][40] , \g10[0][39] , 
        \g10[0][38] , \g10[0][37] , \g10[0][36] , \g10[0][35] , \g10[0][34] , 
        \g10[0][33] , \g10[0][32] , \g10[0][31] , \g10[0][30] , \g10[0][29] , 
        \g10[0][28] , \g10[0][27] , \g10[0][26] , \g10[0][25] , \g10[0][24] , 
        \g10[0][23] , \g10[0][22] , \g10[0][21] , \g10[0][20] , \g10[0][19] , 
        \g10[0][18] , \g10[0][17] , \g10[0][16] , \g10[0][15] , \g10[0][14] , 
        \g10[0][13] , \g10[0][12] , \g10[0][11] , \g10[0][10] , \g10[0][9] , 
        \g10[0][8] , \g10[0][7] , \g10[0][6] , \g10[0][5] , \g10[0][4] , 
        \g10[0][3] , \g10[0][2] , \g10[0][1] , \g10[0][0] }), .cout({
        \g10[1][63] , \g10[1][62] , \g10[1][61] , \g10[1][60] , \g10[1][59] , 
        \g10[1][58] , \g10[1][57] , \g10[1][56] , \g10[1][55] , \g10[1][54] , 
        \g10[1][53] , \g10[1][52] , \g10[1][51] , \g10[1][50] , \g10[1][49] , 
        \g10[1][48] , \g10[1][47] , \g10[1][46] , \g10[1][45] , \g10[1][44] , 
        \g10[1][43] , \g10[1][42] , \g10[1][41] , \g10[1][40] , \g10[1][39] , 
        \g10[1][38] , \g10[1][37] , \g10[1][36] , \g10[1][35] , \g10[1][34] , 
        \g10[1][33] , \g10[1][32] , \g10[1][31] , \g10[1][30] , \g10[1][29] , 
        \g10[1][28] , \g10[1][27] , \g10[1][26] , \g10[1][25] , \g10[1][24] , 
        \g10[1][23] , \g10[1][22] , \g10[1][21] , \g10[1][20] , \g10[1][19] , 
        \g10[1][18] , \g10[1][17] , \g10[1][16] , \g10[1][15] , \g10[1][14] , 
        \g10[1][13] , \g10[1][12] , \g10[1][11] , \g10[1][10] , \g10[1][9] , 
        \g10[1][8] , \g10[1][7] , \g10[1][6] , \g10[1][5] , \g10[1][4] , 
        \g10[1][3] , \g10[1][2] , \g10[1][1] , SYNOPSYS_UNCONNECTED__61}) );
  WallaceTreeMultiplier_DW01_add_0 add_110 ( .A({\g10[1][63] , \g10[1][62] , 
        \g10[1][61] , \g10[1][60] , \g10[1][59] , \g10[1][58] , \g10[1][57] , 
        \g10[1][56] , \g10[1][55] , \g10[1][54] , \g10[1][53] , \g10[1][52] , 
        \g10[1][51] , \g10[1][50] , \g10[1][49] , \g10[1][48] , \g10[1][47] , 
        \g10[1][46] , \g10[1][45] , \g10[1][44] , \g10[1][43] , \g10[1][42] , 
        \g10[1][41] , \g10[1][40] , \g10[1][39] , \g10[1][38] , \g10[1][37] , 
        \g10[1][36] , \g10[1][35] , \g10[1][34] , \g10[1][33] , \g10[1][32] , 
        \g10[1][31] , \g10[1][30] , \g10[1][29] , \g10[1][28] , \g10[1][27] , 
        \g10[1][26] , \g10[1][25] , \g10[1][24] , \g10[1][23] , \g10[1][22] , 
        \g10[1][21] , \g10[1][20] , \g10[1][19] , \g10[1][18] , \g10[1][17] , 
        \g10[1][16] , \g10[1][15] , \g10[1][14] , \g10[1][13] , \g10[1][12] , 
        \g10[1][11] , \g10[1][10] , \g10[1][9] , \g10[1][8] , \g10[1][7] , 
        \g10[1][6] , \g10[1][5] , \g10[1][4] , \g10[1][3] , \g10[1][2] , 
        \g10[1][1] , 1'b0}), .B({\g10[0][63] , \g10[0][62] , \g10[0][61] , 
        \g10[0][60] , \g10[0][59] , \g10[0][58] , \g10[0][57] , \g10[0][56] , 
        \g10[0][55] , \g10[0][54] , \g10[0][53] , \g10[0][52] , \g10[0][51] , 
        \g10[0][50] , \g10[0][49] , \g10[0][48] , \g10[0][47] , \g10[0][46] , 
        \g10[0][45] , \g10[0][44] , \g10[0][43] , \g10[0][42] , \g10[0][41] , 
        \g10[0][40] , \g10[0][39] , \g10[0][38] , \g10[0][37] , \g10[0][36] , 
        \g10[0][35] , \g10[0][34] , \g10[0][33] , \g10[0][32] , \g10[0][31] , 
        \g10[0][30] , \g10[0][29] , \g10[0][28] , \g10[0][27] , \g10[0][26] , 
        \g10[0][25] , \g10[0][24] , \g10[0][23] , \g10[0][22] , \g10[0][21] , 
        \g10[0][20] , \g10[0][19] , \g10[0][18] , \g10[0][17] , \g10[0][16] , 
        \g10[0][15] , \g10[0][14] , \g10[0][13] , \g10[0][12] , \g10[0][11] , 
        \g10[0][10] , \g10[0][9] , \g10[0][8] , \g10[0][7] , \g10[0][6] , 
        \g10[0][5] , \g10[0][4] , \g10[0][3] , \g10[0][2] , \g10[0][1] , 
        \g10[0][0] }), .CI(1'b0), .SUM({N194, N193, N192, N191, N190, N189, 
        N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, 
        N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, 
        N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, 
        N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, 
        N140, N139, N138, N137, N136, N135, N134, N133, N132, N131}) );
  DFFX1 \B_reg_reg[0]  ( .D(N67), .CLK(clk), .Q(B_reg[0]), .QN(n142) );
  DFFX1 \B_reg_reg[1]  ( .D(N68), .CLK(clk), .Q(B_reg[1]), .QN(n141) );
  DFFX2 \A_reg_reg[10]  ( .D(N45), .CLK(clk), .Q(A_reg[10]), .QN(n121) );
  DFFX1 \B_reg_reg[4]  ( .D(N71), .CLK(clk), .Q(B_reg[4]), .QN(n143) );
  DFFX1 \B_reg_reg[3]  ( .D(N70), .CLK(clk), .Q(B_reg[3]), .QN(n145) );
  DFFX1 \B_reg_reg[2]  ( .D(N69), .CLK(clk), .Q(B_reg[2]), .QN(n136) );
  DELLN1X2 U1219 ( .INP(n552), .Z(n274) );
  AND2X4 U1220 ( .IN1(A_reg[3]), .IN2(B_reg[1]), .Q(\p[1][4] ) );
  AND2X4 U1221 ( .IN1(A_reg[3]), .IN2(B_reg[4]), .Q(\p[4][7] ) );
  DELLN2X2 U1222 ( .INP(n560), .Z(n132) );
  DELLN2X2 U1223 ( .INP(n560), .Z(n131) );
  DELLN2X2 U1224 ( .INP(n560), .Z(n355) );
  DELLN2X2 U1225 ( .INP(n555), .Z(n285) );
  DELLN2X2 U1226 ( .INP(n555), .Z(n283) );
  DELLN1X2 U1227 ( .INP(n561), .Z(n117) );
  DELLN1X2 U1228 ( .INP(n561), .Z(n358) );
  DELLN1X2 U1229 ( .INP(n559), .Z(n124) );
  DELLN2X2 U1230 ( .INP(n559), .Z(n354) );
  DELLN1X2 U1231 ( .INP(n559), .Z(n353) );
  DELLN2X2 U1232 ( .INP(n559), .Z(n352) );
  INVX0 U1233 ( .INP(n128), .ZN(n66) );
  DELLN2X2 U1234 ( .INP(n129), .Z(n127) );
  DELLN2X2 U1235 ( .INP(n129), .Z(n343) );
  DELLN2X2 U1236 ( .INP(n547), .Z(n254) );
  DELLN2X2 U1237 ( .INP(n547), .Z(n256) );
  DELLN2X2 U1238 ( .INP(n547), .Z(n257) );
  INVX0 U1239 ( .INP(B_reg[1]), .ZN(n67) );
  INVX0 U1240 ( .INP(B_reg[1]), .ZN(n68) );
  DELLN1X2 U1241 ( .INP(n563), .Z(n368) );
  DELLN2X2 U1242 ( .INP(n553), .Z(n279) );
  DELLN2X2 U1243 ( .INP(n552), .Z(n276) );
  DELLN2X2 U1244 ( .INP(n552), .Z(n275) );
  DELLN2X2 U1245 ( .INP(n548), .Z(n263) );
  DELLN2X2 U1246 ( .INP(n548), .Z(n150) );
  DELLN2X2 U1247 ( .INP(n548), .Z(n261) );
  DELLN2X2 U1248 ( .INP(n548), .Z(n262) );
  DELLN1X2 U1249 ( .INP(n548), .Z(n151) );
  DELLN2X2 U1250 ( .INP(n72), .Z(n344) );
  NBUFFX2 U1251 ( .INP(n71), .Z(n346) );
  NBUFFX4 U1252 ( .INP(n108), .Z(n334) );
  NBUFFX4 U1253 ( .INP(n562), .Z(n134) );
  NBUFFX4 U1254 ( .INP(n562), .Z(n364) );
  DELLN1X2 U1255 ( .INP(n108), .Z(n336) );
  DELLN1X2 U1256 ( .INP(n111), .Z(n340) );
  NBUFFX4 U1257 ( .INP(n111), .Z(n341) );
  NBUFFX4 U1258 ( .INP(n145), .Z(n362) );
  NBUFFX4 U1259 ( .INP(n112), .Z(n258) );
  DELLN1X2 U1260 ( .INP(n110), .Z(n246) );
  DELLN1X2 U1261 ( .INP(n129), .Z(n128) );
  DELLN1X2 U1262 ( .INP(n110), .Z(n249) );
  DELLN1X2 U1263 ( .INP(n107), .Z(n333) );
  NBUFFX4 U1264 ( .INP(n118), .Z(n245) );
  DELLN1X2 U1265 ( .INP(n110), .Z(n248) );
  DELLN1X2 U1266 ( .INP(n116), .Z(n338) );
  DELLN1X2 U1267 ( .INP(n107), .Z(n331) );
  AND2X1 U1268 ( .IN1(A_reg[2]), .IN2(B_reg[3]), .Q(\p[3][5] ) );
  AND2X1 U1269 ( .IN1(A_reg[2]), .IN2(B_reg[2]), .Q(\p[2][4] ) );
  AND2X1 U1270 ( .IN1(B_reg[3]), .IN2(A_reg[1]), .Q(\p[3][4] ) );
  AND2X1 U1271 ( .IN1(A_reg[6]), .IN2(B_reg[1]), .Q(\p[1][7] ) );
  AND2X1 U1272 ( .IN1(A_reg[6]), .IN2(B_reg[3]), .Q(\p[3][9] ) );
  AND2X1 U1273 ( .IN1(A_reg[5]), .IN2(B_reg[4]), .Q(\p[4][9] ) );
  AND2X1 U1274 ( .IN1(A_reg[10]), .IN2(B_reg[1]), .Q(\p[1][11] ) );
  AND2X1 U1275 ( .IN1(n540), .IN2(A_reg[11]), .Q(\p[52][63] ) );
  INVX0 U1276 ( .INP(n139), .ZN(n69) );
  INVX0 U1277 ( .INP(n69), .ZN(n70) );
  INVX0 U1278 ( .INP(n69), .ZN(n71) );
  INVX0 U1279 ( .INP(n69), .ZN(n72) );
  DELLN1X2 U1280 ( .INP(n81), .Z(n319) );
  INVX0 U1281 ( .INP(B_reg[4]), .ZN(n105) );
  AND2X4 U1282 ( .IN1(n540), .IN2(A_reg[3]), .Q(\p[60][63] ) );
  AND2X4 U1283 ( .IN1(B_reg[3]), .IN2(n545), .Q(\p[3][63] ) );
  NBUFFX4 U1284 ( .INP(n80), .Z(n226) );
  NBUFFX4 U1285 ( .INP(n80), .Z(n227) );
  NBUFFX4 U1286 ( .INP(n80), .Z(n228) );
  DELLN1X2 U1287 ( .INP(n562), .Z(n365) );
  DELLN1X2 U1288 ( .INP(n550), .Z(n269) );
  DELLN1X2 U1289 ( .INP(n560), .Z(n356) );
  DELLN1X2 U1290 ( .INP(n88), .Z(n234) );
  DELLN1X2 U1291 ( .INP(n88), .Z(n235) );
  INVX0 U1292 ( .INP(A_reg[1]), .ZN(n106) );
  DELLN1X2 U1293 ( .INP(n554), .Z(n280) );
  DELLN1X2 U1294 ( .INP(n554), .Z(n281) );
  DELLN1X2 U1295 ( .INP(n107), .Z(n332) );
  DELLN1X2 U1296 ( .INP(n108), .Z(n335) );
  INVX0 U1297 ( .INP(B_reg[3]), .ZN(n109) );
  DELLN1X2 U1298 ( .INP(n105), .Z(n360) );
  AND2X4 U1299 ( .IN1(n540), .IN2(A_reg[1]), .Q(\p[62][63] ) );
  DELLN1X2 U1300 ( .INP(n118), .Z(n243) );
  DELLN1X2 U1301 ( .INP(n118), .Z(n242) );
  AND2X4 U1302 ( .IN1(B_reg[0]), .IN2(n543), .Q(\p[0][63] ) );
  AND2X4 U1303 ( .IN1(B_reg[2]), .IN2(n544), .Q(\p[2][63] ) );
  DELLN1X2 U1304 ( .INP(n563), .Z(n367) );
  DELLN1X2 U1305 ( .INP(n563), .Z(n366) );
  AND2X1 U1306 ( .IN1(A_reg[7]), .IN2(B_reg[5]), .Q(\p[5][12] ) );
  DELLN1X2 U1307 ( .INP(n110), .Z(n247) );
  DELLN1X2 U1308 ( .INP(n82), .Z(n328) );
  AND2X4 U1309 ( .IN1(A_reg[5]), .IN2(B_reg[1]), .Q(\p[1][6] ) );
  DELLN1X2 U1310 ( .INP(n89), .Z(n241) );
  DELLN1X2 U1311 ( .INP(n89), .Z(n239) );
  DELLN1X2 U1312 ( .INP(n89), .Z(n238) );
  INVX0 U1313 ( .INP(A_reg[8]), .ZN(n112) );
  DELLN1X2 U1314 ( .INP(n149), .Z(n114) );
  AND2X2 U1315 ( .IN1(n540), .IN2(A_reg[4]), .Q(\p[59][63] ) );
  DELLN1X2 U1316 ( .INP(n551), .Z(n273) );
  DELLN1X2 U1317 ( .INP(n116), .Z(n337) );
  NBUFFX2 U1318 ( .INP(n74), .Z(n208) );
  NBUFFX2 U1319 ( .INP(\p[61][63] ), .Z(n491) );
  NBUFFX2 U1320 ( .INP(n91), .Z(n292) );
  DELLN1X2 U1321 ( .INP(n100), .Z(n305) );
  DELLN1X2 U1322 ( .INP(n102), .Z(n302) );
  DELLN1X2 U1323 ( .INP(n101), .Z(n299) );
  DELLN1X2 U1324 ( .INP(n143), .Z(n359) );
  DELLN1X2 U1325 ( .INP(n564), .Z(n371) );
  DELLN1X2 U1326 ( .INP(n118), .Z(n244) );
  DELLN1X2 U1327 ( .INP(n89), .Z(n240) );
  DELLN1X2 U1328 ( .INP(n88), .Z(n236) );
  DELLN1X2 U1329 ( .INP(n79), .Z(n232) );
  DELLN1X2 U1330 ( .INP(n80), .Z(n229) );
  DELLN1X2 U1331 ( .INP(n79), .Z(n233) );
  DELLN1X2 U1332 ( .INP(n88), .Z(n237) );
  DELLN1X2 U1333 ( .INP(n78), .Z(n224) );
  DELLN1X2 U1334 ( .INP(n77), .Z(n220) );
  DELLN1X2 U1335 ( .INP(n77), .Z(n221) );
  DELLN1X2 U1336 ( .INP(n78), .Z(n225) );
  DELLN1X2 U1337 ( .INP(n75), .Z(n217) );
  DELLN1X2 U1338 ( .INP(n76), .Z(n212) );
  DELLN1X2 U1339 ( .INP(n76), .Z(n213) );
  DELLN1X2 U1340 ( .INP(n74), .Z(n209) );
  DELLN1X2 U1341 ( .INP(n73), .Z(n205) );
  DELLN1X2 U1342 ( .INP(n100), .Z(n304) );
  DELLN1X2 U1343 ( .INP(\p[1][63] ), .Z(n509) );
  DELLN1X2 U1344 ( .INP(\p[0][63] ), .Z(n503) );
  DELLN1X2 U1345 ( .INP(n90), .Z(n201) );
  DELLN1X2 U1346 ( .INP(n99), .Z(n295) );
  DELLN1X2 U1347 ( .INP(n102), .Z(n301) );
  DELLN1X2 U1348 ( .INP(n101), .Z(n298) );
  NBUFFX2 U1349 ( .INP(n91), .Z(n293) );
  NBUFFX2 U1350 ( .INP(n98), .Z(n290) );
  NBUFFX2 U1351 ( .INP(n104), .Z(n287) );
  DELLN1X2 U1352 ( .INP(A_reg[31]), .Z(n543) );
  DELLN1X2 U1353 ( .INP(B_reg[31]), .Z(n540) );
  NOR2X0 U1354 ( .IN1(n278), .IN2(n304), .QN(\p[24][26] ) );
  NOR2X0 U1355 ( .IN1(n280), .IN2(n316), .QN(\p[20][21] ) );
  NOR2X0 U1356 ( .IN1(n283), .IN2(n301), .QN(\p[25][25] ) );
  NOR2X0 U1357 ( .IN1(n281), .IN2(n304), .QN(\p[24][25] ) );
  NOR2X0 U1358 ( .IN1(n284), .IN2(n295), .QN(\p[27][27] ) );
  NOR2X0 U1359 ( .IN1(n284), .IN2(n304), .QN(\p[24][24] ) );
  NOR2X0 U1360 ( .IN1(n242), .IN2(n340), .QN(\p[12][24] ) );
  NOR2X0 U1361 ( .IN1(n278), .IN2(n295), .QN(\p[27][29] ) );
  NOR2X0 U1362 ( .IN1(n285), .IN2(n289), .QN(\p[29][29] ) );
  NOR2X0 U1363 ( .IN1(n347), .IN2(n238), .QN(\p[9][22] ) );
  NOR2X0 U1364 ( .IN1(n349), .IN2(n234), .QN(\p[9][23] ) );
  NOR2X0 U1365 ( .IN1(n285), .IN2(n135), .QN(\p[2][2] ) );
  NOR2X0 U1366 ( .IN1(n283), .IN2(n298), .QN(\p[26][26] ) );
  NOR2X0 U1367 ( .IN1(n281), .IN2(n295), .QN(\p[27][28] ) );
  NOR2X0 U1368 ( .IN1(n278), .IN2(n301), .QN(\p[25][27] ) );
  NOR2X0 U1369 ( .IN1(n279), .IN2(n298), .QN(\p[26][28] ) );
  NOR2X0 U1370 ( .IN1(n285), .IN2(n292), .QN(\p[28][28] ) );
  NOR2X0 U1371 ( .IN1(n281), .IN2(n292), .QN(\p[28][29] ) );
  NOR2X0 U1372 ( .IN1(n218), .IN2(n361), .QN(\p[4][22] ) );
  NOR2X0 U1373 ( .IN1(n218), .IN2(n117), .QN(\p[5][23] ) );
  NOR2X0 U1374 ( .IN1(n222), .IN2(n357), .QN(\p[5][22] ) );
  NOR2X0 U1375 ( .IN1(n214), .IN2(n357), .QN(\p[5][24] ) );
  NOR2X0 U1376 ( .IN1(n210), .IN2(n117), .QN(\p[5][25] ) );
  NOR2X0 U1377 ( .IN1(n272), .IN2(n304), .QN(\p[24][28] ) );
  NOR2X0 U1378 ( .IN1(n281), .IN2(n298), .QN(\p[26][27] ) );
  NOR2X0 U1379 ( .IN1(n282), .IN2(n313), .QN(\p[21][22] ) );
  NOR2X0 U1380 ( .IN1(n348), .IN2(n230), .QN(\p[9][24] ) );
  NOR2X0 U1381 ( .IN1(n281), .IN2(n310), .QN(\p[22][23] ) );
  NOR2X0 U1382 ( .IN1(n280), .IN2(n301), .QN(\p[25][26] ) );
  NOR2X0 U1383 ( .IN1(n207), .IN2(n364), .QN(\p[2][23] ) );
  NOR2X0 U1384 ( .IN1(n211), .IN2(n134), .QN(\p[2][22] ) );
  NOR2X0 U1385 ( .IN1(n230), .IN2(n351), .QN(\p[8][23] ) );
  NOR2X0 U1386 ( .IN1(n234), .IN2(n351), .QN(\p[8][22] ) );
  NOR2X0 U1387 ( .IN1(n210), .IN2(n363), .QN(\p[3][23] ) );
  NOR2X0 U1388 ( .IN1(n214), .IN2(n362), .QN(\p[3][22] ) );
  NOR2X0 U1389 ( .IN1(n226), .IN2(n350), .QN(\p[8][24] ) );
  NOR2X0 U1390 ( .IN1(n241), .IN2(n346), .QN(\p[10][23] ) );
  NOR2X0 U1391 ( .IN1(n222), .IN2(n355), .QN(\p[6][23] ) );
  NOR2X0 U1392 ( .IN1(n244), .IN2(n336), .QN(\p[14][26] ) );
  NOR2X0 U1393 ( .IN1(n241), .IN2(n336), .QN(\p[14][27] ) );
  NOR2X0 U1394 ( .IN1(n276), .IN2(n301), .QN(\p[25][28] ) );
  NOR2X0 U1395 ( .IN1(n242), .IN2(n332), .QN(\p[15][27] ) );
  NOR2X0 U1396 ( .IN1(n241), .IN2(n340), .QN(\p[12][25] ) );
  NOR2X0 U1397 ( .IN1(n237), .IN2(n340), .QN(\p[12][26] ) );
  NOR2X0 U1398 ( .IN1(n275), .IN2(n295), .QN(\p[27][30] ) );
  NOR2X0 U1399 ( .IN1(n275), .IN2(n304), .QN(\p[24][27] ) );
  NOR2X0 U1400 ( .IN1(n226), .IN2(n355), .QN(\p[6][22] ) );
  NOR2X0 U1401 ( .IN1(n270), .IN2(n304), .QN(\p[24][29] ) );
  NOR2X0 U1402 ( .IN1(n244), .IN2(n337), .QN(\p[13][25] ) );
  NOR2X0 U1403 ( .IN1(n241), .IN2(n337), .QN(\p[13][26] ) );
  NOR2X0 U1404 ( .IN1(n237), .IN2(n337), .QN(\p[13][27] ) );
  NOR2X0 U1405 ( .IN1(n226), .IN2(n353), .QN(\p[7][23] ) );
  NOR2X0 U1406 ( .IN1(n347), .IN2(n218), .QN(\p[9][27] ) );
  NOR2X0 U1407 ( .IN1(n265), .IN2(n304), .QN(\p[24][30] ) );
  NOR2X0 U1408 ( .IN1(n283), .IN2(n286), .QN(\p[30][30] ) );
  NOR2X0 U1409 ( .IN1(n278), .IN2(n292), .QN(\p[28][30] ) );
  NOR2X0 U1410 ( .IN1(n279), .IN2(n289), .QN(\p[29][31] ) );
  NOR2X0 U1411 ( .IN1(n271), .IN2(n295), .QN(\p[27][32] ) );
  NOR2X0 U1412 ( .IN1(n262), .IN2(n304), .QN(\p[24][31] ) );
  NOR2X0 U1413 ( .IN1(n280), .IN2(n289), .QN(\p[29][30] ) );
  NOR2X0 U1414 ( .IN1(n203), .IN2(n365), .QN(\p[2][24] ) );
  NOR2X0 U1415 ( .IN1(n199), .IN2(n134), .QN(\p[2][25] ) );
  NOR2X0 U1416 ( .IN1(n195), .IN2(n365), .QN(\p[2][26] ) );
  NOR2X0 U1417 ( .IN1(n266), .IN2(n301), .QN(\p[25][31] ) );
  NOR2X0 U1418 ( .IN1(n237), .IN2(n128), .QN(\p[11][25] ) );
  NOR2X0 U1419 ( .IN1(n210), .IN2(n356), .QN(\p[6][26] ) );
  NOR2X0 U1420 ( .IN1(n202), .IN2(n361), .QN(\p[4][26] ) );
  NOR2X0 U1421 ( .IN1(n237), .IN2(n345), .QN(\p[10][24] ) );
  NOR2X0 U1422 ( .IN1(n230), .IN2(n124), .QN(\p[7][22] ) );
  NOR2X0 U1423 ( .IN1(n244), .IN2(n70), .QN(\p[10][22] ) );
  NOR2X0 U1424 ( .IN1(n233), .IN2(n344), .QN(\p[10][25] ) );
  NOR2X0 U1425 ( .IN1(n214), .IN2(n354), .QN(\p[7][26] ) );
  NOR2X0 U1426 ( .IN1(n214), .IN2(n132), .QN(\p[6][25] ) );
  NOR2X0 U1427 ( .IN1(n198), .IN2(n358), .QN(\p[5][28] ) );
  NOR2X0 U1428 ( .IN1(n206), .IN2(n357), .QN(\p[5][26] ) );
  NOR2X0 U1429 ( .IN1(n202), .IN2(n357), .QN(\p[5][27] ) );
  NOR2X0 U1430 ( .IN1(n273), .IN2(n295), .QN(\p[27][31] ) );
  NOR2X0 U1431 ( .IN1(n348), .IN2(n226), .QN(\p[9][25] ) );
  NOR2X0 U1432 ( .IN1(n348), .IN2(n222), .QN(\p[9][26] ) );
  NOR2X0 U1433 ( .IN1(n272), .IN2(n292), .QN(\p[28][32] ) );
  NOR2X0 U1434 ( .IN1(n206), .IN2(n363), .QN(\p[3][24] ) );
  NOR2X0 U1435 ( .IN1(n202), .IN2(n362), .QN(\p[3][25] ) );
  NOR2X0 U1436 ( .IN1(n198), .IN2(n362), .QN(\p[3][26] ) );
  NOR2X0 U1437 ( .IN1(n262), .IN2(n316), .QN(\p[20][27] ) );
  NOR2X0 U1438 ( .IN1(n276), .IN2(n298), .QN(\p[26][29] ) );
  NOR2X0 U1439 ( .IN1(n218), .IN2(n350), .QN(\p[8][26] ) );
  NOR2X0 U1440 ( .IN1(n222), .IN2(n350), .QN(\p[8][25] ) );
  NOR2X0 U1441 ( .IN1(n151), .IN2(n313), .QN(\p[21][28] ) );
  NOR2X0 U1442 ( .IN1(n240), .IN2(n326), .QN(\p[17][30] ) );
  NOR2X0 U1443 ( .IN1(n243), .IN2(n326), .QN(\p[17][29] ) );
  NOR2X0 U1444 ( .IN1(n218), .IN2(n355), .QN(\p[6][24] ) );
  NOR2X0 U1445 ( .IN1(n244), .IN2(n323), .QN(\p[18][30] ) );
  NOR2X0 U1446 ( .IN1(n240), .IN2(n323), .QN(\p[18][31] ) );
  NOR2X0 U1447 ( .IN1(n210), .IN2(n361), .QN(\p[4][24] ) );
  NOR2X0 U1448 ( .IN1(n206), .IN2(n359), .QN(\p[4][25] ) );
  NOR2X0 U1449 ( .IN1(n229), .IN2(n335), .QN(\p[14][30] ) );
  NOR2X0 U1450 ( .IN1(n233), .IN2(n108), .QN(\p[14][29] ) );
  NOR2X0 U1451 ( .IN1(n237), .IN2(n336), .QN(\p[14][28] ) );
  NOR2X0 U1452 ( .IN1(n275), .IN2(n289), .QN(\p[29][32] ) );
  NOR2X0 U1453 ( .IN1(n270), .IN2(n298), .QN(\p[26][31] ) );
  NOR2X0 U1454 ( .IN1(n276), .IN2(n292), .QN(\p[28][31] ) );
  NOR2X0 U1455 ( .IN1(n218), .IN2(n353), .QN(\p[7][25] ) );
  NOR2X0 U1456 ( .IN1(n233), .IN2(n333), .QN(\p[15][30] ) );
  NOR2X0 U1457 ( .IN1(n225), .IN2(n340), .QN(\p[12][29] ) );
  NOR2X0 U1458 ( .IN1(n237), .IN2(n332), .QN(\p[15][29] ) );
  NOR2X0 U1459 ( .IN1(n241), .IN2(n332), .QN(\p[15][28] ) );
  NOR2X0 U1460 ( .IN1(n229), .IN2(n340), .QN(\p[12][28] ) );
  NOR2X0 U1461 ( .IN1(n233), .IN2(n340), .QN(\p[12][27] ) );
  NOR2X0 U1462 ( .IN1(n236), .IN2(n329), .QN(\p[16][30] ) );
  NOR2X0 U1463 ( .IN1(n240), .IN2(n330), .QN(\p[16][29] ) );
  NOR2X0 U1464 ( .IN1(n243), .IN2(n329), .QN(\p[16][28] ) );
  NOR2X0 U1465 ( .IN1(n222), .IN2(n353), .QN(\p[7][24] ) );
  NOR2X0 U1466 ( .IN1(n225), .IN2(n337), .QN(\p[13][30] ) );
  NOR2X0 U1467 ( .IN1(n229), .IN2(n337), .QN(\p[13][29] ) );
  NOR2X0 U1468 ( .IN1(n233), .IN2(n337), .QN(\p[13][28] ) );
  NOR2X0 U1469 ( .IN1(n137), .IN2(n301), .QN(\p[25][30] ) );
  NOR2X0 U1470 ( .IN1(n254), .IN2(n316), .QN(\p[20][29] ) );
  NOR2X0 U1471 ( .IN1(n254), .IN2(n313), .QN(\p[21][30] ) );
  NOR2X0 U1472 ( .IN1(n347), .IN2(n206), .QN(\p[9][30] ) );
  NOR2X0 U1473 ( .IN1(n349), .IN2(n210), .QN(\p[9][29] ) );
  NOR2X0 U1474 ( .IN1(n265), .IN2(n295), .QN(\p[27][33] ) );
  NOR2X0 U1475 ( .IN1(n254), .IN2(n310), .QN(\p[22][31] ) );
  NOR2X0 U1476 ( .IN1(n225), .IN2(n342), .QN(\p[11][28] ) );
  NOR2X0 U1477 ( .IN1(n229), .IN2(n128), .QN(\p[11][27] ) );
  NOR2X0 U1478 ( .IN1(n267), .IN2(n289), .QN(\p[29][35] ) );
  NOR2X0 U1479 ( .IN1(n267), .IN2(n298), .QN(\p[26][32] ) );
  NOR2X0 U1480 ( .IN1(n271), .IN2(n286), .QN(\p[30][35] ) );
  NOR2X0 U1481 ( .IN1(n256), .IN2(n301), .QN(\p[25][34] ) );
  NOR2X0 U1482 ( .IN1(n261), .IN2(n295), .QN(\p[27][34] ) );
  NOR2X0 U1483 ( .IN1(n263), .IN2(n292), .QN(\p[28][35] ) );
  NOR2X0 U1484 ( .IN1(n151), .IN2(n310), .QN(\p[22][29] ) );
  NOR2X0 U1485 ( .IN1(n257), .IN2(n304), .QN(\p[24][33] ) );
  NOR2X0 U1486 ( .IN1(n183), .IN2(n365), .QN(\p[2][29] ) );
  NOR2X0 U1487 ( .IN1(n266), .IN2(n292), .QN(\p[28][34] ) );
  NOR2X0 U1488 ( .IN1(n151), .IN2(n301), .QN(\p[25][32] ) );
  NOR2X0 U1489 ( .IN1(n190), .IN2(n359), .QN(\p[4][29] ) );
  NOR2X0 U1490 ( .IN1(n194), .IN2(n361), .QN(\p[4][28] ) );
  NOR2X0 U1491 ( .IN1(n198), .IN2(n359), .QN(\p[4][27] ) );
  NOR2X0 U1492 ( .IN1(n202), .IN2(n124), .QN(\p[7][29] ) );
  NOR2X0 U1493 ( .IN1(n206), .IN2(n354), .QN(\p[7][28] ) );
  NOR2X0 U1494 ( .IN1(n190), .IN2(n357), .QN(\p[5][30] ) );
  NOR2X0 U1495 ( .IN1(n186), .IN2(n358), .QN(\p[5][31] ) );
  NOR2X0 U1496 ( .IN1(n194), .IN2(n117), .QN(\p[5][29] ) );
  NOR2X0 U1497 ( .IN1(n187), .IN2(n364), .QN(\p[2][28] ) );
  NOR2X0 U1498 ( .IN1(n198), .IN2(n131), .QN(\p[6][29] ) );
  NOR2X0 U1499 ( .IN1(n272), .IN2(n286), .QN(\p[30][34] ) );
  NOR2X0 U1500 ( .IN1(n348), .IN2(n214), .QN(\p[9][28] ) );
  NOR2X0 U1501 ( .IN1(n258), .IN2(n298), .QN(\p[26][34] ) );
  NOR2X0 U1502 ( .IN1(n259), .IN2(n295), .QN(\p[27][35] ) );
  NOR2X0 U1503 ( .IN1(n260), .IN2(n304), .QN(\p[24][32] ) );
  NOR2X0 U1504 ( .IN1(n210), .IN2(n351), .QN(\p[8][28] ) );
  NOR2X0 U1505 ( .IN1(n214), .IN2(n351), .QN(\p[8][27] ) );
  NOR2X0 U1506 ( .IN1(n191), .IN2(n365), .QN(\p[2][27] ) );
  NOR2X0 U1507 ( .IN1(n202), .IN2(n355), .QN(\p[6][28] ) );
  NOR2X0 U1508 ( .IN1(n206), .IN2(n355), .QN(\p[6][27] ) );
  NOR2X0 U1509 ( .IN1(n246), .IN2(n316), .QN(\p[20][31] ) );
  NOR2X0 U1510 ( .IN1(n251), .IN2(n316), .QN(\p[20][30] ) );
  NOR2X0 U1511 ( .IN1(n251), .IN2(n313), .QN(\p[21][31] ) );
  NOR2X0 U1512 ( .IN1(n243), .IN2(n317), .QN(\p[20][32] ) );
  NOR2X0 U1513 ( .IN1(n232), .IN2(n326), .QN(\p[17][32] ) );
  NOR2X0 U1514 ( .IN1(n240), .IN2(n317), .QN(\p[20][33] ) );
  NOR2X0 U1515 ( .IN1(n228), .IN2(n326), .QN(\p[17][33] ) );
  NOR2X0 U1516 ( .IN1(n236), .IN2(n326), .QN(\p[17][31] ) );
  NOR2X0 U1517 ( .IN1(n260), .IN2(n301), .QN(\p[25][33] ) );
  NOR2X0 U1518 ( .IN1(n150), .IN2(n298), .QN(\p[26][33] ) );
  NOR2X0 U1519 ( .IN1(n252), .IN2(n304), .QN(\p[24][34] ) );
  NOR2X0 U1520 ( .IN1(n186), .IN2(n144), .QN(\p[3][29] ) );
  NOR2X0 U1521 ( .IN1(n190), .IN2(n363), .QN(\p[3][28] ) );
  NOR2X0 U1522 ( .IN1(n194), .IN2(n144), .QN(\p[3][27] ) );
  NOR2X0 U1523 ( .IN1(n245), .IN2(n314), .QN(\p[21][33] ) );
  NOR2X0 U1524 ( .IN1(n236), .IN2(n323), .QN(\p[18][32] ) );
  NOR2X0 U1525 ( .IN1(n232), .IN2(n323), .QN(\p[18][33] ) );
  NOR2X0 U1526 ( .IN1(n240), .IN2(n314), .QN(\p[21][34] ) );
  NOR2X0 U1527 ( .IN1(n228), .IN2(n323), .QN(\p[18][34] ) );
  NOR2X0 U1528 ( .IN1(n210), .IN2(n353), .QN(\p[7][27] ) );
  NOR2X0 U1529 ( .IN1(n221), .IN2(n335), .QN(\p[14][32] ) );
  NOR2X0 U1530 ( .IN1(n217), .IN2(n335), .QN(\p[14][33] ) );
  NOR2X0 U1531 ( .IN1(n225), .IN2(n335), .QN(\p[14][31] ) );
  NOR2X0 U1532 ( .IN1(n233), .IN2(n127), .QN(\p[11][26] ) );
  NOR2X0 U1533 ( .IN1(n137), .IN2(n289), .QN(\p[29][34] ) );
  NOR2X0 U1534 ( .IN1(n213), .IN2(n341), .QN(\p[12][32] ) );
  NOR2X0 U1535 ( .IN1(n225), .IN2(n333), .QN(\p[15][32] ) );
  NOR2X0 U1536 ( .IN1(n217), .IN2(n340), .QN(\p[12][31] ) );
  NOR2X0 U1537 ( .IN1(n229), .IN2(n332), .QN(\p[15][31] ) );
  NOR2X0 U1538 ( .IN1(n221), .IN2(n333), .QN(\p[15][33] ) );
  NOR2X0 U1539 ( .IN1(n221), .IN2(n339), .QN(\p[12][30] ) );
  NOR2X0 U1540 ( .IN1(n240), .IN2(n320), .QN(\p[19][32] ) );
  NOR2X0 U1541 ( .IN1(n242), .IN2(n320), .QN(\p[19][31] ) );
  NOR2X0 U1542 ( .IN1(n228), .IN2(n329), .QN(\p[16][32] ) );
  NOR2X0 U1543 ( .IN1(n232), .IN2(n330), .QN(\p[16][31] ) );
  NOR2X0 U1544 ( .IN1(n236), .IN2(n320), .QN(\p[19][33] ) );
  NOR2X0 U1545 ( .IN1(n224), .IN2(n330), .QN(\p[16][33] ) );
  NOR2X0 U1546 ( .IN1(n217), .IN2(n337), .QN(\p[13][32] ) );
  NOR2X0 U1547 ( .IN1(n221), .IN2(n337), .QN(\p[13][31] ) );
  NOR2X0 U1548 ( .IN1(n213), .IN2(n337), .QN(\p[13][33] ) );
  NOR2X0 U1549 ( .IN1(n268), .IN2(n292), .QN(\p[28][33] ) );
  NBUFFX2 U1550 ( .INP(\p[58][63] ), .Z(n474) );
  NBUFFX2 U1551 ( .INP(\p[58][63] ), .Z(n476) );
  NOR2X0 U1552 ( .IN1(n254), .IN2(n295), .QN(\p[27][36] ) );
  NOR2X0 U1553 ( .IN1(n256), .IN2(n307), .QN(\p[23][32] ) );
  NOR2X0 U1554 ( .IN1(n349), .IN2(n198), .QN(\p[9][32] ) );
  NOR2X0 U1555 ( .IN1(n250), .IN2(n286), .QN(\p[30][40] ) );
  NOR2X0 U1556 ( .IN1(n247), .IN2(n308), .QN(\p[23][34] ) );
  NOR2X0 U1557 ( .IN1(n252), .IN2(n308), .QN(\p[23][33] ) );
  NOR2X0 U1558 ( .IN1(n244), .IN2(n308), .QN(\p[23][35] ) );
  NOR2X0 U1559 ( .IN1(n261), .IN2(n286), .QN(\p[30][37] ) );
  NOR2X0 U1560 ( .IN1(n209), .IN2(n342), .QN(\p[11][32] ) );
  NOR2X0 U1561 ( .IN1(n151), .IN2(n289), .QN(\p[29][36] ) );
  NOR2X0 U1562 ( .IN1(n253), .IN2(n301), .QN(\p[25][35] ) );
  NOR2X0 U1563 ( .IN1(n253), .IN2(n292), .QN(\p[28][38] ) );
  NOR2X0 U1564 ( .IN1(n213), .IN2(n128), .QN(\p[11][31] ) );
  NOR2X0 U1565 ( .IN1(n194), .IN2(n356), .QN(\p[6][30] ) );
  NOR2X0 U1566 ( .IN1(n174), .IN2(n356), .QN(\p[6][35] ) );
  NOR2X0 U1567 ( .IN1(n186), .IN2(n361), .QN(\p[4][30] ) );
  NOR2X0 U1568 ( .IN1(n182), .IN2(n359), .QN(\p[4][31] ) );
  NOR2X0 U1569 ( .IN1(n178), .IN2(n361), .QN(\p[4][32] ) );
  NOR2X0 U1570 ( .IN1(n209), .IN2(n345), .QN(\p[10][31] ) );
  NOR2X0 U1571 ( .IN1(n197), .IN2(n344), .QN(\p[10][34] ) );
  NOR2X0 U1572 ( .IN1(n193), .IN2(n344), .QN(\p[10][35] ) );
  NOR2X0 U1573 ( .IN1(n186), .IN2(n124), .QN(\p[7][33] ) );
  NOR2X0 U1574 ( .IN1(n205), .IN2(n127), .QN(\p[11][33] ) );
  NOR2X0 U1575 ( .IN1(n201), .IN2(n128), .QN(\p[11][34] ) );
  NOR2X0 U1576 ( .IN1(n213), .IN2(n344), .QN(\p[10][30] ) );
  NOR2X0 U1577 ( .IN1(n198), .IN2(n354), .QN(\p[7][30] ) );
  NOR2X0 U1578 ( .IN1(n182), .IN2(n354), .QN(\p[7][34] ) );
  NOR2X0 U1579 ( .IN1(n190), .IN2(n132), .QN(\p[6][31] ) );
  NOR2X0 U1580 ( .IN1(n186), .IN2(n132), .QN(\p[6][32] ) );
  NOR2X0 U1581 ( .IN1(n182), .IN2(n117), .QN(\p[5][32] ) );
  NOR2X0 U1582 ( .IN1(n178), .IN2(n358), .QN(\p[5][33] ) );
  NOR2X0 U1583 ( .IN1(n179), .IN2(n365), .QN(\p[2][30] ) );
  NOR2X0 U1584 ( .IN1(n194), .IN2(n352), .QN(\p[7][31] ) );
  NOR2X0 U1585 ( .IN1(n178), .IN2(n131), .QN(\p[6][34] ) );
  NOR2X0 U1586 ( .IN1(n259), .IN2(n309), .QN(\p[23][31] ) );
  NOR2X0 U1587 ( .IN1(n348), .IN2(n202), .QN(\p[9][31] ) );
  NOR2X0 U1588 ( .IN1(n260), .IN2(n289), .QN(\p[29][37] ) );
  NOR2X0 U1589 ( .IN1(n255), .IN2(n298), .QN(\p[26][35] ) );
  NOR2X0 U1590 ( .IN1(n255), .IN2(n289), .QN(\p[29][38] ) );
  NOR2X0 U1591 ( .IN1(n259), .IN2(n286), .QN(\p[30][38] ) );
  NOR2X0 U1592 ( .IN1(n255), .IN2(n286), .QN(\p[30][39] ) );
  NOR2X0 U1593 ( .IN1(n198), .IN2(n351), .QN(\p[8][31] ) );
  NOR2X0 U1594 ( .IN1(n175), .IN2(n365), .QN(\p[2][31] ) );
  NOR2X0 U1595 ( .IN1(n252), .IN2(n298), .QN(\p[26][36] ) );
  NOR2X0 U1596 ( .IN1(n251), .IN2(n289), .QN(\p[29][39] ) );
  NOR2X0 U1597 ( .IN1(n190), .IN2(n350), .QN(\p[8][33] ) );
  NOR2X0 U1598 ( .IN1(n194), .IN2(n350), .QN(\p[8][32] ) );
  NOR2X0 U1599 ( .IN1(n255), .IN2(n292), .QN(\p[28][37] ) );
  NOR2X0 U1600 ( .IN1(n249), .IN2(n313), .QN(\p[21][32] ) );
  NOR2X0 U1601 ( .IN1(n236), .IN2(n317), .QN(\p[20][34] ) );
  NOR2X0 U1602 ( .IN1(n224), .IN2(n326), .QN(\p[17][34] ) );
  NOR2X0 U1603 ( .IN1(n232), .IN2(n317), .QN(\p[20][35] ) );
  NOR2X0 U1604 ( .IN1(n220), .IN2(n326), .QN(\p[17][35] ) );
  NOR2X0 U1605 ( .IN1(n228), .IN2(n317), .QN(\p[20][36] ) );
  NOR2X0 U1606 ( .IN1(n216), .IN2(n326), .QN(\p[17][36] ) );
  NOR2X0 U1607 ( .IN1(n224), .IN2(n317), .QN(\p[20][37] ) );
  NOR2X0 U1608 ( .IN1(n212), .IN2(n326), .QN(\p[17][37] ) );
  NOR2X0 U1609 ( .IN1(n208), .IN2(n326), .QN(\p[17][38] ) );
  NOR2X0 U1610 ( .IN1(n220), .IN2(n317), .QN(\p[20][38] ) );
  NOR2X0 U1611 ( .IN1(n204), .IN2(n326), .QN(\p[17][39] ) );
  NOR2X0 U1612 ( .IN1(n245), .IN2(n299), .QN(\p[26][38] ) );
  NOR2X0 U1613 ( .IN1(n216), .IN2(n317), .QN(\p[20][39] ) );
  NOR2X0 U1614 ( .IN1(n239), .IN2(n299), .QN(\p[26][39] ) );
  NOR2X0 U1615 ( .IN1(n243), .IN2(n290), .QN(\p[29][41] ) );
  NOR2X0 U1616 ( .IN1(n235), .IN2(n299), .QN(\p[26][40] ) );
  NOR2X0 U1617 ( .IN1(n249), .IN2(n298), .QN(\p[26][37] ) );
  NOR2X0 U1618 ( .IN1(n248), .IN2(n289), .QN(\p[29][40] ) );
  NOR2X0 U1619 ( .IN1(n260), .IN2(n292), .QN(\p[28][36] ) );
  NOR2X0 U1620 ( .IN1(n251), .IN2(n295), .QN(\p[27][37] ) );
  NOR2X0 U1621 ( .IN1(n182), .IN2(n362), .QN(\p[3][30] ) );
  NOR2X0 U1622 ( .IN1(n182), .IN2(n355), .QN(\p[6][33] ) );
  NOR2X0 U1623 ( .IN1(n245), .IN2(n296), .QN(\p[27][39] ) );
  NOR2X0 U1624 ( .IN1(n242), .IN2(n305), .QN(\p[24][36] ) );
  NOR2X0 U1625 ( .IN1(n236), .IN2(n314), .QN(\p[21][35] ) );
  NOR2X0 U1626 ( .IN1(n224), .IN2(n323), .QN(\p[18][35] ) );
  NOR2X0 U1627 ( .IN1(n220), .IN2(n323), .QN(\p[18][36] ) );
  NOR2X0 U1628 ( .IN1(n232), .IN2(n314), .QN(\p[21][36] ) );
  NOR2X0 U1629 ( .IN1(n239), .IN2(n305), .QN(\p[24][37] ) );
  NOR2X0 U1630 ( .IN1(n235), .IN2(n305), .QN(\p[24][38] ) );
  NOR2X0 U1631 ( .IN1(n216), .IN2(n323), .QN(\p[18][37] ) );
  NOR2X0 U1632 ( .IN1(n228), .IN2(n314), .QN(\p[21][37] ) );
  NOR2X0 U1633 ( .IN1(n212), .IN2(n323), .QN(\p[18][38] ) );
  NOR2X0 U1634 ( .IN1(n224), .IN2(n314), .QN(\p[21][38] ) );
  NOR2X0 U1635 ( .IN1(n239), .IN2(n296), .QN(\p[27][40] ) );
  NOR2X0 U1636 ( .IN1(n208), .IN2(n323), .QN(\p[18][39] ) );
  NOR2X0 U1637 ( .IN1(n220), .IN2(n314), .QN(\p[21][39] ) );
  NOR2X0 U1638 ( .IN1(n231), .IN2(n305), .QN(\p[24][39] ) );
  NOR2X0 U1639 ( .IN1(n235), .IN2(n296), .QN(\p[27][41] ) );
  NOR2X0 U1640 ( .IN1(n204), .IN2(n323), .QN(\p[18][40] ) );
  NOR2X0 U1641 ( .IN1(n227), .IN2(n305), .QN(\p[24][40] ) );
  NOR2X0 U1642 ( .IN1(n246), .IN2(n304), .QN(\p[24][35] ) );
  NOR2X0 U1643 ( .IN1(n249), .IN2(n295), .QN(\p[27][38] ) );
  NOR2X0 U1644 ( .IN1(n205), .IN2(n344), .QN(\p[10][32] ) );
  NOR2X0 U1645 ( .IN1(n201), .IN2(n345), .QN(\p[10][33] ) );
  NOR2X0 U1646 ( .IN1(n252), .IN2(n310), .QN(\p[22][32] ) );
  NOR2X0 U1647 ( .IN1(n249), .IN2(n310), .QN(\p[22][33] ) );
  NOR2X0 U1648 ( .IN1(n213), .IN2(n335), .QN(\p[14][34] ) );
  NOR2X0 U1649 ( .IN1(n209), .IN2(n335), .QN(\p[14][35] ) );
  NOR2X0 U1650 ( .IN1(n217), .IN2(n342), .QN(\p[11][30] ) );
  NOR2X0 U1651 ( .IN1(n221), .IN2(n342), .QN(\p[11][29] ) );
  NOR2X0 U1652 ( .IN1(n205), .IN2(n335), .QN(\p[14][36] ) );
  NOR2X0 U1653 ( .IN1(n201), .IN2(n335), .QN(\p[14][37] ) );
  NOR2X0 U1654 ( .IN1(n209), .IN2(n339), .QN(\p[12][33] ) );
  NOR2X0 U1655 ( .IN1(n217), .IN2(n332), .QN(\p[15][34] ) );
  NOR2X0 U1656 ( .IN1(n205), .IN2(n332), .QN(\p[15][37] ) );
  NOR2X0 U1657 ( .IN1(n205), .IN2(n339), .QN(\p[12][34] ) );
  NOR2X0 U1658 ( .IN1(n213), .IN2(n331), .QN(\p[15][35] ) );
  NOR2X0 U1659 ( .IN1(n209), .IN2(n331), .QN(\p[15][36] ) );
  NOR2X0 U1660 ( .IN1(n201), .IN2(n339), .QN(\p[12][35] ) );
  NOR2X0 U1661 ( .IN1(n201), .IN2(n333), .QN(\p[15][38] ) );
  NOR2X0 U1662 ( .IN1(n190), .IN2(n353), .QN(\p[7][32] ) );
  NOR2X0 U1663 ( .IN1(n242), .IN2(n311), .QN(\p[22][34] ) );
  NOR2X0 U1664 ( .IN1(n232), .IN2(n320), .QN(\p[19][34] ) );
  NOR2X0 U1665 ( .IN1(n240), .IN2(n311), .QN(\p[22][35] ) );
  NOR2X0 U1666 ( .IN1(n220), .IN2(n329), .QN(\p[16][34] ) );
  NOR2X0 U1667 ( .IN1(n228), .IN2(n320), .QN(\p[19][35] ) );
  NOR2X0 U1668 ( .IN1(n236), .IN2(n311), .QN(\p[22][36] ) );
  NOR2X0 U1669 ( .IN1(n224), .IN2(n320), .QN(\p[19][36] ) );
  NOR2X0 U1670 ( .IN1(n216), .IN2(n330), .QN(\p[16][35] ) );
  NOR2X0 U1671 ( .IN1(n239), .IN2(n302), .QN(\p[25][38] ) );
  NOR2X0 U1672 ( .IN1(n243), .IN2(n302), .QN(\p[25][37] ) );
  NOR2X0 U1673 ( .IN1(n212), .IN2(n329), .QN(\p[16][36] ) );
  NOR2X0 U1674 ( .IN1(n220), .IN2(n320), .QN(\p[19][37] ) );
  NOR2X0 U1675 ( .IN1(n232), .IN2(n311), .QN(\p[22][37] ) );
  NOR2X0 U1676 ( .IN1(n208), .IN2(n330), .QN(\p[16][37] ) );
  NOR2X0 U1677 ( .IN1(n204), .IN2(n329), .QN(\p[16][38] ) );
  NOR2X0 U1678 ( .IN1(n216), .IN2(n320), .QN(\p[19][38] ) );
  NOR2X0 U1679 ( .IN1(n228), .IN2(n311), .QN(\p[22][38] ) );
  NOR2X0 U1680 ( .IN1(n200), .IN2(n330), .QN(\p[16][39] ) );
  NOR2X0 U1681 ( .IN1(n245), .IN2(n293), .QN(\p[28][40] ) );
  NOR2X0 U1682 ( .IN1(n212), .IN2(n320), .QN(\p[19][39] ) );
  NOR2X0 U1683 ( .IN1(n224), .IN2(n311), .QN(\p[22][39] ) );
  NOR2X0 U1684 ( .IN1(n235), .IN2(n302), .QN(\p[25][39] ) );
  NOR2X0 U1685 ( .IN1(n239), .IN2(n293), .QN(\p[28][41] ) );
  NOR2X0 U1686 ( .IN1(n231), .IN2(n302), .QN(\p[25][40] ) );
  NOR2X0 U1687 ( .IN1(n247), .IN2(n292), .QN(\p[28][39] ) );
  NOR2X0 U1688 ( .IN1(n246), .IN2(n301), .QN(\p[25][36] ) );
  NOR2X0 U1689 ( .IN1(n174), .IN2(n359), .QN(\p[4][33] ) );
  NOR2X0 U1690 ( .IN1(n209), .IN2(n337), .QN(\p[13][34] ) );
  NOR2X0 U1691 ( .IN1(n201), .IN2(n337), .QN(\p[13][36] ) );
  NOR2X0 U1692 ( .IN1(n205), .IN2(n337), .QN(\p[13][35] ) );
  NOR2X0 U1693 ( .IN1(n247), .IN2(n286), .QN(\p[30][41] ) );
  NBUFFX2 U1694 ( .INP(\p[58][63] ), .Z(n475) );
  NOR2X0 U1695 ( .IN1(n235), .IN2(n308), .QN(\p[23][37] ) );
  NOR2X0 U1696 ( .IN1(n227), .IN2(n308), .QN(\p[23][39] ) );
  NOR2X0 U1697 ( .IN1(n193), .IN2(n127), .QN(\p[11][36] ) );
  NOR2X0 U1698 ( .IN1(n197), .IN2(n128), .QN(\p[11][35] ) );
  NOR2X0 U1699 ( .IN1(n239), .IN2(n307), .QN(\p[23][36] ) );
  NOR2X0 U1700 ( .IN1(n174), .IN2(n124), .QN(\p[7][36] ) );
  NOR2X0 U1701 ( .IN1(n189), .IN2(n342), .QN(\p[11][37] ) );
  NOR2X0 U1702 ( .IN1(n189), .IN2(n345), .QN(\p[10][36] ) );
  NOR2X0 U1703 ( .IN1(n178), .IN2(n352), .QN(\p[7][35] ) );
  NOR2X0 U1704 ( .IN1(n170), .IN2(n352), .QN(\p[7][37] ) );
  NOR2X0 U1705 ( .IN1(n182), .IN2(n351), .QN(\p[8][35] ) );
  NOR2X0 U1706 ( .IN1(n174), .IN2(n351), .QN(\p[8][37] ) );
  NOR2X0 U1707 ( .IN1(n170), .IN2(n350), .QN(\p[8][38] ) );
  NOR2X0 U1708 ( .IN1(n200), .IN2(n326), .QN(\p[17][40] ) );
  NOR2X0 U1709 ( .IN1(n212), .IN2(n317), .QN(\p[20][40] ) );
  NOR2X0 U1710 ( .IN1(n239), .IN2(n290), .QN(\p[29][42] ) );
  NOR2X0 U1711 ( .IN1(n208), .IN2(n317), .QN(\p[20][41] ) );
  NOR2X0 U1712 ( .IN1(n231), .IN2(n299), .QN(\p[26][41] ) );
  NOR2X0 U1713 ( .IN1(n235), .IN2(n290), .QN(\p[29][43] ) );
  NOR2X0 U1714 ( .IN1(n204), .IN2(n317), .QN(\p[20][42] ) );
  NOR2X0 U1715 ( .IN1(n227), .IN2(n299), .QN(\p[26][42] ) );
  NOR2X0 U1716 ( .IN1(n216), .IN2(n314), .QN(\p[21][40] ) );
  NOR2X0 U1717 ( .IN1(n231), .IN2(n296), .QN(\p[27][42] ) );
  NOR2X0 U1718 ( .IN1(n200), .IN2(n323), .QN(\p[18][41] ) );
  NOR2X0 U1719 ( .IN1(n212), .IN2(n314), .QN(\p[21][41] ) );
  NOR2X0 U1720 ( .IN1(n223), .IN2(n305), .QN(\p[24][41] ) );
  NOR2X0 U1721 ( .IN1(n227), .IN2(n296), .QN(\p[27][43] ) );
  NOR2X0 U1722 ( .IN1(n208), .IN2(n314), .QN(\p[21][42] ) );
  NOR2X0 U1723 ( .IN1(n219), .IN2(n305), .QN(\p[24][42] ) );
  NOR2X0 U1724 ( .IN1(n223), .IN2(n296), .QN(\p[27][44] ) );
  NOR2X0 U1725 ( .IN1(n215), .IN2(n305), .QN(\p[24][43] ) );
  NOR2X0 U1726 ( .IN1(n185), .IN2(n344), .QN(\p[10][37] ) );
  NOR2X0 U1727 ( .IN1(n181), .IN2(n345), .QN(\p[10][38] ) );
  NOR2X0 U1728 ( .IN1(n197), .IN2(n339), .QN(\p[12][36] ) );
  NOR2X0 U1729 ( .IN1(n193), .IN2(n339), .QN(\p[12][37] ) );
  NOR2X0 U1730 ( .IN1(n208), .IN2(n320), .QN(\p[19][40] ) );
  NOR2X0 U1731 ( .IN1(n220), .IN2(n311), .QN(\p[22][40] ) );
  NOR2X0 U1732 ( .IN1(n235), .IN2(n293), .QN(\p[28][42] ) );
  NOR2X0 U1733 ( .IN1(n204), .IN2(n320), .QN(\p[19][41] ) );
  NOR2X0 U1734 ( .IN1(n216), .IN2(n311), .QN(\p[22][41] ) );
  NOR2X0 U1735 ( .IN1(n227), .IN2(n302), .QN(\p[25][41] ) );
  NOR2X0 U1736 ( .IN1(n231), .IN2(n293), .QN(\p[28][43] ) );
  NOR2X0 U1737 ( .IN1(n212), .IN2(n311), .QN(\p[22][42] ) );
  NOR2X0 U1738 ( .IN1(n200), .IN2(n320), .QN(\p[19][42] ) );
  NOR2X0 U1739 ( .IN1(n223), .IN2(n302), .QN(\p[25][42] ) );
  NOR2X0 U1740 ( .IN1(n227), .IN2(n293), .QN(\p[28][44] ) );
  NOR2X0 U1741 ( .IN1(n219), .IN2(n302), .QN(\p[25][43] ) );
  NOR2X0 U1742 ( .IN1(n197), .IN2(n338), .QN(\p[13][37] ) );
  NOR2X0 U1743 ( .IN1(n193), .IN2(n338), .QN(\p[13][38] ) );
  NOR2X0 U1744 ( .IN1(n234), .IN2(n287), .QN(\p[30][44] ) );
  NOR2X0 U1745 ( .IN1(n244), .IN2(n287), .QN(\p[30][42] ) );
  NOR2X0 U1746 ( .IN1(n238), .IN2(n287), .QN(\p[30][43] ) );
  NBUFFX2 U1747 ( .INP(\p[58][63] ), .Z(n473) );
  NOR2X0 U1748 ( .IN1(n215), .IN2(n308), .QN(\p[23][42] ) );
  NOR2X0 U1749 ( .IN1(n181), .IN2(n343), .QN(\p[11][39] ) );
  NOR2X0 U1750 ( .IN1(n231), .IN2(n307), .QN(\p[23][38] ) );
  NOR2X0 U1751 ( .IN1(n223), .IN2(n309), .QN(\p[23][40] ) );
  NOR2X0 U1752 ( .IN1(n211), .IN2(n305), .QN(\p[24][44] ) );
  NOR2X0 U1753 ( .IN1(n207), .IN2(n305), .QN(\p[24][45] ) );
  NOR2X0 U1754 ( .IN1(n211), .IN2(n296), .QN(\p[27][47] ) );
  NOR2X0 U1755 ( .IN1(n203), .IN2(n305), .QN(\p[24][46] ) );
  NOR2X0 U1756 ( .IN1(n196), .IN2(n327), .QN(\p[17][41] ) );
  NOR2X0 U1757 ( .IN1(n231), .IN2(n290), .QN(\p[29][44] ) );
  NOR2X0 U1758 ( .IN1(n200), .IN2(n317), .QN(\p[20][43] ) );
  NOR2X0 U1759 ( .IN1(n223), .IN2(n299), .QN(\p[26][43] ) );
  NOR2X0 U1760 ( .IN1(n227), .IN2(n290), .QN(\p[29][45] ) );
  NOR2X0 U1761 ( .IN1(n219), .IN2(n299), .QN(\p[26][44] ) );
  NOR2X0 U1762 ( .IN1(n223), .IN2(n290), .QN(\p[29][46] ) );
  NOR2X0 U1763 ( .IN1(n215), .IN2(n299), .QN(\p[26][45] ) );
  NOR2X0 U1764 ( .IN1(n204), .IN2(n314), .QN(\p[21][43] ) );
  NOR2X0 U1765 ( .IN1(n219), .IN2(n296), .QN(\p[27][45] ) );
  NOR2X0 U1766 ( .IN1(n200), .IN2(n314), .QN(\p[21][44] ) );
  NOR2X0 U1767 ( .IN1(n215), .IN2(n296), .QN(\p[27][46] ) );
  NOR2X0 U1768 ( .IN1(n177), .IN2(n344), .QN(\p[10][39] ) );
  NOR2X0 U1769 ( .IN1(n173), .IN2(n345), .QN(\p[10][40] ) );
  NOR2X0 U1770 ( .IN1(n222), .IN2(n287), .QN(\p[30][47] ) );
  NOR2X0 U1771 ( .IN1(n211), .IN2(n302), .QN(\p[25][45] ) );
  NOR2X0 U1772 ( .IN1(n207), .IN2(n302), .QN(\p[25][46] ) );
  NOR2X0 U1773 ( .IN1(n185), .IN2(n127), .QN(\p[11][38] ) );
  NOR2X0 U1774 ( .IN1(n197), .IN2(n335), .QN(\p[14][38] ) );
  NOR2X0 U1775 ( .IN1(n193), .IN2(n335), .QN(\p[14][39] ) );
  NOR2X0 U1776 ( .IN1(n177), .IN2(n127), .QN(\p[11][40] ) );
  NOR2X0 U1777 ( .IN1(n189), .IN2(n335), .QN(\p[14][40] ) );
  NOR2X0 U1778 ( .IN1(n189), .IN2(n339), .QN(\p[12][38] ) );
  NOR2X0 U1779 ( .IN1(n185), .IN2(n339), .QN(\p[12][39] ) );
  NOR2X0 U1780 ( .IN1(n197), .IN2(n333), .QN(\p[15][39] ) );
  NOR2X0 U1781 ( .IN1(n181), .IN2(n339), .QN(\p[12][40] ) );
  NOR2X0 U1782 ( .IN1(n193), .IN2(n333), .QN(\p[15][40] ) );
  NOR2X0 U1783 ( .IN1(n189), .IN2(n332), .QN(\p[15][41] ) );
  NOR2X0 U1784 ( .IN1(n226), .IN2(n287), .QN(\p[30][46] ) );
  NOR2X0 U1785 ( .IN1(n196), .IN2(n329), .QN(\p[16][40] ) );
  NOR2X0 U1786 ( .IN1(n208), .IN2(n311), .QN(\p[22][43] ) );
  NOR2X0 U1787 ( .IN1(n223), .IN2(n293), .QN(\p[28][45] ) );
  NOR2X0 U1788 ( .IN1(n204), .IN2(n311), .QN(\p[22][44] ) );
  NOR2X0 U1789 ( .IN1(n215), .IN2(n302), .QN(\p[25][44] ) );
  NOR2X0 U1790 ( .IN1(n219), .IN2(n293), .QN(\p[28][46] ) );
  NOR2X0 U1791 ( .IN1(n200), .IN2(n311), .QN(\p[22][45] ) );
  NOR2X0 U1792 ( .IN1(n215), .IN2(n293), .QN(\p[28][47] ) );
  NOR2X0 U1793 ( .IN1(n230), .IN2(n287), .QN(\p[30][45] ) );
  NOR2X0 U1794 ( .IN1(n189), .IN2(n338), .QN(\p[13][39] ) );
  NOR2X0 U1795 ( .IN1(n185), .IN2(n338), .QN(\p[13][40] ) );
  NOR2X0 U1796 ( .IN1(n181), .IN2(n338), .QN(\p[13][41] ) );
  NOR2X0 U1797 ( .IN1(n173), .IN2(n342), .QN(\p[11][41] ) );
  NOR2X0 U1798 ( .IN1(n219), .IN2(n307), .QN(\p[23][41] ) );
  NOR2X0 U1799 ( .IN1(n211), .IN2(n299), .QN(\p[26][46] ) );
  NOR2X0 U1800 ( .IN1(n207), .IN2(n299), .QN(\p[26][47] ) );
  NOR2X0 U1801 ( .IN1(n211), .IN2(n290), .QN(\p[29][49] ) );
  NOR2X0 U1802 ( .IN1(n203), .IN2(n299), .QN(\p[26][48] ) );
  NOR2X0 U1803 ( .IN1(n214), .IN2(n287), .QN(\p[30][49] ) );
  NOR2X0 U1804 ( .IN1(n210), .IN2(n287), .QN(\p[30][50] ) );
  NOR2X0 U1805 ( .IN1(n207), .IN2(n296), .QN(\p[27][48] ) );
  NOR2X0 U1806 ( .IN1(n199), .IN2(n305), .QN(\p[24][47] ) );
  NOR2X0 U1807 ( .IN1(n203), .IN2(n296), .QN(\p[27][49] ) );
  NOR2X0 U1808 ( .IN1(n199), .IN2(n296), .QN(\p[27][50] ) );
  NOR2X0 U1809 ( .IN1(n192), .IN2(n327), .QN(\p[17][42] ) );
  NOR2X0 U1810 ( .IN1(n188), .IN2(n327), .QN(\p[17][43] ) );
  NOR2X0 U1811 ( .IN1(n196), .IN2(n318), .QN(\p[20][44] ) );
  NOR2X0 U1812 ( .IN1(n219), .IN2(n290), .QN(\p[29][47] ) );
  NOR2X0 U1813 ( .IN1(n215), .IN2(n290), .QN(\p[29][48] ) );
  NOR2X0 U1814 ( .IN1(n218), .IN2(n287), .QN(\p[30][48] ) );
  NOR2X0 U1815 ( .IN1(n196), .IN2(n324), .QN(\p[18][42] ) );
  NOR2X0 U1816 ( .IN1(n192), .IN2(n324), .QN(\p[18][43] ) );
  NOR2X0 U1817 ( .IN1(n188), .IN2(n324), .QN(\p[18][44] ) );
  NOR2X0 U1818 ( .IN1(n211), .IN2(n293), .QN(\p[28][48] ) );
  NOR2X0 U1819 ( .IN1(n203), .IN2(n302), .QN(\p[25][47] ) );
  NOR2X0 U1820 ( .IN1(n207), .IN2(n293), .QN(\p[28][49] ) );
  NOR2X0 U1821 ( .IN1(n199), .IN2(n302), .QN(\p[25][48] ) );
  NOR2X0 U1822 ( .IN1(n203), .IN2(n293), .QN(\p[28][50] ) );
  NOR2X0 U1823 ( .IN1(n185), .IN2(n335), .QN(\p[14][41] ) );
  NOR2X0 U1824 ( .IN1(n181), .IN2(n335), .QN(\p[14][42] ) );
  NOR2X0 U1825 ( .IN1(n177), .IN2(n335), .QN(\p[14][43] ) );
  NOR2X0 U1826 ( .IN1(n177), .IN2(n339), .QN(\p[12][41] ) );
  NOR2X0 U1827 ( .IN1(n173), .IN2(n339), .QN(\p[12][42] ) );
  NOR2X0 U1828 ( .IN1(n185), .IN2(n331), .QN(\p[15][42] ) );
  NOR2X0 U1829 ( .IN1(n181), .IN2(n331), .QN(\p[15][43] ) );
  NOR2X0 U1830 ( .IN1(n192), .IN2(n330), .QN(\p[16][41] ) );
  NOR2X0 U1831 ( .IN1(n188), .IN2(n329), .QN(\p[16][42] ) );
  NOR2X0 U1832 ( .IN1(n184), .IN2(n330), .QN(\p[16][43] ) );
  NOR2X0 U1833 ( .IN1(n196), .IN2(n321), .QN(\p[19][43] ) );
  NOR2X0 U1834 ( .IN1(n177), .IN2(n338), .QN(\p[13][42] ) );
  NOR2X0 U1835 ( .IN1(n173), .IN2(n338), .QN(\p[13][43] ) );
  NOR2X0 U1836 ( .IN1(n207), .IN2(n290), .QN(\p[29][50] ) );
  NOR2X0 U1837 ( .IN1(n199), .IN2(n299), .QN(\p[26][49] ) );
  NOR2X0 U1838 ( .IN1(n203), .IN2(n290), .QN(\p[29][51] ) );
  NOR2X0 U1839 ( .IN1(n199), .IN2(n290), .QN(\p[29][52] ) );
  NOR2X0 U1840 ( .IN1(n206), .IN2(n287), .QN(\p[30][51] ) );
  NOR2X0 U1841 ( .IN1(n202), .IN2(n287), .QN(\p[30][52] ) );
  NOR2X0 U1842 ( .IN1(n198), .IN2(n287), .QN(\p[30][53] ) );
  NOR2X0 U1843 ( .IN1(n195), .IN2(n306), .QN(\p[24][48] ) );
  NOR2X0 U1844 ( .IN1(n184), .IN2(n327), .QN(\p[17][44] ) );
  NOR2X0 U1845 ( .IN1(n180), .IN2(n327), .QN(\p[17][45] ) );
  NOR2X0 U1846 ( .IN1(n192), .IN2(n318), .QN(\p[20][45] ) );
  NOR2X0 U1847 ( .IN1(n176), .IN2(n327), .QN(\p[17][46] ) );
  NOR2X0 U1848 ( .IN1(n188), .IN2(n318), .QN(\p[20][46] ) );
  NOR2X0 U1849 ( .IN1(n184), .IN2(n318), .QN(\p[20][47] ) );
  NOR2X0 U1850 ( .IN1(n196), .IN2(n315), .QN(\p[21][45] ) );
  NOR2X0 U1851 ( .IN1(n184), .IN2(n324), .QN(\p[18][45] ) );
  NOR2X0 U1852 ( .IN1(n192), .IN2(n315), .QN(\p[21][46] ) );
  NOR2X0 U1853 ( .IN1(n180), .IN2(n324), .QN(\p[18][46] ) );
  NOR2X0 U1854 ( .IN1(n188), .IN2(n315), .QN(\p[21][47] ) );
  NOR2X0 U1855 ( .IN1(n176), .IN2(n324), .QN(\p[18][47] ) );
  NOR2X0 U1856 ( .IN1(n199), .IN2(n293), .QN(\p[28][51] ) );
  NOR2X0 U1857 ( .IN1(n173), .IN2(n335), .QN(\p[14][44] ) );
  NOR2X0 U1858 ( .IN1(n177), .IN2(n107), .QN(\p[15][44] ) );
  NOR2X0 U1859 ( .IN1(n173), .IN2(n332), .QN(\p[15][45] ) );
  NOR2X0 U1860 ( .IN1(n180), .IN2(n329), .QN(\p[16][44] ) );
  NOR2X0 U1861 ( .IN1(n192), .IN2(n321), .QN(\p[19][44] ) );
  NOR2X0 U1862 ( .IN1(n176), .IN2(n330), .QN(\p[16][45] ) );
  NOR2X0 U1863 ( .IN1(n188), .IN2(n321), .QN(\p[19][45] ) );
  NOR2X0 U1864 ( .IN1(n172), .IN2(n329), .QN(\p[16][46] ) );
  NOR2X0 U1865 ( .IN1(n196), .IN2(n312), .QN(\p[22][46] ) );
  NOR2X0 U1866 ( .IN1(n184), .IN2(n321), .QN(\p[19][46] ) );
  NOR2X0 U1867 ( .IN1(n192), .IN2(n312), .QN(\p[22][47] ) );
  NOR2X0 U1868 ( .IN1(n195), .IN2(n300), .QN(\p[26][50] ) );
  NOR2X0 U1869 ( .IN1(n191), .IN2(n306), .QN(\p[24][49] ) );
  NOR2X0 U1870 ( .IN1(n195), .IN2(n297), .QN(\p[27][51] ) );
  NOR2X0 U1871 ( .IN1(n187), .IN2(n306), .QN(\p[24][50] ) );
  NOR2X0 U1872 ( .IN1(n191), .IN2(n297), .QN(\p[27][52] ) );
  NOR2X0 U1873 ( .IN1(n183), .IN2(n306), .QN(\p[24][51] ) );
  NOR2X0 U1874 ( .IN1(n172), .IN2(n327), .QN(\p[17][47] ) );
  NOR2X0 U1875 ( .IN1(n180), .IN2(n318), .QN(\p[20][48] ) );
  NOR2X0 U1876 ( .IN1(n176), .IN2(n318), .QN(\p[20][49] ) );
  NOR2X0 U1877 ( .IN1(n172), .IN2(n318), .QN(\p[20][50] ) );
  NOR2X0 U1878 ( .IN1(n184), .IN2(n315), .QN(\p[21][48] ) );
  NOR2X0 U1879 ( .IN1(n172), .IN2(n324), .QN(\p[18][48] ) );
  NOR2X0 U1880 ( .IN1(n180), .IN2(n315), .QN(\p[21][49] ) );
  NOR2X0 U1881 ( .IN1(n176), .IN2(n315), .QN(\p[21][50] ) );
  NOR2X0 U1882 ( .IN1(n195), .IN2(n303), .QN(\p[25][49] ) );
  NOR2X0 U1883 ( .IN1(n191), .IN2(n303), .QN(\p[25][50] ) );
  NOR2X0 U1884 ( .IN1(n180), .IN2(n321), .QN(\p[19][47] ) );
  NOR2X0 U1885 ( .IN1(n188), .IN2(n312), .QN(\p[22][48] ) );
  NOR2X0 U1886 ( .IN1(n176), .IN2(n321), .QN(\p[19][48] ) );
  NOR2X0 U1887 ( .IN1(n184), .IN2(n312), .QN(\p[22][49] ) );
  NOR2X0 U1888 ( .IN1(n172), .IN2(n321), .QN(\p[19][49] ) );
  NOR2X0 U1889 ( .IN1(n180), .IN2(n312), .QN(\p[22][50] ) );
  NOR2X0 U1890 ( .IN1(n191), .IN2(n300), .QN(\p[26][51] ) );
  NOR2X0 U1891 ( .IN1(n195), .IN2(n291), .QN(\p[29][53] ) );
  NOR2X0 U1892 ( .IN1(n187), .IN2(n300), .QN(\p[26][52] ) );
  NOR2X0 U1893 ( .IN1(n191), .IN2(n291), .QN(\p[29][54] ) );
  NOR2X0 U1894 ( .IN1(n183), .IN2(n300), .QN(\p[26][53] ) );
  NOR2X0 U1895 ( .IN1(n187), .IN2(n297), .QN(\p[27][53] ) );
  NOR2X0 U1896 ( .IN1(n179), .IN2(n306), .QN(\p[24][52] ) );
  NOR2X0 U1897 ( .IN1(n183), .IN2(n297), .QN(\p[27][54] ) );
  NOR2X0 U1898 ( .IN1(n175), .IN2(n306), .QN(\p[24][53] ) );
  NOR2X0 U1899 ( .IN1(n179), .IN2(n297), .QN(\p[27][55] ) );
  NOR2X0 U1900 ( .IN1(n171), .IN2(n306), .QN(\p[24][54] ) );
  NOR2X0 U1901 ( .IN1(n194), .IN2(n288), .QN(\p[30][54] ) );
  NOR2X0 U1902 ( .IN1(n172), .IN2(n315), .QN(\p[21][51] ) );
  NOR2X0 U1903 ( .IN1(n195), .IN2(n294), .QN(\p[28][52] ) );
  NOR2X0 U1904 ( .IN1(n187), .IN2(n303), .QN(\p[25][51] ) );
  NOR2X0 U1905 ( .IN1(n191), .IN2(n294), .QN(\p[28][53] ) );
  NOR2X0 U1906 ( .IN1(n183), .IN2(n303), .QN(\p[25][52] ) );
  NOR2X0 U1907 ( .IN1(n187), .IN2(n294), .QN(\p[28][54] ) );
  NOR2X0 U1908 ( .IN1(n179), .IN2(n303), .QN(\p[25][53] ) );
  NOR2X0 U1909 ( .IN1(n176), .IN2(n312), .QN(\p[22][51] ) );
  NOR2X0 U1910 ( .IN1(n172), .IN2(n312), .QN(\p[22][52] ) );
  NOR2X0 U1911 ( .IN1(n187), .IN2(n291), .QN(\p[29][55] ) );
  NOR2X0 U1912 ( .IN1(n179), .IN2(n300), .QN(\p[26][54] ) );
  NOR2X0 U1913 ( .IN1(n183), .IN2(n291), .QN(\p[29][56] ) );
  NOR2X0 U1914 ( .IN1(n175), .IN2(n300), .QN(\p[26][55] ) );
  NOR2X0 U1915 ( .IN1(n179), .IN2(n291), .QN(\p[29][57] ) );
  NOR2X0 U1916 ( .IN1(n171), .IN2(n300), .QN(\p[26][56] ) );
  NOR2X0 U1917 ( .IN1(n175), .IN2(n297), .QN(\p[27][56] ) );
  NOR2X0 U1918 ( .IN1(n171), .IN2(n297), .QN(\p[27][57] ) );
  NOR2X0 U1919 ( .IN1(n190), .IN2(n288), .QN(\p[30][55] ) );
  NOR2X0 U1920 ( .IN1(n186), .IN2(n288), .QN(\p[30][56] ) );
  NOR2X0 U1921 ( .IN1(n182), .IN2(n288), .QN(\p[30][57] ) );
  NOR2X0 U1922 ( .IN1(n183), .IN2(n294), .QN(\p[28][55] ) );
  NOR2X0 U1923 ( .IN1(n175), .IN2(n303), .QN(\p[25][54] ) );
  NOR2X0 U1924 ( .IN1(n179), .IN2(n294), .QN(\p[28][56] ) );
  NOR2X0 U1925 ( .IN1(n171), .IN2(n303), .QN(\p[25][55] ) );
  NOR2X0 U1926 ( .IN1(n175), .IN2(n294), .QN(\p[28][57] ) );
  NOR2X0 U1927 ( .IN1(n175), .IN2(n291), .QN(\p[29][58] ) );
  NOR2X0 U1928 ( .IN1(n171), .IN2(n291), .QN(\p[29][59] ) );
  NOR2X0 U1929 ( .IN1(n178), .IN2(n288), .QN(\p[30][58] ) );
  NOR2X0 U1930 ( .IN1(n171), .IN2(n294), .QN(\p[28][58] ) );
  NOR2X0 U1931 ( .IN1(n174), .IN2(n288), .QN(\p[30][59] ) );
  NOR2X0 U1932 ( .IN1(n170), .IN2(n288), .QN(\p[30][60] ) );
  NBUFFX2 U1933 ( .INP(\p[58][63] ), .Z(n477) );
  DELLN1X2 U1934 ( .INP(n143), .Z(n361) );
  NOR2X0 U1935 ( .IN1(n348), .IN2(n112), .QN(\p[9][17] ) );
  DELLN1X2 U1936 ( .INP(n553), .Z(n278) );
  DELLN1X2 U1937 ( .INP(n549), .Z(n265) );
  DELLN1X2 U1938 ( .INP(n549), .Z(n266) );
  DELLN1X2 U1939 ( .INP(n550), .Z(n271) );
  DELLN1X2 U1940 ( .INP(n549), .Z(n267) );
  NBUFFX2 U1941 ( .INP(n76), .Z(n210) );
  NBUFFX2 U1942 ( .INP(n75), .Z(n214) );
  NBUFFX2 U1943 ( .INP(n74), .Z(n207) );
  NBUFFX2 U1944 ( .INP(n76), .Z(n211) );
  NBUFFX2 U1945 ( .INP(n77), .Z(n218) );
  NBUFFX2 U1946 ( .INP(n79), .Z(n231) );
  NBUFFX2 U1947 ( .INP(n78), .Z(n222) );
  NBUFFX2 U1948 ( .INP(n79), .Z(n230) );
  NOR2X0 U1949 ( .IN1(n348), .IN2(n244), .QN(\p[9][21] ) );
  NBUFFX4 U1950 ( .INP(n98), .Z(n289) );
  NBUFFX2 U1951 ( .INP(n557), .Z(n349) );
  NBUFFX2 U1952 ( .INP(n557), .Z(n347) );
  NBUFFX2 U1953 ( .INP(n74), .Z(n206) );
  NBUFFX2 U1954 ( .INP(n73), .Z(n202) );
  NBUFFX2 U1955 ( .INP(n90), .Z(n198) );
  NBUFFX2 U1956 ( .INP(n73), .Z(n203) );
  NBUFFX2 U1957 ( .INP(n90), .Z(n199) );
  NBUFFX2 U1958 ( .INP(n96), .Z(n195) );
  NBUFFX2 U1959 ( .INP(n75), .Z(n216) );
  NBUFFX2 U1960 ( .INP(n78), .Z(n223) );
  NBUFFX2 U1961 ( .INP(n77), .Z(n219) );
  NBUFFX2 U1962 ( .INP(n75), .Z(n215) );
  NBUFFX4 U1963 ( .INP(n86), .Z(n323) );
  NBUFFX4 U1964 ( .INP(n87), .Z(n326) );
  NBUFFX4 U1965 ( .INP(n104), .Z(n286) );
  NBUFFX2 U1966 ( .INP(n121), .Z(n250) );
  DELLN1X2 U1967 ( .INP(n121), .Z(n253) );
  NBUFFX2 U1968 ( .INP(n95), .Z(n191) );
  NBUFFX2 U1969 ( .INP(n94), .Z(n187) );
  NBUFFX2 U1970 ( .INP(n93), .Z(n183) );
  NBUFFX2 U1971 ( .INP(n95), .Z(n190) );
  NBUFFX2 U1972 ( .INP(n96), .Z(n194) );
  NBUFFX2 U1973 ( .INP(n94), .Z(n186) );
  NBUFFX2 U1974 ( .INP(n73), .Z(n204) );
  NBUFFX2 U1975 ( .INP(n90), .Z(n200) );
  NBUFFX2 U1976 ( .INP(n96), .Z(n196) );
  NBUFFX2 U1977 ( .INP(n95), .Z(n193) );
  NBUFFX2 U1978 ( .INP(n96), .Z(n197) );
  NBUFFX4 U1979 ( .INP(n85), .Z(n317) );
  NBUFFX4 U1980 ( .INP(n84), .Z(n314) );
  NOR2X0 U1981 ( .IN1(n221), .IN2(n344), .QN(\p[10][28] ) );
  NBUFFX2 U1982 ( .INP(n556), .Z(n308) );
  NBUFFX2 U1983 ( .INP(n556), .Z(n307) );
  NBUFFX2 U1984 ( .INP(n556), .Z(n309) );
  NBUFFX2 U1985 ( .INP(\p[61][63] ), .Z(n489) );
  NBUFFX2 U1986 ( .INP(\p[63][63] ), .Z(n501) );
  NBUFFX2 U1987 ( .INP(\p[62][63] ), .Z(n496) );
  NBUFFX4 U1988 ( .INP(\p[63][63] ), .Z(n498) );
  NBUFFX2 U1989 ( .INP(\p[62][63] ), .Z(n493) );
  NBUFFX2 U1990 ( .INP(\p[61][63] ), .Z(n488) );
  NBUFFX2 U1991 ( .INP(\p[3][63] ), .Z(n518) );
  NBUFFX2 U1992 ( .INP(\p[62][63] ), .Z(n497) );
  NBUFFX2 U1993 ( .INP(n92), .Z(n179) );
  NBUFFX2 U1994 ( .INP(n97), .Z(n175) );
  NBUFFX2 U1995 ( .INP(n103), .Z(n171) );
  NBUFFX2 U1996 ( .INP(n93), .Z(n182) );
  NBUFFX2 U1997 ( .INP(n92), .Z(n178) );
  NBUFFX2 U1998 ( .INP(n95), .Z(n192) );
  NBUFFX2 U1999 ( .INP(n94), .Z(n188) );
  NBUFFX2 U2000 ( .INP(n92), .Z(n180) );
  NBUFFX2 U2001 ( .INP(n93), .Z(n184) );
  NBUFFX2 U2002 ( .INP(n97), .Z(n176) );
  NBUFFX2 U2003 ( .INP(n103), .Z(n172) );
  NBUFFX2 U2004 ( .INP(n97), .Z(n174) );
  NBUFFX2 U2005 ( .INP(n94), .Z(n189) );
  NBUFFX2 U2006 ( .INP(n93), .Z(n185) );
  NBUFFX2 U2007 ( .INP(n97), .Z(n177) );
  NBUFFX2 U2008 ( .INP(n92), .Z(n181) );
  NBUFFX2 U2009 ( .INP(n103), .Z(n173) );
  NBUFFX2 U2010 ( .INP(n103), .Z(n170) );
  NOR2X0 U2011 ( .IN1(n265), .IN2(n122), .QN(\p[23][29] ) );
  NOR2X0 U2012 ( .IN1(n170), .IN2(n362), .QN(\p[3][33] ) );
  NOR2X0 U2013 ( .IN1(n178), .IN2(n362), .QN(\p[3][31] ) );
  NOR2X0 U2014 ( .IN1(n174), .IN2(n362), .QN(\p[3][32] ) );
  NOR2X0 U2015 ( .IN1(n171), .IN2(n365), .QN(\p[2][32] ) );
  NBUFFX4 U2016 ( .INP(n83), .Z(n311) );
  NBUFFX4 U2017 ( .INP(n99), .Z(n296) );
  NOR2X0 U2018 ( .IN1(n275), .IN2(n122), .QN(\p[23][26] ) );
  NOR2X0 U2019 ( .IN1(n262), .IN2(n122), .QN(\p[23][30] ) );
  NOR2X0 U2020 ( .IN1(n137), .IN2(n122), .QN(\p[23][28] ) );
  NOR2X0 U2021 ( .IN1(n549), .IN2(n286), .QN(\p[30][36] ) );
  AND2X1 U2022 ( .IN1(n540), .IN2(A_reg[5]), .Q(\p[58][63] ) );
  NBUFFX2 U2023 ( .INP(\p[59][63] ), .Z(n479) );
  NBUFFX2 U2024 ( .INP(\p[60][63] ), .Z(n486) );
  NBUFFX2 U2025 ( .INP(\p[56][63] ), .Z(n463) );
  NBUFFX2 U2026 ( .INP(\p[5][63] ), .Z(n526) );
  NBUFFX2 U2027 ( .INP(\p[60][63] ), .Z(n483) );
  NBUFFX2 U2028 ( .INP(\p[59][63] ), .Z(n478) );
  NBUFFX2 U2029 ( .INP(\p[6][63] ), .Z(n531) );
  NBUFFX2 U2030 ( .INP(\p[60][63] ), .Z(n485) );
  NBUFFX2 U2031 ( .INP(\p[0][63] ), .Z(n504) );
  NBUFFX2 U2032 ( .INP(\p[2][63] ), .Z(n515) );
  NBUFFX2 U2033 ( .INP(\p[60][63] ), .Z(n487) );
  NOR2X0 U2034 ( .IN1(n170), .IN2(n131), .QN(\p[6][36] ) );
  NBUFFX4 U2035 ( .INP(\p[14][63] ), .Z(n395) );
  NOR2X0 U2036 ( .IN1(n211), .IN2(n556), .QN(\p[23][43] ) );
  NBUFFX2 U2037 ( .INP(\p[57][63] ), .Z(n466) );
  NBUFFX2 U2038 ( .INP(\p[57][63] ), .Z(n467) );
  NBUFFX2 U2039 ( .INP(\p[57][63] ), .Z(n472) );
  NBUFFX2 U2040 ( .INP(\p[54][63] ), .Z(n454) );
  NBUFFX2 U2041 ( .INP(\p[60][63] ), .Z(n484) );
  NBUFFX2 U2042 ( .INP(\p[55][63] ), .Z(n457) );
  NBUFFX2 U2043 ( .INP(\p[56][63] ), .Z(n461) );
  NBUFFX2 U2044 ( .INP(\p[7][63] ), .Z(n536) );
  NBUFFX2 U2045 ( .INP(\p[59][63] ), .Z(n481) );
  NBUFFX2 U2046 ( .INP(\p[1][63] ), .Z(n510) );
  NBUFFX2 U2047 ( .INP(\p[10][63] ), .Z(n380) );
  NBUFFX2 U2048 ( .INP(\p[56][63] ), .Z(n460) );
  NBUFFX2 U2049 ( .INP(\p[8][63] ), .Z(n372) );
  NBUFFX2 U2050 ( .INP(\p[3][63] ), .Z(n519) );
  NBUFFX2 U2051 ( .INP(\p[9][63] ), .Z(n376) );
  NBUFFX2 U2052 ( .INP(\p[62][63] ), .Z(n495) );
  NBUFFX2 U2053 ( .INP(\p[61][63] ), .Z(n490) );
  NBUFFX2 U2054 ( .INP(\p[55][63] ), .Z(n458) );
  NBUFFX2 U2055 ( .INP(\p[61][63] ), .Z(n492) );
  NBUFFX2 U2056 ( .INP(\p[59][63] ), .Z(n482) );
  NBUFFX2 U2057 ( .INP(n87), .Z(n327) );
  NOR2X0 U2058 ( .IN1(n207), .IN2(n556), .QN(\p[23][44] ) );
  NOR2X0 U2059 ( .IN1(n203), .IN2(n556), .QN(\p[23][45] ) );
  NOR2X0 U2060 ( .IN1(n199), .IN2(n556), .QN(\p[23][46] ) );
  NBUFFX2 U2061 ( .INP(\p[57][63] ), .Z(n464) );
  NBUFFX2 U2062 ( .INP(\p[57][63] ), .Z(n471) );
  NBUFFX2 U2063 ( .INP(\p[54][63] ), .Z(n453) );
  NBUFFX2 U2064 ( .INP(\p[63][63] ), .Z(n499) );
  NBUFFX2 U2065 ( .INP(\p[53][63] ), .Z(n449) );
  NBUFFX2 U2066 ( .INP(\p[13][63] ), .Z(n392) );
  NBUFFX2 U2067 ( .INP(\p[11][63] ), .Z(n384) );
  NBUFFX2 U2068 ( .INP(\p[5][63] ), .Z(n527) );
  NBUFFX2 U2069 ( .INP(\p[12][63] ), .Z(n388) );
  NBUFFX2 U2070 ( .INP(\p[63][63] ), .Z(n500) );
  NBUFFX2 U2071 ( .INP(\p[0][63] ), .Z(n505) );
  NBUFFX2 U2072 ( .INP(\p[59][63] ), .Z(n480) );
  NBUFFX2 U2073 ( .INP(n86), .Z(n324) );
  NBUFFX2 U2074 ( .INP(n85), .Z(n318) );
  NOR2X0 U2075 ( .IN1(n195), .IN2(n556), .QN(\p[23][47] ) );
  NOR2X0 U2076 ( .IN1(n191), .IN2(n556), .QN(\p[23][48] ) );
  NOR2X0 U2077 ( .IN1(n187), .IN2(n556), .QN(\p[23][49] ) );
  NBUFFX2 U2078 ( .INP(\p[57][63] ), .Z(n470) );
  NBUFFX2 U2079 ( .INP(\p[51][63] ), .Z(n438) );
  NBUFFX2 U2080 ( .INP(\p[51][63] ), .Z(n439) );
  NBUFFX2 U2081 ( .INP(\p[51][63] ), .Z(n443) );
  NBUFFX2 U2082 ( .INP(\p[52][63] ), .Z(n445) );
  NBUFFX2 U2083 ( .INP(\p[52][63] ), .Z(n446) );
  NBUFFX2 U2084 ( .INP(\p[62][63] ), .Z(n494) );
  NBUFFX2 U2085 ( .INP(\p[50][63] ), .Z(n435) );
  NBUFFX2 U2086 ( .INP(\p[50][63] ), .Z(n436) );
  NBUFFX2 U2087 ( .INP(\p[7][63] ), .Z(n537) );
  NBUFFX2 U2088 ( .INP(\p[1][63] ), .Z(n511) );
  NBUFFX2 U2089 ( .INP(\p[50][63] ), .Z(n434) );
  NBUFFX2 U2090 ( .INP(\p[52][63] ), .Z(n444) );
  NBUFFX2 U2091 ( .INP(\p[55][63] ), .Z(n456) );
  NBUFFX2 U2092 ( .INP(\p[54][63] ), .Z(n452) );
  NBUFFX2 U2093 ( .INP(\p[53][63] ), .Z(n448) );
  NBUFFX2 U2094 ( .INP(\p[8][63] ), .Z(n373) );
  NBUFFX2 U2095 ( .INP(\p[15][63] ), .Z(n397) );
  NBUFFX2 U2096 ( .INP(\p[6][63] ), .Z(n532) );
  NBUFFX2 U2097 ( .INP(\p[3][63] ), .Z(n520) );
  NBUFFX2 U2098 ( .INP(\p[49][63] ), .Z(n433) );
  NBUFFX2 U2099 ( .INP(\p[55][63] ), .Z(n459) );
  NBUFFX2 U2100 ( .INP(\p[2][63] ), .Z(n516) );
  NBUFFX2 U2101 ( .INP(\p[53][63] ), .Z(n451) );
  NBUFFX2 U2102 ( .INP(\p[52][63] ), .Z(n447) );
  NBUFFX2 U2103 ( .INP(n84), .Z(n315) );
  NBUFFX2 U2104 ( .INP(n83), .Z(n312) );
  NBUFFX2 U2105 ( .INP(n100), .Z(n306) );
  NBUFFX2 U2106 ( .INP(\p[42][63] ), .Z(n156) );
  NBUFFX2 U2107 ( .INP(\p[42][63] ), .Z(n158) );
  NBUFFX2 U2108 ( .INP(\p[21][63] ), .Z(n153) );
  NBUFFX2 U2109 ( .INP(\p[42][63] ), .Z(n157) );
  NOR2X0 U2110 ( .IN1(n183), .IN2(n556), .QN(\p[23][50] ) );
  NOR2X0 U2111 ( .IN1(n179), .IN2(n556), .QN(\p[23][51] ) );
  NOR2X0 U2112 ( .IN1(n175), .IN2(n556), .QN(\p[23][52] ) );
  NBUFFX2 U2113 ( .INP(\p[57][63] ), .Z(n465) );
  NBUFFX2 U2114 ( .INP(\p[51][63] ), .Z(n437) );
  NBUFFX2 U2115 ( .INP(\p[57][63] ), .Z(n468) );
  NBUFFX2 U2116 ( .INP(\p[51][63] ), .Z(n442) );
  NBUFFX2 U2117 ( .INP(\p[49][63] ), .Z(n432) );
  NBUFFX2 U2118 ( .INP(\p[47][63] ), .Z(n425) );
  NBUFFX2 U2119 ( .INP(\p[53][63] ), .Z(n450) );
  NBUFFX2 U2120 ( .INP(\p[48][63] ), .Z(n429) );
  NBUFFX2 U2121 ( .INP(\p[16][63] ), .Z(n400) );
  NBUFFX2 U2122 ( .INP(\p[10][63] ), .Z(n381) );
  NBUFFX2 U2123 ( .INP(\p[17][63] ), .Z(n403) );
  NBUFFX2 U2124 ( .INP(\p[49][63] ), .Z(n431) );
  NBUFFX2 U2125 ( .INP(\p[48][63] ), .Z(n428) );
  NBUFFX2 U2126 ( .INP(\p[11][63] ), .Z(n385) );
  NBUFFX2 U2127 ( .INP(\p[5][63] ), .Z(n528) );
  NBUFFX2 U2128 ( .INP(\p[18][63] ), .Z(n406) );
  NBUFFX2 U2129 ( .INP(\p[12][63] ), .Z(n389) );
  NBUFFX2 U2130 ( .INP(\p[9][63] ), .Z(n377) );
  NBUFFX2 U2131 ( .INP(\p[0][63] ), .Z(n506) );
  NBUFFX2 U2132 ( .INP(\p[56][63] ), .Z(n462) );
  NBUFFX2 U2133 ( .INP(\p[20][63] ), .Z(n411) );
  NBUFFX2 U2134 ( .INP(\p[48][63] ), .Z(n430) );
  NBUFFX2 U2135 ( .INP(n102), .Z(n303) );
  NBUFFX2 U2136 ( .INP(n99), .Z(n297) );
  NBUFFX2 U2137 ( .INP(n101), .Z(n300) );
  NBUFFX2 U2138 ( .INP(\p[21][63] ), .Z(n155) );
  NBUFFX2 U2139 ( .INP(\p[21][63] ), .Z(n154) );
  NOR2X0 U2140 ( .IN1(n171), .IN2(n556), .QN(\p[23][53] ) );
  NBUFFX2 U2141 ( .INP(\p[45][63] ), .Z(n418) );
  NBUFFX2 U2142 ( .INP(\p[51][63] ), .Z(n440) );
  NBUFFX2 U2143 ( .INP(\p[45][63] ), .Z(n421) );
  NBUFFX2 U2144 ( .INP(\p[43][63] ), .Z(n413) );
  NBUFFX2 U2145 ( .INP(\p[44][63] ), .Z(n416) );
  NBUFFX2 U2146 ( .INP(\p[44][63] ), .Z(n415) );
  NBUFFX2 U2147 ( .INP(\p[46][63] ), .Z(n423) );
  NBUFFX2 U2148 ( .INP(\p[19][63] ), .Z(n409) );
  NBUFFX2 U2149 ( .INP(\p[13][63] ), .Z(n393) );
  NBUFFX2 U2150 ( .INP(\p[1][63] ), .Z(n512) );
  NBUFFX2 U2151 ( .INP(\p[46][63] ), .Z(n422) );
  NBUFFX2 U2152 ( .INP(\p[6][63] ), .Z(n533) );
  NBUFFX2 U2153 ( .INP(\p[47][63] ), .Z(n426) );
  NBUFFX2 U2154 ( .INP(\p[43][63] ), .Z(n414) );
  NBUFFX2 U2155 ( .INP(\p[47][63] ), .Z(n427) );
  NBUFFX2 U2156 ( .INP(\p[46][63] ), .Z(n424) );
  NBUFFX2 U2157 ( .INP(n91), .Z(n294) );
  NBUFFX2 U2158 ( .INP(n98), .Z(n291) );
  NBUFFX2 U2159 ( .INP(n104), .Z(n288) );
  NBUFFX2 U2160 ( .INP(\p[51][63] ), .Z(n441) );
  NBUFFX2 U2161 ( .INP(\p[45][63] ), .Z(n417) );
  NBUFFX2 U2162 ( .INP(\p[45][63] ), .Z(n419) );
  NBUFFX2 U2163 ( .INP(\p[57][63] ), .Z(n469) );
  NBUFFX2 U2164 ( .INP(\p[16][63] ), .Z(n401) );
  NBUFFX2 U2165 ( .INP(\p[7][63] ), .Z(n538) );
  NBUFFX2 U2166 ( .INP(\p[10][63] ), .Z(n382) );
  NBUFFX2 U2167 ( .INP(\p[17][63] ), .Z(n404) );
  NBUFFX2 U2168 ( .INP(\p[11][63] ), .Z(n386) );
  NBUFFX2 U2169 ( .INP(\p[8][63] ), .Z(n374) );
  NBUFFX2 U2170 ( .INP(\p[5][63] ), .Z(n529) );
  NBUFFX2 U2171 ( .INP(\p[15][63] ), .Z(n398) );
  NBUFFX2 U2172 ( .INP(\p[18][63] ), .Z(n407) );
  NBUFFX2 U2173 ( .INP(\p[12][63] ), .Z(n390) );
  NBUFFX2 U2174 ( .INP(\p[3][63] ), .Z(n521) );
  NBUFFX2 U2175 ( .INP(\p[9][63] ), .Z(n378) );
  NBUFFX2 U2176 ( .INP(\p[0][63] ), .Z(n507) );
  NBUFFX2 U2177 ( .INP(\p[4][63] ), .Z(n525) );
  NBUFFX2 U2178 ( .INP(\p[14][63] ), .Z(n396) );
  NBUFFX2 U2179 ( .INP(\p[45][63] ), .Z(n420) );
  NBUFFX2 U2180 ( .INP(\p[19][63] ), .Z(n410) );
  NBUFFX2 U2181 ( .INP(\p[6][63] ), .Z(n534) );
  NBUFFX2 U2182 ( .INP(\p[2][63] ), .Z(n517) );
  NBUFFX2 U2183 ( .INP(\p[54][63] ), .Z(n455) );
  NBUFFX2 U2184 ( .INP(\p[8][63] ), .Z(n375) );
  NBUFFX2 U2185 ( .INP(\p[15][63] ), .Z(n399) );
  NBUFFX2 U2186 ( .INP(\p[3][63] ), .Z(n522) );
  NBUFFX2 U2187 ( .INP(\p[9][63] ), .Z(n379) );
  NBUFFX2 U2188 ( .INP(\p[13][63] ), .Z(n394) );
  NBUFFX2 U2189 ( .INP(\p[7][63] ), .Z(n539) );
  NBUFFX2 U2190 ( .INP(\p[5][63] ), .Z(n530) );
  NBUFFX2 U2191 ( .INP(\p[11][63] ), .Z(n387) );
  NBUFFX2 U2192 ( .INP(\p[17][63] ), .Z(n405) );
  NBUFFX2 U2193 ( .INP(\p[1][63] ), .Z(n513) );
  NBUFFX2 U2194 ( .INP(\p[0][63] ), .Z(n508) );
  NBUFFX2 U2195 ( .INP(\p[20][63] ), .Z(n412) );
  NBUFFX2 U2196 ( .INP(\p[6][63] ), .Z(n535) );
  NBUFFX2 U2197 ( .INP(\p[12][63] ), .Z(n391) );
  NBUFFX2 U2198 ( .INP(\p[18][63] ), .Z(n408) );
  NBUFFX2 U2199 ( .INP(\p[16][63] ), .Z(n402) );
  NBUFFX2 U2200 ( .INP(\p[10][63] ), .Z(n383) );
  NBUFFX2 U2201 ( .INP(n546), .Z(n168) );
  NBUFFX2 U2202 ( .INP(n546), .Z(n167) );
  NBUFFX2 U2203 ( .INP(n546), .Z(n166) );
  NBUFFX2 U2204 ( .INP(n546), .Z(n165) );
  NBUFFX2 U2205 ( .INP(n546), .Z(n160) );
  NBUFFX2 U2206 ( .INP(n546), .Z(n159) );
  NBUFFX2 U2207 ( .INP(n546), .Z(n164) );
  NBUFFX2 U2208 ( .INP(n546), .Z(n163) );
  NBUFFX2 U2209 ( .INP(n546), .Z(n162) );
  NBUFFX2 U2210 ( .INP(n546), .Z(n161) );
  NBUFFX2 U2211 ( .INP(n546), .Z(n169) );
  NOR2X0 U2212 ( .IN1(n123), .IN2(n248), .QN(\p[9][20] ) );
  NOR2X0 U2213 ( .IN1(n123), .IN2(n148), .QN(\p[9][15] ) );
  NOR2X0 U2214 ( .IN1(n120), .IN2(n363), .QN(\p[3][3] ) );
  NOR2X0 U2215 ( .IN1(n123), .IN2(n152), .QN(\p[9][16] ) );
  NOR2X0 U2216 ( .IN1(n214), .IN2(n359), .QN(\p[4][23] ) );
  NOR2X0 U2217 ( .IN1(n123), .IN2(n119), .QN(\p[9][18] ) );
  NOR2X0 U2218 ( .IN1(n123), .IN2(n121), .QN(\p[9][19] ) );
  NOR2X0 U2219 ( .IN1(n281), .IN2(n122), .QN(\p[23][24] ) );
  NOR2X0 U2220 ( .IN1(n284), .IN2(n122), .QN(\p[23][23] ) );
  NOR2X0 U2221 ( .IN1(n277), .IN2(n122), .QN(\p[23][25] ) );
  NOR2X0 U2222 ( .IN1(n243), .IN2(n127), .QN(\p[11][23] ) );
  NOR2X0 U2223 ( .IN1(n241), .IN2(n127), .QN(\p[11][24] ) );
  NOR2X0 U2224 ( .IN1(n229), .IN2(n345), .QN(\p[10][26] ) );
  NOR2X0 U2225 ( .IN1(n225), .IN2(n345), .QN(\p[10][27] ) );
  NBUFFX2 U2226 ( .INP(A_reg[31]), .Z(n545) );
  NOR2X0 U2227 ( .IN1(n202), .IN2(n126), .QN(\p[8][30] ) );
  NOR2X0 U2228 ( .IN1(n206), .IN2(n126), .QN(\p[8][29] ) );
  NOR2X0 U2229 ( .IN1(n186), .IN2(n126), .QN(\p[8][34] ) );
  NOR2X0 U2230 ( .IN1(n217), .IN2(n345), .QN(\p[10][29] ) );
  AND2X1 U2231 ( .IN1(B_reg[4]), .IN2(n545), .Q(\p[4][63] ) );
  AND2X1 U2232 ( .IN1(B_reg[1]), .IN2(n543), .Q(\p[1][63] ) );
  AND2X1 U2233 ( .IN1(n540), .IN2(A_reg[2]), .Q(\p[61][63] ) );
  NOR2X0 U2234 ( .IN1(n178), .IN2(n126), .QN(\p[8][36] ) );
  AND2X1 U2235 ( .IN1(n540), .IN2(A_reg[6]), .Q(\p[57][63] ) );
  AND2X1 U2236 ( .IN1(B_reg[10]), .IN2(n543), .Q(\p[10][63] ) );
  AND2X1 U2237 ( .IN1(n545), .IN2(B_reg[9]), .Q(\p[9][63] ) );
  NBUFFX2 U2238 ( .INP(B_reg[31]), .Z(n541) );
  AND2X1 U2239 ( .IN1(n541), .IN2(A_reg[21]), .Q(\p[42][63] ) );
  AND2X1 U2240 ( .IN1(B_reg[21]), .IN2(n544), .Q(\p[21][63] ) );
  AND2X1 U2241 ( .IN1(n541), .IN2(A_reg[22]), .Q(\p[41][63] ) );
  AND2X1 U2242 ( .IN1(B_reg[22]), .IN2(n544), .Q(\p[22][63] ) );
  AND2X1 U2243 ( .IN1(B_reg[23]), .IN2(n544), .Q(\p[23][63] ) );
  AND2X1 U2244 ( .IN1(n541), .IN2(A_reg[23]), .Q(\p[40][63] ) );
  AND2X1 U2245 ( .IN1(B_reg[24]), .IN2(n544), .Q(\p[24][63] ) );
  AND2X1 U2246 ( .IN1(n542), .IN2(A_reg[24]), .Q(\p[39][63] ) );
  NBUFFX2 U2247 ( .INP(B_reg[31]), .Z(n542) );
  INVX0 U2248 ( .INP(rst), .ZN(n546) );
  DELLN1X2 U2249 ( .INP(n547), .Z(n255) );
  DELLN1X2 U2250 ( .INP(n555), .Z(n284) );
  DELLN1X2 U2251 ( .INP(n121), .Z(n252) );
  DELLN1X2 U2252 ( .INP(n121), .Z(n251) );
  INVX0 U2253 ( .INP(B_reg[23]), .ZN(n556) );
  NOR2X0 U2254 ( .IN1(n246), .IN2(n325), .QN(\p[17][28] ) );
  NOR2X0 U2255 ( .IN1(n250), .IN2(n325), .QN(\p[17][27] ) );
  NOR2X0 U2256 ( .IN1(n255), .IN2(n325), .QN(\p[17][26] ) );
  NOR2X0 U2257 ( .IN1(n261), .IN2(n325), .QN(\p[17][24] ) );
  NOR2X0 U2258 ( .IN1(n282), .IN2(n325), .QN(\p[17][18] ) );
  DELLN1X2 U2259 ( .INP(n558), .Z(n350) );
  NOR2X0 U2260 ( .IN1(n247), .IN2(n322), .QN(\p[18][29] ) );
  NOR2X0 U2261 ( .IN1(n250), .IN2(n322), .QN(\p[18][28] ) );
  NOR2X0 U2262 ( .IN1(n255), .IN2(n322), .QN(\p[18][27] ) );
  NOR2X0 U2263 ( .IN1(n151), .IN2(n322), .QN(\p[18][25] ) );
  NOR2X0 U2264 ( .IN1(n554), .IN2(n322), .QN(\p[18][19] ) );
  DELLN1X2 U2265 ( .INP(n554), .Z(n282) );
  DELLN1X2 U2266 ( .INP(n562), .Z(n135) );
  DELLN1X2 U2267 ( .INP(n550), .Z(n137) );
  DELLN1X2 U2268 ( .INP(n141), .Z(n140) );
  DELLN1X2 U2269 ( .INP(n109), .Z(n144) );
  DELLN1X2 U2270 ( .INP(n145), .Z(n363) );
  NOR2X0 U2271 ( .IN1(n284), .IN2(n310), .QN(\p[22][22] ) );
  DELLN1X2 U2272 ( .INP(n83), .Z(n310) );
  NOR2X0 U2273 ( .IN1(n557), .IN2(n271), .QN(\p[9][14] ) );
  NOR2X0 U2274 ( .IN1(n114), .IN2(n289), .QN(\p[29][33] ) );
  NOR2X0 U2275 ( .IN1(n114), .IN2(n298), .QN(\p[26][30] ) );
  NOR2X0 U2276 ( .IN1(n114), .IN2(n301), .QN(\p[25][29] ) );
  NOR2X0 U2277 ( .IN1(n273), .IN2(n122), .QN(\p[23][27] ) );
  NOR2X0 U2278 ( .IN1(n557), .IN2(n272), .QN(\p[9][13] ) );
  DELLN1X2 U2279 ( .INP(n72), .Z(n345) );
  DELLN1X2 U2280 ( .INP(n564), .Z(n369) );
  NOR2X0 U2281 ( .IN1(n284), .IN2(n313), .QN(\p[21][21] ) );
  DELLN1X2 U2282 ( .INP(n84), .Z(n313) );
  NOR2X0 U2283 ( .IN1(n270), .IN2(n310), .QN(\p[22][27] ) );
  NOR2X0 U2284 ( .IN1(n268), .IN2(n313), .QN(\p[21][26] ) );
  NOR2X0 U2285 ( .IN1(n269), .IN2(n316), .QN(\p[20][25] ) );
  NOR2X0 U2286 ( .IN1(n269), .IN2(n322), .QN(\p[18][23] ) );
  NOR2X0 U2287 ( .IN1(n268), .IN2(n325), .QN(\p[17][22] ) );
  DELLN1X2 U2288 ( .INP(n129), .Z(n342) );
  NOR2X0 U2289 ( .IN1(n277), .IN2(n310), .QN(\p[22][24] ) );
  NOR2X0 U2290 ( .IN1(n277), .IN2(n313), .QN(\p[21][23] ) );
  NOR2X0 U2291 ( .IN1(n277), .IN2(n316), .QN(\p[20][22] ) );
  NOR2X0 U2292 ( .IN1(n277), .IN2(n322), .QN(\p[18][20] ) );
  NOR2X0 U2293 ( .IN1(n277), .IN2(n325), .QN(\p[17][19] ) );
  NOR2X0 U2294 ( .IN1(n553), .IN2(n563), .QN(\p[1][3] ) );
  NOR2X0 U2295 ( .IN1(n173), .IN2(n369), .QN(\p[0][30] ) );
  NOR2X0 U2296 ( .IN1(n177), .IN2(n371), .QN(\p[0][29] ) );
  NOR2X0 U2297 ( .IN1(n181), .IN2(n371), .QN(\p[0][28] ) );
  NOR2X0 U2298 ( .IN1(n185), .IN2(n369), .QN(\p[0][27] ) );
  NOR2X0 U2299 ( .IN1(n189), .IN2(n369), .QN(\p[0][26] ) );
  NOR2X0 U2300 ( .IN1(n193), .IN2(n371), .QN(\p[0][25] ) );
  NOR2X0 U2301 ( .IN1(n197), .IN2(n369), .QN(\p[0][24] ) );
  NOR2X0 U2302 ( .IN1(n201), .IN2(n371), .QN(\p[0][23] ) );
  NOR2X0 U2303 ( .IN1(n205), .IN2(n369), .QN(\p[0][22] ) );
  NOR2X0 U2304 ( .IN1(n209), .IN2(n371), .QN(\p[0][21] ) );
  NOR2X0 U2305 ( .IN1(n213), .IN2(n369), .QN(\p[0][20] ) );
  NOR2X0 U2306 ( .IN1(n279), .IN2(n370), .QN(\p[0][2] ) );
  INVX0 U2307 ( .INP(A_reg[0]), .ZN(n555) );
  DELLN1X2 U2308 ( .INP(n549), .Z(n264) );
  NOR2X0 U2309 ( .IN1(n284), .IN2(n316), .QN(\p[20][20] ) );
  DELLN1X2 U2310 ( .INP(n85), .Z(n316) );
  INVX0 U2311 ( .INP(A_reg[1]), .ZN(n554) );
  NOR2X0 U2312 ( .IN1(n172), .IN2(n68), .QN(\p[1][31] ) );
  NOR2X0 U2313 ( .IN1(n176), .IN2(n366), .QN(\p[1][30] ) );
  NOR2X0 U2314 ( .IN1(n180), .IN2(n367), .QN(\p[1][29] ) );
  NOR2X0 U2315 ( .IN1(n184), .IN2(n368), .QN(\p[1][28] ) );
  NOR2X0 U2316 ( .IN1(n188), .IN2(n368), .QN(\p[1][27] ) );
  NOR2X0 U2317 ( .IN1(n192), .IN2(n368), .QN(\p[1][26] ) );
  NOR2X0 U2318 ( .IN1(n196), .IN2(n563), .QN(\p[1][25] ) );
  NOR2X0 U2319 ( .IN1(n200), .IN2(n67), .QN(\p[1][24] ) );
  NOR2X0 U2320 ( .IN1(n204), .IN2(n368), .QN(\p[1][23] ) );
  NOR2X0 U2321 ( .IN1(n208), .IN2(n67), .QN(\p[1][22] ) );
  NOR2X0 U2322 ( .IN1(n212), .IN2(n366), .QN(\p[1][21] ) );
  NOR2X0 U2323 ( .IN1(n554), .IN2(n68), .QN(\p[1][2] ) );
  INVX0 U2324 ( .INP(A_reg[7]), .ZN(n548) );
  NOR2X0 U2325 ( .IN1(n276), .IN2(n310), .QN(\p[22][25] ) );
  NOR2X0 U2326 ( .IN1(n275), .IN2(n313), .QN(\p[21][24] ) );
  NOR2X0 U2327 ( .IN1(n276), .IN2(n316), .QN(\p[20][23] ) );
  NOR2X0 U2328 ( .IN1(n274), .IN2(n322), .QN(\p[18][21] ) );
  NOR2X0 U2329 ( .IN1(n274), .IN2(n325), .QN(\p[17][20] ) );
  DELLN1X2 U2330 ( .INP(n564), .Z(n370) );
  NBUFFX2 U2331 ( .INP(n81), .Z(n321) );
  NOR2X0 U2332 ( .IN1(n247), .IN2(n319), .QN(\p[19][30] ) );
  NOR2X0 U2333 ( .IN1(n250), .IN2(n319), .QN(\p[19][29] ) );
  NOR2X0 U2334 ( .IN1(n255), .IN2(n319), .QN(\p[19][28] ) );
  NOR2X0 U2335 ( .IN1(n151), .IN2(n319), .QN(\p[19][26] ) );
  NOR2X0 U2336 ( .IN1(n270), .IN2(n319), .QN(\p[19][24] ) );
  NOR2X0 U2337 ( .IN1(n275), .IN2(n319), .QN(\p[19][22] ) );
  NOR2X0 U2338 ( .IN1(n277), .IN2(n319), .QN(\p[19][21] ) );
  NOR2X0 U2339 ( .IN1(n282), .IN2(n319), .QN(\p[19][20] ) );
  NBUFFX2 U2340 ( .INP(n81), .Z(n320) );
  NOR2X0 U2341 ( .IN1(n283), .IN2(n319), .QN(\p[19][19] ) );
  NOR2X0 U2342 ( .IN1(n285), .IN2(n325), .QN(\p[17][17] ) );
  DELLN1X2 U2343 ( .INP(n87), .Z(n325) );
  NOR2X0 U2344 ( .IN1(n285), .IN2(n322), .QN(\p[18][18] ) );
  DELLN1X2 U2345 ( .INP(n86), .Z(n322) );
  NOR2X0 U2346 ( .IN1(n277), .IN2(n286), .QN(\p[30][32] ) );
  NOR2X0 U2347 ( .IN1(n123), .IN2(n147), .QN(\p[9][11] ) );
  NOR2X0 U2348 ( .IN1(n147), .IN2(n125), .QN(\p[7][9] ) );
  NOR2X0 U2349 ( .IN1(n147), .IN2(n133), .QN(\p[6][8] ) );
  NOR2X0 U2350 ( .IN1(n258), .IN2(n310), .QN(\p[22][30] ) );
  NOR2X0 U2351 ( .IN1(n260), .IN2(n313), .QN(\p[21][29] ) );
  NOR2X0 U2352 ( .IN1(n258), .IN2(n316), .QN(\p[20][28] ) );
  NOR2X0 U2353 ( .IN1(n259), .IN2(n319), .QN(\p[19][27] ) );
  NOR2X0 U2354 ( .IN1(n260), .IN2(n322), .QN(\p[18][26] ) );
  NOR2X0 U2355 ( .IN1(n259), .IN2(n325), .QN(\p[17][25] ) );
  NOR2X0 U2356 ( .IN1(n113), .IN2(n141), .QN(\p[1][9] ) );
  DELLN1X2 U2357 ( .INP(n112), .Z(n259) );
  NBUFFX2 U2358 ( .INP(n82), .Z(n330) );
  NOR2X0 U2359 ( .IN1(n249), .IN2(n330), .QN(\p[16][27] ) );
  NOR2X0 U2360 ( .IN1(n250), .IN2(n329), .QN(\p[16][26] ) );
  NOR2X0 U2361 ( .IN1(n256), .IN2(n330), .QN(\p[16][25] ) );
  NOR2X0 U2362 ( .IN1(n260), .IN2(n329), .QN(\p[16][24] ) );
  NOR2X0 U2363 ( .IN1(n151), .IN2(n330), .QN(\p[16][23] ) );
  NOR2X0 U2364 ( .IN1(n268), .IN2(n328), .QN(\p[16][21] ) );
  NOR2X0 U2365 ( .IN1(n274), .IN2(n328), .QN(\p[16][19] ) );
  NOR2X0 U2366 ( .IN1(n277), .IN2(n328), .QN(\p[16][18] ) );
  NOR2X0 U2367 ( .IN1(n282), .IN2(n328), .QN(\p[16][17] ) );
  NBUFFX2 U2368 ( .INP(n82), .Z(n329) );
  NOR2X0 U2369 ( .IN1(n146), .IN2(n370), .QN(\p[0][3] ) );
  NOR2X0 U2370 ( .IN1(n551), .IN2(n142), .QN(\p[0][4] ) );
  NOR2X0 U2371 ( .IN1(n138), .IN2(n142), .QN(\p[0][5] ) );
  NOR2X0 U2372 ( .IN1(n148), .IN2(n142), .QN(\p[0][6] ) );
  NOR2X0 U2373 ( .IN1(n276), .IN2(n286), .QN(\p[30][33] ) );
  NOR2X0 U2374 ( .IN1(n557), .IN2(n146), .QN(\p[9][12] ) );
  NOR2X0 U2375 ( .IN1(n146), .IN2(n133), .QN(\p[6][9] ) );
  NOR2X0 U2376 ( .IN1(n146), .IN2(n145), .QN(\p[3][6] ) );
  NOR2X0 U2377 ( .IN1(n349), .IN2(n170), .QN(\p[9][39] ) );
  NOR2X0 U2378 ( .IN1(n348), .IN2(n174), .QN(\p[9][38] ) );
  NOR2X0 U2379 ( .IN1(n349), .IN2(n178), .QN(\p[9][37] ) );
  NOR2X0 U2380 ( .IN1(n347), .IN2(n182), .QN(\p[9][36] ) );
  NOR2X0 U2381 ( .IN1(n347), .IN2(n186), .QN(\p[9][35] ) );
  NOR2X0 U2382 ( .IN1(n348), .IN2(n190), .QN(\p[9][34] ) );
  NOR2X0 U2383 ( .IN1(n348), .IN2(n194), .QN(\p[9][33] ) );
  NOR2X0 U2384 ( .IN1(n120), .IN2(n123), .QN(\p[9][9] ) );
  DELLN1X2 U2385 ( .INP(n557), .Z(n348) );
  NOR2X0 U2386 ( .IN1(n138), .IN2(n145), .QN(\p[3][8] ) );
  DELLN1X2 U2387 ( .INP(n550), .Z(n268) );
  NOR2X0 U2388 ( .IN1(n246), .IN2(n341), .QN(\p[12][23] ) );
  NOR2X0 U2389 ( .IN1(n251), .IN2(n111), .QN(\p[12][22] ) );
  NOR2X0 U2390 ( .IN1(n256), .IN2(n111), .QN(\p[12][21] ) );
  NOR2X0 U2391 ( .IN1(n258), .IN2(n111), .QN(\p[12][20] ) );
  NOR2X0 U2392 ( .IN1(n150), .IN2(n111), .QN(\p[12][19] ) );
  NOR2X0 U2393 ( .IN1(n264), .IN2(n111), .QN(\p[12][18] ) );
  NOR2X0 U2394 ( .IN1(n269), .IN2(n111), .QN(\p[12][17] ) );
  NOR2X0 U2395 ( .IN1(n114), .IN2(n111), .QN(\p[12][16] ) );
  NOR2X0 U2396 ( .IN1(n552), .IN2(n111), .QN(\p[12][15] ) );
  NOR2X0 U2397 ( .IN1(n120), .IN2(n111), .QN(\p[12][12] ) );
  NOR2X0 U2398 ( .IN1(n278), .IN2(n111), .QN(\p[12][14] ) );
  NOR2X0 U2399 ( .IN1(n554), .IN2(n111), .QN(\p[12][13] ) );
  NOR2X0 U2400 ( .IN1(n113), .IN2(n142), .QN(\p[0][8] ) );
  NOR2X0 U2401 ( .IN1(n119), .IN2(n142), .QN(\p[0][9] ) );
  INVX0 U2402 ( .INP(A_reg[9]), .ZN(n547) );
  NOR2X0 U2403 ( .IN1(n170), .IN2(n361), .QN(\p[4][34] ) );
  NOR2X0 U2404 ( .IN1(n120), .IN2(n143), .QN(\p[4][4] ) );
  NOR2X0 U2405 ( .IN1(n555), .IN2(n328), .QN(\p[16][16] ) );
  NOR2X0 U2406 ( .IN1(n149), .IN2(n143), .QN(\p[4][8] ) );
  INVX0 U2407 ( .INP(A_reg[4]), .ZN(n551) );
  NOR2X0 U2408 ( .IN1(n114), .IN2(n310), .QN(\p[22][26] ) );
  NOR2X0 U2409 ( .IN1(n273), .IN2(n313), .QN(\p[21][25] ) );
  NOR2X0 U2410 ( .IN1(n114), .IN2(n316), .QN(\p[20][24] ) );
  NOR2X0 U2411 ( .IN1(n273), .IN2(n319), .QN(\p[19][23] ) );
  NOR2X0 U2412 ( .IN1(n273), .IN2(n322), .QN(\p[18][22] ) );
  NOR2X0 U2413 ( .IN1(n114), .IN2(n325), .QN(\p[17][21] ) );
  NOR2X0 U2414 ( .IN1(n273), .IN2(n328), .QN(\p[16][20] ) );
  NOR2X0 U2415 ( .IN1(n149), .IN2(n141), .QN(\p[1][5] ) );
  NOR2X0 U2416 ( .IN1(n226), .IN2(n357), .QN(\p[5][21] ) );
  NOR2X0 U2417 ( .IN1(n230), .IN2(n358), .QN(\p[5][20] ) );
  NOR2X0 U2418 ( .IN1(n234), .IN2(n117), .QN(\p[5][19] ) );
  NOR2X0 U2419 ( .IN1(n238), .IN2(n357), .QN(\p[5][18] ) );
  NOR2X0 U2420 ( .IN1(n245), .IN2(n561), .QN(\p[5][17] ) );
  NOR2X0 U2421 ( .IN1(n110), .IN2(n358), .QN(\p[5][16] ) );
  NOR2X0 U2422 ( .IN1(n121), .IN2(n115), .QN(\p[5][15] ) );
  NOR2X0 U2423 ( .IN1(n547), .IN2(n115), .QN(\p[5][14] ) );
  NOR2X0 U2424 ( .IN1(n112), .IN2(n561), .QN(\p[5][13] ) );
  NOR2X0 U2425 ( .IN1(n148), .IN2(n561), .QN(\p[5][11] ) );
  NOR2X0 U2426 ( .IN1(n138), .IN2(n115), .QN(\p[5][10] ) );
  NOR2X0 U2427 ( .IN1(n170), .IN2(n358), .QN(\p[5][35] ) );
  NOR2X0 U2428 ( .IN1(n174), .IN2(n117), .QN(\p[5][34] ) );
  NOR2X0 U2429 ( .IN1(n120), .IN2(n115), .QN(\p[5][5] ) );
  NOR2X0 U2430 ( .IN1(n551), .IN2(n115), .QN(\p[5][9] ) );
  NOR2X0 U2431 ( .IN1(n147), .IN2(n115), .QN(\p[5][7] ) );
  DELLN1X2 U2432 ( .INP(n558), .Z(n351) );
  INVX0 U2433 ( .INP(B_reg[8]), .ZN(n558) );
  NOR2X0 U2434 ( .IN1(n120), .IN2(n126), .QN(\p[8][8] ) );
  INVX0 U2435 ( .INP(A_reg[6]), .ZN(n549) );
  NOR2X0 U2436 ( .IN1(n554), .IN2(n135), .QN(\p[2][3] ) );
  NOR2X0 U2437 ( .IN1(n146), .IN2(n136), .QN(\p[2][5] ) );
  NOR2X0 U2438 ( .IN1(n152), .IN2(n136), .QN(\p[2][9] ) );
  NOR2X0 U2439 ( .IN1(n551), .IN2(n136), .QN(\p[2][6] ) );
  NOR2X0 U2440 ( .IN1(n138), .IN2(n136), .QN(\p[2][7] ) );
  DELLN1X2 U2441 ( .INP(n112), .Z(n260) );
  NOR2X0 U2442 ( .IN1(n222), .IN2(n359), .QN(\p[4][21] ) );
  NOR2X0 U2443 ( .IN1(n226), .IN2(n361), .QN(\p[4][20] ) );
  NOR2X0 U2444 ( .IN1(n230), .IN2(n359), .QN(\p[4][19] ) );
  NOR2X0 U2445 ( .IN1(n234), .IN2(n361), .QN(\p[4][18] ) );
  NOR2X0 U2446 ( .IN1(n238), .IN2(n360), .QN(\p[4][17] ) );
  NOR2X0 U2447 ( .IN1(n245), .IN2(n360), .QN(\p[4][16] ) );
  NOR2X0 U2448 ( .IN1(n110), .IN2(n360), .QN(\p[4][15] ) );
  NOR2X0 U2449 ( .IN1(n121), .IN2(n360), .QN(\p[4][14] ) );
  NOR2X0 U2450 ( .IN1(n547), .IN2(n360), .QN(\p[4][13] ) );
  NOR2X0 U2451 ( .IN1(n112), .IN2(n105), .QN(\p[4][12] ) );
  NOR2X0 U2452 ( .IN1(n152), .IN2(n105), .QN(\p[4][11] ) );
  NOR2X0 U2453 ( .IN1(n148), .IN2(n143), .QN(\p[4][10] ) );
  NOR2X0 U2454 ( .IN1(n147), .IN2(n143), .QN(\p[4][6] ) );
  DELLN1X2 U2455 ( .INP(n553), .Z(n277) );
  INVX0 U2456 ( .INP(A_reg[2]), .ZN(n553) );
  NOR2X0 U2457 ( .IN1(n282), .IN2(n286), .QN(\p[30][31] ) );
  NOR2X0 U2458 ( .IN1(n123), .IN2(n130), .QN(\p[9][10] ) );
  NOR2X0 U2459 ( .IN1(n130), .IN2(n126), .QN(\p[8][9] ) );
  NOR2X0 U2460 ( .IN1(n130), .IN2(n143), .QN(\p[4][5] ) );
  NOR2X0 U2461 ( .IN1(n106), .IN2(n125), .QN(\p[7][8] ) );
  NOR2X0 U2462 ( .IN1(n130), .IN2(n115), .QN(\p[5][6] ) );
  NOR2X0 U2463 ( .IN1(n130), .IN2(n133), .QN(\p[6][7] ) );
  INVX0 U2464 ( .INP(A_reg[3]), .ZN(n552) );
  NOR2X0 U2465 ( .IN1(n120), .IN2(n125), .QN(\p[7][7] ) );
  INVX0 U2466 ( .INP(B_reg[7]), .ZN(n559) );
  DELLN1X2 U2467 ( .INP(n550), .Z(n270) );
  INVX0 U2468 ( .INP(A_reg[5]), .ZN(n550) );
  NOR2X0 U2469 ( .IN1(n266), .IN2(n310), .QN(\p[22][28] ) );
  NOR2X0 U2470 ( .IN1(n264), .IN2(n313), .QN(\p[21][27] ) );
  NOR2X0 U2471 ( .IN1(n264), .IN2(n316), .QN(\p[20][26] ) );
  NOR2X0 U2472 ( .IN1(n265), .IN2(n319), .QN(\p[19][25] ) );
  NOR2X0 U2473 ( .IN1(n264), .IN2(n322), .QN(\p[18][24] ) );
  NOR2X0 U2474 ( .IN1(n264), .IN2(n325), .QN(\p[17][23] ) );
  NOR2X0 U2475 ( .IN1(n264), .IN2(n329), .QN(\p[16][22] ) );
  NOR2X0 U2476 ( .IN1(n246), .IN2(n332), .QN(\p[15][26] ) );
  NOR2X0 U2477 ( .IN1(n250), .IN2(n332), .QN(\p[15][25] ) );
  NOR2X0 U2478 ( .IN1(n256), .IN2(n332), .QN(\p[15][24] ) );
  NOR2X0 U2479 ( .IN1(n259), .IN2(n333), .QN(\p[15][23] ) );
  NOR2X0 U2480 ( .IN1(n261), .IN2(n331), .QN(\p[15][22] ) );
  NOR2X0 U2481 ( .IN1(n264), .IN2(n107), .QN(\p[15][21] ) );
  NOR2X0 U2482 ( .IN1(n269), .IN2(n107), .QN(\p[15][20] ) );
  NOR2X0 U2483 ( .IN1(n114), .IN2(n107), .QN(\p[15][19] ) );
  NOR2X0 U2484 ( .IN1(n274), .IN2(n107), .QN(\p[15][18] ) );
  NOR2X0 U2485 ( .IN1(n278), .IN2(n107), .QN(\p[15][17] ) );
  NOR2X0 U2486 ( .IN1(n281), .IN2(n107), .QN(\p[15][16] ) );
  NOR2X0 U2487 ( .IN1(n555), .IN2(n107), .QN(\p[15][15] ) );
  NOR2X0 U2488 ( .IN1(n120), .IN2(n133), .QN(\p[6][6] ) );
  INVX0 U2489 ( .INP(B_reg[6]), .ZN(n560) );
  NOR2X0 U2490 ( .IN1(n149), .IN2(n145), .QN(\p[3][7] ) );
  DELLN1X2 U2491 ( .INP(n149), .Z(n272) );
  NOR2X0 U2492 ( .IN1(n247), .IN2(n336), .QN(\p[14][25] ) );
  NOR2X0 U2493 ( .IN1(n250), .IN2(n336), .QN(\p[14][24] ) );
  NOR2X0 U2494 ( .IN1(n256), .IN2(n334), .QN(\p[14][23] ) );
  NOR2X0 U2495 ( .IN1(n260), .IN2(n334), .QN(\p[14][22] ) );
  NOR2X0 U2496 ( .IN1(n262), .IN2(n108), .QN(\p[14][21] ) );
  NOR2X0 U2497 ( .IN1(n264), .IN2(n108), .QN(\p[14][20] ) );
  NOR2X0 U2498 ( .IN1(n268), .IN2(n108), .QN(\p[14][19] ) );
  NOR2X0 U2499 ( .IN1(n273), .IN2(n108), .QN(\p[14][18] ) );
  NOR2X0 U2500 ( .IN1(n274), .IN2(n108), .QN(\p[14][17] ) );
  NOR2X0 U2501 ( .IN1(n553), .IN2(n108), .QN(\p[14][16] ) );
  NOR2X0 U2502 ( .IN1(n554), .IN2(n108), .QN(\p[14][15] ) );
  NOR2X0 U2503 ( .IN1(n555), .IN2(n108), .QN(\p[14][14] ) );
  INVX0 U2504 ( .INP(B_reg[9]), .ZN(n557) );
  NOR2X0 U2505 ( .IN1(n152), .IN2(n141), .QN(\p[1][8] ) );
  INVX0 U2506 ( .INP(B_reg[1]), .ZN(n563) );
  NOR2X0 U2507 ( .IN1(n152), .IN2(n142), .QN(\p[0][7] ) );
  INVX0 U2508 ( .INP(B_reg[0]), .ZN(n564) );
  NOR2X0 U2509 ( .IN1(n249), .IN2(n337), .QN(\p[13][24] ) );
  NOR2X0 U2510 ( .IN1(n252), .IN2(n337), .QN(\p[13][23] ) );
  NOR2X0 U2511 ( .IN1(n255), .IN2(n338), .QN(\p[13][22] ) );
  NOR2X0 U2512 ( .IN1(n259), .IN2(n338), .QN(\p[13][21] ) );
  NOR2X0 U2513 ( .IN1(n263), .IN2(n116), .QN(\p[13][20] ) );
  NOR2X0 U2514 ( .IN1(n264), .IN2(n116), .QN(\p[13][19] ) );
  NOR2X0 U2515 ( .IN1(n269), .IN2(n116), .QN(\p[13][18] ) );
  NOR2X0 U2516 ( .IN1(n273), .IN2(n116), .QN(\p[13][17] ) );
  NOR2X0 U2517 ( .IN1(n552), .IN2(n116), .QN(\p[13][16] ) );
  NOR2X0 U2518 ( .IN1(n553), .IN2(n116), .QN(\p[13][15] ) );
  NOR2X0 U2519 ( .IN1(n554), .IN2(n116), .QN(\p[13][14] ) );
  NOR2X0 U2520 ( .IN1(n120), .IN2(n116), .QN(\p[13][13] ) );
  DELLN1X2 U2521 ( .INP(n111), .Z(n339) );
  NOR2X0 U2522 ( .IN1(n238), .IN2(n350), .QN(\p[8][21] ) );
  NOR2X0 U2523 ( .IN1(n242), .IN2(n350), .QN(\p[8][20] ) );
  NOR2X0 U2524 ( .IN1(n246), .IN2(n350), .QN(\p[8][19] ) );
  NOR2X0 U2525 ( .IN1(n121), .IN2(n350), .QN(\p[8][18] ) );
  NOR2X0 U2526 ( .IN1(n257), .IN2(n351), .QN(\p[8][17] ) );
  NOR2X0 U2527 ( .IN1(n260), .IN2(n351), .QN(\p[8][16] ) );
  NOR2X0 U2528 ( .IN1(n548), .IN2(n558), .QN(\p[8][15] ) );
  NOR2X0 U2529 ( .IN1(n265), .IN2(n558), .QN(\p[8][14] ) );
  NOR2X0 U2530 ( .IN1(n268), .IN2(n558), .QN(\p[8][13] ) );
  NOR2X0 U2531 ( .IN1(n551), .IN2(n558), .QN(\p[8][12] ) );
  NOR2X0 U2532 ( .IN1(n552), .IN2(n558), .QN(\p[8][11] ) );
  NOR2X0 U2533 ( .IN1(n147), .IN2(n558), .QN(\p[8][10] ) );
  NOR2X0 U2534 ( .IN1(n247), .IN2(n128), .QN(\p[11][22] ) );
  NOR2X0 U2535 ( .IN1(n253), .IN2(n128), .QN(\p[11][21] ) );
  NOR2X0 U2536 ( .IN1(n254), .IN2(n127), .QN(\p[11][20] ) );
  NOR2X0 U2537 ( .IN1(n260), .IN2(n342), .QN(\p[11][19] ) );
  NOR2X0 U2538 ( .IN1(n262), .IN2(n342), .QN(\p[11][18] ) );
  NOR2X0 U2539 ( .IN1(n264), .IN2(n128), .QN(\p[11][17] ) );
  NOR2X0 U2540 ( .IN1(n269), .IN2(n342), .QN(\p[11][16] ) );
  NOR2X0 U2541 ( .IN1(n272), .IN2(n129), .QN(\p[11][15] ) );
  NOR2X0 U2542 ( .IN1(n552), .IN2(n129), .QN(\p[11][14] ) );
  NOR2X0 U2543 ( .IN1(n147), .IN2(n129), .QN(\p[11][13] ) );
  NOR2X0 U2544 ( .IN1(n554), .IN2(n129), .QN(\p[11][12] ) );
  NOR2X0 U2545 ( .IN1(n120), .IN2(n129), .QN(\p[11][11] ) );
  DELLN1X2 U2546 ( .INP(n561), .Z(n357) );
  NOR2X0 U2547 ( .IN1(n146), .IN2(n115), .QN(\p[5][8] ) );
  INVX0 U2548 ( .INP(B_reg[5]), .ZN(n561) );
  NOR2X0 U2549 ( .IN1(n234), .IN2(n353), .QN(\p[7][21] ) );
  NOR2X0 U2550 ( .IN1(n238), .IN2(n124), .QN(\p[7][20] ) );
  NOR2X0 U2551 ( .IN1(n243), .IN2(n124), .QN(\p[7][19] ) );
  NOR2X0 U2552 ( .IN1(n247), .IN2(n354), .QN(\p[7][18] ) );
  NOR2X0 U2553 ( .IN1(n121), .IN2(n352), .QN(\p[7][17] ) );
  NOR2X0 U2554 ( .IN1(n119), .IN2(n559), .QN(\p[7][16] ) );
  NOR2X0 U2555 ( .IN1(n113), .IN2(n559), .QN(\p[7][15] ) );
  NOR2X0 U2556 ( .IN1(n548), .IN2(n559), .QN(\p[7][14] ) );
  NOR2X0 U2557 ( .IN1(n267), .IN2(n559), .QN(\p[7][13] ) );
  NOR2X0 U2558 ( .IN1(n137), .IN2(n125), .QN(\p[7][12] ) );
  NOR2X0 U2559 ( .IN1(n149), .IN2(n125), .QN(\p[7][11] ) );
  NOR2X0 U2560 ( .IN1(n552), .IN2(n125), .QN(\p[7][10] ) );
  NOR2X0 U2561 ( .IN1(n148), .IN2(n136), .QN(\p[2][8] ) );
  INVX0 U2562 ( .INP(B_reg[2]), .ZN(n562) );
  NOR2X0 U2563 ( .IN1(n215), .IN2(n365), .QN(\p[2][21] ) );
  NOR2X0 U2564 ( .IN1(n219), .IN2(n364), .QN(\p[2][20] ) );
  NOR2X0 U2565 ( .IN1(n223), .IN2(n134), .QN(\p[2][19] ) );
  NOR2X0 U2566 ( .IN1(n227), .IN2(n135), .QN(\p[2][18] ) );
  NOR2X0 U2567 ( .IN1(n231), .IN2(n135), .QN(\p[2][17] ) );
  NOR2X0 U2568 ( .IN1(n235), .IN2(n135), .QN(\p[2][16] ) );
  NOR2X0 U2569 ( .IN1(n239), .IN2(n562), .QN(\p[2][15] ) );
  NOR2X0 U2570 ( .IN1(n118), .IN2(n562), .QN(\p[2][14] ) );
  NOR2X0 U2571 ( .IN1(n113), .IN2(n136), .QN(\p[2][10] ) );
  NOR2X0 U2572 ( .IN1(n110), .IN2(n562), .QN(\p[2][13] ) );
  NOR2X0 U2573 ( .IN1(n121), .IN2(n562), .QN(\p[2][12] ) );
  NOR2X0 U2574 ( .IN1(n119), .IN2(n136), .QN(\p[2][11] ) );
  NOR2X0 U2575 ( .IN1(n230), .IN2(n356), .QN(\p[6][21] ) );
  NOR2X0 U2576 ( .IN1(n234), .IN2(n356), .QN(\p[6][20] ) );
  NOR2X0 U2577 ( .IN1(n238), .IN2(n356), .QN(\p[6][19] ) );
  NOR2X0 U2578 ( .IN1(n243), .IN2(n132), .QN(\p[6][18] ) );
  NOR2X0 U2579 ( .IN1(n248), .IN2(n131), .QN(\p[6][17] ) );
  NOR2X0 U2580 ( .IN1(n121), .IN2(n560), .QN(\p[6][16] ) );
  NOR2X0 U2581 ( .IN1(n547), .IN2(n560), .QN(\p[6][15] ) );
  NOR2X0 U2582 ( .IN1(n112), .IN2(n560), .QN(\p[6][14] ) );
  NOR2X0 U2583 ( .IN1(n548), .IN2(n560), .QN(\p[6][13] ) );
  NOR2X0 U2584 ( .IN1(n148), .IN2(n133), .QN(\p[6][12] ) );
  NOR2X0 U2585 ( .IN1(n138), .IN2(n560), .QN(\p[6][11] ) );
  NOR2X0 U2586 ( .IN1(n149), .IN2(n133), .QN(\p[6][10] ) );
  NOR2X0 U2587 ( .IN1(n218), .IN2(n363), .QN(\p[3][21] ) );
  NOR2X0 U2588 ( .IN1(n222), .IN2(n363), .QN(\p[3][20] ) );
  NOR2X0 U2589 ( .IN1(n226), .IN2(n363), .QN(\p[3][19] ) );
  NOR2X0 U2590 ( .IN1(n230), .IN2(n363), .QN(\p[3][18] ) );
  NOR2X0 U2591 ( .IN1(n234), .IN2(n363), .QN(\p[3][17] ) );
  NOR2X0 U2592 ( .IN1(n238), .IN2(n362), .QN(\p[3][16] ) );
  NOR2X0 U2593 ( .IN1(n118), .IN2(n363), .QN(\p[3][15] ) );
  NOR2X0 U2594 ( .IN1(n110), .IN2(n144), .QN(\p[3][14] ) );
  NOR2X0 U2595 ( .IN1(n121), .IN2(n145), .QN(\p[3][13] ) );
  NOR2X0 U2596 ( .IN1(n113), .IN2(n145), .QN(\p[3][11] ) );
  NOR2X0 U2597 ( .IN1(n119), .IN2(n109), .QN(\p[3][12] ) );
  NOR2X0 U2598 ( .IN1(n152), .IN2(n109), .QN(\p[3][10] ) );
  NOR2X0 U2599 ( .IN1(n249), .IN2(n72), .QN(\p[10][21] ) );
  NOR2X0 U2600 ( .IN1(n121), .IN2(n70), .QN(\p[10][20] ) );
  NOR2X0 U2601 ( .IN1(n257), .IN2(n71), .QN(\p[10][19] ) );
  NOR2X0 U2602 ( .IN1(n259), .IN2(n72), .QN(\p[10][18] ) );
  NOR2X0 U2603 ( .IN1(n261), .IN2(n71), .QN(\p[10][17] ) );
  NOR2X0 U2604 ( .IN1(n266), .IN2(n72), .QN(\p[10][16] ) );
  NOR2X0 U2605 ( .IN1(n270), .IN2(n139), .QN(\p[10][15] ) );
  NOR2X0 U2606 ( .IN1(n272), .IN2(n139), .QN(\p[10][14] ) );
  NOR2X0 U2607 ( .IN1(n552), .IN2(n139), .QN(\p[10][13] ) );
  NOR2X0 U2608 ( .IN1(n130), .IN2(n139), .QN(\p[10][11] ) );
  NOR2X0 U2609 ( .IN1(n553), .IN2(n139), .QN(\p[10][12] ) );
  NOR2X0 U2610 ( .IN1(n555), .IN2(n139), .QN(\p[10][10] ) );
  NOR2X0 U2611 ( .IN1(n284), .IN2(n368), .QN(\p[1][1] ) );
  NOR2X0 U2612 ( .IN1(n216), .IN2(n67), .QN(\p[1][20] ) );
  NOR2X0 U2613 ( .IN1(n220), .IN2(n563), .QN(\p[1][19] ) );
  NOR2X0 U2614 ( .IN1(n224), .IN2(n367), .QN(\p[1][18] ) );
  NOR2X0 U2615 ( .IN1(n228), .IN2(n366), .QN(\p[1][17] ) );
  NOR2X0 U2616 ( .IN1(n232), .IN2(n68), .QN(\p[1][16] ) );
  NOR2X0 U2617 ( .IN1(n236), .IN2(n67), .QN(\p[1][15] ) );
  NOR2X0 U2618 ( .IN1(n240), .IN2(n68), .QN(\p[1][14] ) );
  NOR2X0 U2619 ( .IN1(n118), .IN2(n68), .QN(\p[1][13] ) );
  NOR2X0 U2620 ( .IN1(n110), .IN2(n140), .QN(\p[1][12] ) );
  NOR2X0 U2621 ( .IN1(n119), .IN2(n140), .QN(\p[1][10] ) );
  NOR2X0 U2622 ( .IN1(n284), .IN2(n371), .QN(\p[0][0] ) );
  NOR2X0 U2623 ( .IN1(n281), .IN2(n369), .QN(\p[0][1] ) );
  NOR2X0 U2624 ( .IN1(n217), .IN2(n371), .QN(\p[0][19] ) );
  NOR2X0 U2625 ( .IN1(n221), .IN2(n371), .QN(\p[0][18] ) );
  NOR2X0 U2626 ( .IN1(n225), .IN2(n369), .QN(\p[0][17] ) );
  NOR2X0 U2627 ( .IN1(n229), .IN2(n370), .QN(\p[0][16] ) );
  NOR2X0 U2628 ( .IN1(n233), .IN2(n370), .QN(\p[0][15] ) );
  NOR2X0 U2629 ( .IN1(n237), .IN2(n370), .QN(\p[0][14] ) );
  NOR2X0 U2630 ( .IN1(n241), .IN2(n370), .QN(\p[0][13] ) );
  NOR2X0 U2631 ( .IN1(n118), .IN2(n564), .QN(\p[0][12] ) );
  NOR2X0 U2632 ( .IN1(n110), .IN2(n564), .QN(\p[0][11] ) );
  NOR2X0 U2633 ( .IN1(n121), .IN2(n142), .QN(\p[0][10] ) );
  DELLN1X2 U2634 ( .INP(\p[63][63] ), .Z(n502) );
  NBUFFX4 U2635 ( .INP(\p[2][63] ), .Z(n514) );
  NBUFFX4 U2636 ( .INP(\p[4][63] ), .Z(n523) );
  NBUFFX4 U2637 ( .INP(\p[4][63] ), .Z(n524) );
  DELLN1X2 U2638 ( .INP(A_reg[31]), .Z(n544) );
endmodule

