
module SeqMult_DW01_inc_0 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;

  wire   [31:2] carry;

  HA_X1 U1_1_30 ( .A(A[30]), .B(carry[30]), .CO(carry[31]), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[31]), .B(A[31]), .Z(SUM[31]) );
endmodule


module SeqMult_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [0:0] B;
  output [32:0] PRODUCT;
  input TC;
  wire   n1, n2, n3;

  BUF_X1 U2 ( .A(B[0]), .Z(n3) );
  CLKBUF_X3 U3 ( .A(n1), .Z(n2) );
  BUF_X2 U4 ( .A(B[0]), .Z(n1) );
  AND2_X1 U5 ( .A1(A[0]), .A2(n3), .ZN(PRODUCT[0]) );
  AND2_X1 U6 ( .A1(A[1]), .A2(n3), .ZN(PRODUCT[1]) );
  AND2_X1 U7 ( .A1(A[2]), .A2(n3), .ZN(PRODUCT[2]) );
  AND2_X1 U8 ( .A1(A[3]), .A2(n1), .ZN(PRODUCT[3]) );
  AND2_X1 U9 ( .A1(A[4]), .A2(n3), .ZN(PRODUCT[4]) );
  AND2_X1 U10 ( .A1(B[0]), .A2(A[5]), .ZN(PRODUCT[5]) );
  AND2_X1 U11 ( .A1(A[6]), .A2(n3), .ZN(PRODUCT[6]) );
  AND2_X1 U12 ( .A1(A[7]), .A2(n1), .ZN(PRODUCT[7]) );
  AND2_X1 U13 ( .A1(A[8]), .A2(n1), .ZN(PRODUCT[8]) );
  AND2_X1 U14 ( .A1(A[9]), .A2(n3), .ZN(PRODUCT[9]) );
  AND2_X1 U15 ( .A1(A[10]), .A2(n1), .ZN(PRODUCT[10]) );
  AND2_X1 U16 ( .A1(A[11]), .A2(n1), .ZN(PRODUCT[11]) );
  AND2_X1 U17 ( .A1(A[12]), .A2(n2), .ZN(PRODUCT[12]) );
  AND2_X1 U18 ( .A1(A[13]), .A2(n1), .ZN(PRODUCT[13]) );
  AND2_X1 U19 ( .A1(A[14]), .A2(n2), .ZN(PRODUCT[14]) );
  AND2_X1 U20 ( .A1(A[15]), .A2(n2), .ZN(PRODUCT[15]) );
  AND2_X1 U21 ( .A1(A[16]), .A2(n2), .ZN(PRODUCT[16]) );
  AND2_X1 U22 ( .A1(A[17]), .A2(n2), .ZN(PRODUCT[17]) );
  AND2_X1 U23 ( .A1(A[18]), .A2(n1), .ZN(PRODUCT[18]) );
  AND2_X1 U24 ( .A1(A[19]), .A2(n2), .ZN(PRODUCT[19]) );
  AND2_X1 U25 ( .A1(A[20]), .A2(n2), .ZN(PRODUCT[20]) );
  AND2_X1 U26 ( .A1(A[21]), .A2(n2), .ZN(PRODUCT[21]) );
  AND2_X1 U27 ( .A1(A[22]), .A2(n2), .ZN(PRODUCT[22]) );
  AND2_X1 U28 ( .A1(A[23]), .A2(n2), .ZN(PRODUCT[23]) );
  AND2_X1 U29 ( .A1(A[24]), .A2(n2), .ZN(PRODUCT[24]) );
  AND2_X1 U30 ( .A1(A[25]), .A2(n2), .ZN(PRODUCT[25]) );
  AND2_X1 U31 ( .A1(A[26]), .A2(n2), .ZN(PRODUCT[26]) );
  AND2_X1 U32 ( .A1(A[27]), .A2(n2), .ZN(PRODUCT[27]) );
  AND2_X1 U33 ( .A1(A[28]), .A2(n2), .ZN(PRODUCT[28]) );
  AND2_X1 U34 ( .A1(A[29]), .A2(n2), .ZN(PRODUCT[29]) );
  AND2_X1 U35 ( .A1(A[30]), .A2(n2), .ZN(PRODUCT[30]) );
  AND2_X1 U36 ( .A1(A[31]), .A2(n2), .ZN(PRODUCT[31]) );
endmodule


module SeqMult_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND3_X1 U3 ( .A1(n98), .A2(n99), .A3(n2), .ZN(n1) );
  AND3_X1 U4 ( .A1(n100), .A2(n128), .A3(n101), .ZN(n2) );
  NOR2_X1 U5 ( .A1(B[61]), .A2(n9), .ZN(n3) );
  OR2_X2 U6 ( .A1(B[60]), .A2(n8), .ZN(n9) );
  AND4_X1 U7 ( .A1(n61), .A2(n62), .A3(n63), .A4(n64), .ZN(n6) );
  OR2_X1 U8 ( .A1(B[58]), .A2(n11), .ZN(n10) );
  AND2_X1 U9 ( .A1(n140), .A2(n141), .ZN(n4) );
  XOR2_X1 U10 ( .A(n68), .B(B[47]), .Z(DIFF[47]) );
  NOR2_X1 U11 ( .A1(B[33]), .A2(n96), .ZN(n95) );
  NOR2_X1 U12 ( .A1(n79), .A2(n66), .ZN(n78) );
  OR2_X1 U13 ( .A1(n70), .A2(n65), .ZN(n5) );
  AND2_X1 U14 ( .A1(n71), .A2(n77), .ZN(n76) );
  NOR2_X1 U15 ( .A1(B[36]), .A2(n79), .ZN(n88) );
  NAND4_X1 U16 ( .A1(n90), .A2(n91), .A3(n92), .A4(n93), .ZN(n67) );
  NOR2_X1 U17 ( .A1(B[61]), .A2(n9), .ZN(n38) );
  NOR2_X1 U18 ( .A1(B[40]), .A2(n70), .ZN(n77) );
  NOR2_X1 U19 ( .A1(B[45]), .A2(n7), .ZN(n69) );
  OR2_X1 U20 ( .A1(B[44]), .A2(n5), .ZN(n7) );
  NOR2_X1 U21 ( .A1(n42), .A2(n67), .ZN(n89) );
  OR2_X1 U22 ( .A1(B[59]), .A2(n10), .ZN(n8) );
  OR2_X1 U23 ( .A1(B[57]), .A2(n24), .ZN(n11) );
  AND2_X1 U24 ( .A1(n6), .A2(n59), .ZN(n12) );
  AND2_X1 U25 ( .A1(n51), .A2(n22), .ZN(n13) );
  AND2_X1 U26 ( .A1(n15), .A2(n46), .ZN(n14) );
  AND2_X1 U27 ( .A1(n13), .A2(n48), .ZN(n15) );
  AND2_X1 U28 ( .A1(n12), .A2(n56), .ZN(n16) );
  NAND2_X1 U29 ( .A1(n45), .A2(n90), .ZN(n96) );
  AND2_X1 U30 ( .A1(n14), .A2(n43), .ZN(n17) );
  AND2_X1 U31 ( .A1(n88), .A2(n80), .ZN(n18) );
  NAND2_X1 U32 ( .A1(n76), .A2(n73), .ZN(n75) );
  NAND2_X1 U33 ( .A1(n95), .A2(n92), .ZN(n94) );
  NAND2_X1 U34 ( .A1(n14), .A2(n45), .ZN(n44) );
  NAND2_X1 U35 ( .A1(n15), .A2(n45), .ZN(n47) );
  NAND2_X1 U36 ( .A1(n13), .A2(n45), .ZN(n49) );
  NAND2_X1 U37 ( .A1(n23), .A2(n45), .ZN(n50) );
  NAND2_X1 U38 ( .A1(n51), .A2(n45), .ZN(n52) );
  NAND2_X1 U39 ( .A1(n16), .A2(n45), .ZN(n55) );
  NAND2_X1 U40 ( .A1(n12), .A2(n45), .ZN(n58) );
  NAND2_X1 U41 ( .A1(n6), .A2(n45), .ZN(n60) );
  NAND2_X1 U42 ( .A1(n45), .A2(n25), .ZN(n24) );
  NAND2_X1 U43 ( .A1(n18), .A2(n82), .ZN(n87) );
  NAND2_X1 U44 ( .A1(n17), .A2(n45), .ZN(n41) );
  NAND2_X1 U45 ( .A1(n69), .A2(n63), .ZN(n68) );
  INV_X1 U46 ( .A(n42), .ZN(n45) );
  NOR2_X1 U47 ( .A1(n112), .A2(n102), .ZN(n111) );
  NOR2_X1 U48 ( .A1(n103), .A2(n104), .ZN(n120) );
  NOR2_X1 U49 ( .A1(B[13]), .A2(n19), .ZN(n153) );
  NOR2_X1 U50 ( .A1(B[17]), .A2(n139), .ZN(n137) );
  NOR2_X1 U51 ( .A1(n151), .A2(n150), .ZN(n28) );
  NOR2_X1 U52 ( .A1(n157), .A2(n149), .ZN(n155) );
  OR2_X1 U53 ( .A1(B[12]), .A2(n154), .ZN(n19) );
  NOR2_X1 U54 ( .A1(n150), .A2(n151), .ZN(n147) );
  INV_X1 U55 ( .A(B[34]), .ZN(n92) );
  INV_X1 U56 ( .A(B[32]), .ZN(n90) );
  INV_X1 U57 ( .A(B[46]), .ZN(n63) );
  INV_X1 U58 ( .A(B[42]), .ZN(n73) );
  INV_X1 U59 ( .A(B[38]), .ZN(n82) );
  INV_X1 U60 ( .A(B[40]), .ZN(n72) );
  INV_X1 U61 ( .A(B[41]), .ZN(n71) );
  INV_X1 U62 ( .A(B[37]), .ZN(n80) );
  INV_X1 U63 ( .A(B[35]), .ZN(n93) );
  INV_X1 U64 ( .A(n151), .ZN(n57) );
  INV_X1 U65 ( .A(B[36]), .ZN(n81) );
  INV_X1 U66 ( .A(n103), .ZN(n128) );
  INV_X1 U67 ( .A(B[55]), .ZN(n43) );
  INV_X1 U68 ( .A(B[54]), .ZN(n46) );
  INV_X1 U69 ( .A(B[53]), .ZN(n48) );
  INV_X1 U70 ( .A(B[50]), .ZN(n54) );
  INV_X1 U71 ( .A(B[49]), .ZN(n56) );
  INV_X1 U72 ( .A(B[48]), .ZN(n59) );
  INV_X1 U73 ( .A(B[43]), .ZN(n74) );
  INV_X1 U74 ( .A(B[47]), .ZN(n64) );
  INV_X1 U75 ( .A(B[39]), .ZN(n83) );
  INV_X1 U76 ( .A(B[56]), .ZN(n40) );
  INV_X1 U77 ( .A(B[33]), .ZN(n91) );
  NAND4_X1 U78 ( .A1(n36), .A2(n39), .A3(n33), .A4(n31), .ZN(n150) );
  NAND4_X1 U79 ( .A1(n110), .A2(n135), .A3(n86), .A4(n84), .ZN(n151) );
  AND2_X1 U80 ( .A1(n113), .A2(n119), .ZN(n118) );
  AND2_X1 U81 ( .A1(n121), .A2(n127), .ZN(n126) );
  NAND4_X1 U82 ( .A1(n113), .A2(n114), .A3(n115), .A4(n116), .ZN(n102) );
  NAND4_X1 U83 ( .A1(n121), .A2(n122), .A3(n123), .A4(n124), .ZN(n104) );
  NAND4_X1 U84 ( .A1(n27), .A2(n29), .A3(n158), .A4(n159), .ZN(n149) );
  NAND4_X1 U85 ( .A1(n129), .A2(n130), .A3(n131), .A4(n132), .ZN(n103) );
  NOR2_X1 U86 ( .A1(B[16]), .A2(n133), .ZN(n129) );
  NOR2_X1 U87 ( .A1(B[20]), .A2(n103), .ZN(n127) );
  AND2_X1 U88 ( .A1(n98), .A2(n111), .ZN(n109) );
  NOR2_X1 U89 ( .A1(B[24]), .A2(n112), .ZN(n119) );
  AND2_X1 U90 ( .A1(n99), .A2(n109), .ZN(n106) );
  AND2_X1 U91 ( .A1(n36), .A2(n35), .ZN(n32) );
  NOR2_X1 U92 ( .A1(n157), .A2(B[8]), .ZN(n26) );
  NOR2_X1 U93 ( .A1(n151), .A2(B[4]), .ZN(n35) );
  NAND2_X1 U94 ( .A1(n97), .A2(n1), .ZN(n42) );
  NOR2_X1 U95 ( .A1(B[31]), .A2(B[30]), .ZN(n97) );
  NOR2_X1 U96 ( .A1(n142), .A2(B[14]), .ZN(n140) );
  NAND2_X1 U97 ( .A1(n4), .A2(n134), .ZN(n139) );
  INV_X1 U98 ( .A(B[62]), .ZN(n37) );
  NAND2_X1 U99 ( .A1(n118), .A2(n115), .ZN(n117) );
  NAND2_X1 U100 ( .A1(n126), .A2(n123), .ZN(n125) );
  NAND2_X1 U101 ( .A1(n153), .A2(n143), .ZN(n152) );
  NAND2_X1 U102 ( .A1(n137), .A2(n131), .ZN(n136) );
  NAND2_X1 U103 ( .A1(n106), .A2(n107), .ZN(n105) );
  NAND2_X1 U104 ( .A1(n32), .A2(n33), .ZN(n30) );
  AND2_X1 U105 ( .A1(n26), .A2(n27), .ZN(n160) );
  NAND2_X1 U106 ( .A1(n144), .A2(n145), .ZN(n142) );
  NOR2_X1 U107 ( .A1(n146), .A2(B[12]), .ZN(n144) );
  NAND2_X1 U108 ( .A1(n147), .A2(n148), .ZN(n146) );
  AND2_X1 U109 ( .A1(n160), .A2(n158), .ZN(n20) );
  AND2_X1 U110 ( .A1(n85), .A2(n86), .ZN(n21) );
  INV_X1 U111 ( .A(B[2]), .ZN(n86) );
  INV_X1 U112 ( .A(\B[0] ), .ZN(n135) );
  INV_X1 U113 ( .A(B[6]), .ZN(n33) );
  INV_X1 U114 ( .A(B[10]), .ZN(n158) );
  INV_X1 U115 ( .A(B[14]), .ZN(n143) );
  INV_X1 U116 ( .A(B[8]), .ZN(n29) );
  INV_X1 U117 ( .A(B[4]), .ZN(n39) );
  INV_X1 U118 ( .A(B[20]), .ZN(n122) );
  INV_X1 U119 ( .A(B[29]), .ZN(n99) );
  INV_X1 U120 ( .A(B[26]), .ZN(n115) );
  INV_X1 U121 ( .A(B[22]), .ZN(n123) );
  INV_X1 U122 ( .A(B[16]), .ZN(n134) );
  INV_X1 U123 ( .A(B[9]), .ZN(n27) );
  INV_X1 U124 ( .A(B[18]), .ZN(n131) );
  INV_X1 U125 ( .A(B[15]), .ZN(n141) );
  INV_X1 U126 ( .A(B[12]), .ZN(n156) );
  INV_X1 U127 ( .A(B[24]), .ZN(n114) );
  INV_X1 U128 ( .A(B[3]), .ZN(n84) );
  INV_X1 U129 ( .A(B[28]), .ZN(n98) );
  INV_X1 U130 ( .A(B[25]), .ZN(n113) );
  INV_X1 U131 ( .A(B[5]), .ZN(n36) );
  INV_X1 U132 ( .A(B[1]), .ZN(n110) );
  INV_X1 U133 ( .A(B[21]), .ZN(n121) );
  INV_X1 U134 ( .A(B[11]), .ZN(n159) );
  INV_X1 U135 ( .A(B[19]), .ZN(n132) );
  INV_X1 U136 ( .A(B[17]), .ZN(n130) );
  INV_X1 U137 ( .A(B[27]), .ZN(n116) );
  INV_X1 U138 ( .A(B[23]), .ZN(n124) );
  INV_X1 U139 ( .A(B[7]), .ZN(n31) );
  INV_X1 U140 ( .A(B[13]), .ZN(n145) );
  INV_X1 U141 ( .A(B[30]), .ZN(n107) );
  NOR2_X1 U142 ( .A1(B[1]), .A2(\B[0] ), .ZN(n85) );
  XOR2_X1 U143 ( .A(n28), .B(n29), .Z(DIFF[8]) );
  XOR2_X1 U144 ( .A(n35), .B(n36), .Z(DIFF[5]) );
  XOR2_X1 U145 ( .A(n63), .B(n69), .Z(DIFF[46]) );
  XOR2_X1 U146 ( .A(n75), .B(B[43]), .Z(DIFF[43]) );
  XOR2_X1 U147 ( .A(n7), .B(B[45]), .Z(DIFF[45]) );
  XOR2_X1 U148 ( .A(n73), .B(n76), .Z(DIFF[42]) );
  XOR2_X1 U149 ( .A(n87), .B(B[39]), .Z(DIFF[39]) );
  XOR2_X1 U150 ( .A(n5), .B(B[44]), .Z(DIFF[44]) );
  XOR2_X1 U151 ( .A(n11), .B(B[58]), .Z(DIFF[58]) );
  XOR2_X1 U152 ( .A(n9), .B(B[61]), .Z(DIFF[61]) );
  XOR2_X1 U153 ( .A(n8), .B(B[60]), .Z(DIFF[60]) );
  XOR2_X1 U154 ( .A(n10), .B(B[59]), .Z(DIFF[59]) );
  XOR2_X1 U155 ( .A(n109), .B(n99), .Z(DIFF[29]) );
  XOR2_X1 U156 ( .A(n111), .B(n98), .Z(DIFF[28]) );
  XOR2_X1 U157 ( .A(n117), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U158 ( .A(n115), .B(n118), .Z(DIFF[26]) );
  XOR2_X1 U159 ( .A(n119), .B(n113), .Z(DIFF[25]) );
  XOR2_X1 U160 ( .A(n120), .B(n114), .Z(DIFF[24]) );
  XOR2_X1 U161 ( .A(n125), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U162 ( .A(n123), .B(n126), .Z(DIFF[22]) );
  XOR2_X1 U163 ( .A(n127), .B(n121), .Z(DIFF[21]) );
  XOR2_X1 U164 ( .A(n128), .B(n122), .Z(DIFF[20]) );
  XOR2_X1 U165 ( .A(n136), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U166 ( .A(n138), .B(B[18]), .Z(DIFF[18]) );
  XOR2_X1 U167 ( .A(n139), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U168 ( .A(n4), .B(n134), .Z(DIFF[16]) );
  XOR2_X1 U169 ( .A(n152), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U170 ( .A(n153), .B(n143), .Z(DIFF[14]) );
  XOR2_X1 U171 ( .A(n19), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U172 ( .A(n155), .B(n156), .Z(DIFF[12]) );
  XOR2_X1 U173 ( .A(n20), .B(n159), .Z(DIFF[11]) );
  XOR2_X1 U174 ( .A(n160), .B(n158), .Z(DIFF[10]) );
  XOR2_X1 U175 ( .A(n26), .B(n27), .Z(DIFF[9]) );
  XOR2_X1 U176 ( .A(n30), .B(B[7]), .Z(DIFF[7]) );
  XOR2_X1 U177 ( .A(n34), .B(B[6]), .Z(DIFF[6]) );
  XOR2_X1 U178 ( .A(n108), .B(B[30]), .Z(DIFF[30]) );
  XOR2_X1 U179 ( .A(n44), .B(B[55]), .Z(DIFF[55]) );
  XOR2_X1 U180 ( .A(n47), .B(B[54]), .Z(DIFF[54]) );
  XOR2_X1 U181 ( .A(n49), .B(B[53]), .Z(DIFF[53]) );
  XOR2_X1 U182 ( .A(n50), .B(B[52]), .Z(DIFF[52]) );
  XOR2_X1 U183 ( .A(n52), .B(B[51]), .Z(DIFF[51]) );
  XOR2_X1 U184 ( .A(n55), .B(B[50]), .Z(DIFF[50]) );
  XOR2_X1 U185 ( .A(n58), .B(B[49]), .Z(DIFF[49]) );
  XOR2_X1 U186 ( .A(n60), .B(B[48]), .Z(DIFF[48]) );
  XOR2_X1 U187 ( .A(n78), .B(n72), .Z(DIFF[40]) );
  XOR2_X1 U188 ( .A(n80), .B(n88), .Z(DIFF[37]) );
  XOR2_X1 U189 ( .A(n89), .B(n81), .Z(DIFF[36]) );
  XOR2_X1 U190 ( .A(n94), .B(B[35]), .Z(DIFF[35]) );
  XOR2_X1 U191 ( .A(n92), .B(n95), .Z(DIFF[34]) );
  XOR2_X1 U192 ( .A(n96), .B(B[33]), .Z(DIFF[33]) );
  XOR2_X1 U193 ( .A(n45), .B(n90), .Z(DIFF[32]) );
  XOR2_X1 U194 ( .A(n105), .B(B[31]), .Z(DIFF[31]) );
  XOR2_X1 U195 ( .A(n41), .B(B[56]), .Z(DIFF[56]) );
  XOR2_X1 U196 ( .A(n77), .B(n71), .Z(DIFF[41]) );
  XOR2_X1 U197 ( .A(n24), .B(B[57]), .Z(DIFF[57]) );
  XOR2_X1 U198 ( .A(n82), .B(n18), .Z(DIFF[38]) );
  NAND2_X1 U199 ( .A1(n37), .A2(n3), .ZN(DIFF[63]) );
  XOR2_X1 U200 ( .A(n57), .B(n39), .Z(DIFF[4]) );
  XOR2_X1 U201 ( .A(n21), .B(n84), .Z(DIFF[3]) );
  XOR2_X1 U202 ( .A(n85), .B(n86), .Z(DIFF[2]) );
  XOR2_X1 U203 ( .A(n135), .B(n110), .Z(DIFF[1]) );
  NOR2_X1 U204 ( .A1(B[51]), .A2(B[52]), .ZN(n22) );
  NOR2_X1 U205 ( .A1(n53), .A2(B[51]), .ZN(n23) );
  NAND4_X1 U206 ( .A1(n80), .A2(n81), .A3(n82), .A4(n83), .ZN(n66) );
  AND2_X1 U207 ( .A1(n17), .A2(n40), .ZN(n25) );
  NAND4_X1 U208 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(n65) );
  XNOR2_X1 U209 ( .A(B[62]), .B(n38), .ZN(DIFF[62]) );
  NAND2_X1 U210 ( .A1(n16), .A2(n54), .ZN(n53) );
  NOR3_X1 U211 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n61) );
  INV_X1 U212 ( .A(n32), .ZN(n34) );
  INV_X1 U213 ( .A(n53), .ZN(n51) );
  NOR2_X1 U214 ( .A1(B[45]), .A2(B[44]), .ZN(n62) );
  INV_X1 U215 ( .A(n78), .ZN(n70) );
  INV_X1 U216 ( .A(n89), .ZN(n79) );
  INV_X1 U217 ( .A(n102), .ZN(n101) );
  INV_X1 U218 ( .A(n104), .ZN(n100) );
  INV_X1 U219 ( .A(n106), .ZN(n108) );
  INV_X1 U220 ( .A(n120), .ZN(n112) );
  INV_X1 U221 ( .A(n4), .ZN(n133) );
  INV_X1 U222 ( .A(n137), .ZN(n138) );
  INV_X1 U223 ( .A(n149), .ZN(n148) );
  INV_X1 U224 ( .A(n155), .ZN(n154) );
  INV_X1 U225 ( .A(n28), .ZN(n157) );
endmodule


module SeqMult_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND4_X1 U3 ( .A1(n49), .A2(n15), .A3(n50), .A4(n51), .ZN(n1) );
  NAND2_X1 U4 ( .A1(n8), .A2(n9), .ZN(n2) );
  OR2_X1 U5 ( .A1(n54), .A2(n52), .ZN(n3) );
  NOR2_X1 U6 ( .A1(n3), .A2(n53), .ZN(n64) );
  NOR2_X1 U7 ( .A1(B[13]), .A2(n63), .ZN(n62) );
  XOR2_X1 U8 ( .A(n63), .B(B[13]), .Z(DIFF[13]) );
  NOR2_X1 U9 ( .A1(n3), .A2(B[8]), .ZN(n8) );
  NOR2_X1 U10 ( .A1(B[5]), .A2(n4), .ZN(n11) );
  NOR2_X1 U11 ( .A1(B[10]), .A2(n2), .ZN(n68) );
  AND2_X1 U12 ( .A1(n23), .A2(n22), .ZN(n20) );
  AND2_X1 U13 ( .A1(n44), .A2(n43), .ZN(n41) );
  AND2_X1 U14 ( .A1(n42), .A2(n41), .ZN(n39) );
  AND2_X1 U15 ( .A1(n40), .A2(n39), .ZN(n37) );
  AND2_X1 U16 ( .A1(n38), .A2(n37), .ZN(n35) );
  AND2_X1 U17 ( .A1(n36), .A2(n35), .ZN(n33) );
  AND2_X1 U18 ( .A1(n34), .A2(n33), .ZN(n31) );
  AND2_X1 U19 ( .A1(n32), .A2(n31), .ZN(n29) );
  AND2_X1 U20 ( .A1(n46), .A2(n45), .ZN(n43) );
  AND2_X1 U21 ( .A1(n47), .A2(n6), .ZN(n45) );
  OR2_X1 U22 ( .A1(n54), .A2(B[4]), .ZN(n4) );
  INV_X1 U23 ( .A(n54), .ZN(n15) );
  AND2_X1 U24 ( .A1(n11), .A2(n12), .ZN(n5) );
  NAND2_X1 U25 ( .A1(n64), .A2(n57), .ZN(n63) );
  NAND2_X1 U26 ( .A1(n62), .A2(n59), .ZN(n61) );
  NOR2_X1 U27 ( .A1(n55), .A2(n56), .ZN(n49) );
  AND2_X1 U28 ( .A1(n30), .A2(n29), .ZN(n27) );
  AND2_X1 U29 ( .A1(n28), .A2(n27), .ZN(n25) );
  AND2_X1 U30 ( .A1(n26), .A2(n25), .ZN(n22) );
  AND2_X1 U31 ( .A1(n1), .A2(n48), .ZN(n6) );
  NAND2_X1 U32 ( .A1(n20), .A2(n21), .ZN(n19) );
  NAND2_X1 U33 ( .A1(n57), .A2(n58), .ZN(n56) );
  NAND2_X1 U34 ( .A1(n59), .A2(n60), .ZN(n55) );
  XOR2_X1 U35 ( .A(\B[0] ), .B(B[1]), .Z(DIFF[1]) );
  XNOR2_X1 U36 ( .A(n61), .B(n60), .ZN(DIFF[15]) );
  XOR2_X1 U37 ( .A(n20), .B(n21), .Z(DIFF[30]) );
  XOR2_X1 U38 ( .A(n8), .B(n9), .Z(DIFF[9]) );
  XOR2_X1 U39 ( .A(n5), .B(n10), .Z(DIFF[7]) );
  XOR2_X1 U40 ( .A(n4), .B(B[5]), .Z(DIFF[5]) );
  XOR2_X1 U41 ( .A(n7), .B(n16), .Z(DIFF[3]) );
  XOR2_X1 U42 ( .A(n39), .B(n40), .Z(DIFF[21]) );
  XOR2_X1 U43 ( .A(n68), .B(n65), .Z(DIFF[11]) );
  XOR2_X1 U44 ( .A(n2), .B(B[10]), .Z(DIFF[10]) );
  XOR2_X1 U45 ( .A(n15), .B(n14), .Z(DIFF[4]) );
  XOR2_X1 U46 ( .A(n41), .B(n42), .Z(DIFF[20]) );
  XOR2_X1 U47 ( .A(n45), .B(n46), .Z(DIFF[18]) );
  XOR2_X1 U48 ( .A(n6), .B(n47), .Z(DIFF[17]) );
  XOR2_X1 U49 ( .A(n25), .B(n26), .Z(DIFF[28]) );
  XOR2_X1 U50 ( .A(n27), .B(n28), .Z(DIFF[27]) );
  XOR2_X1 U51 ( .A(n29), .B(n30), .Z(DIFF[26]) );
  XOR2_X1 U52 ( .A(n35), .B(n36), .Z(DIFF[23]) );
  XOR2_X1 U53 ( .A(n33), .B(n34), .Z(DIFF[24]) );
  XOR2_X1 U54 ( .A(n22), .B(n23), .Z(DIFF[29]) );
  XOR2_X1 U55 ( .A(n31), .B(n32), .Z(DIFF[25]) );
  XOR2_X1 U56 ( .A(n11), .B(n12), .Z(DIFF[6]) );
  XOR2_X1 U57 ( .A(n18), .B(n24), .Z(DIFF[2]) );
  XOR2_X1 U58 ( .A(n64), .B(n57), .Z(DIFF[12]) );
  XOR2_X1 U59 ( .A(n3), .B(B[8]), .Z(DIFF[8]) );
  XOR2_X1 U60 ( .A(n37), .B(n38), .Z(DIFF[22]) );
  XOR2_X1 U61 ( .A(n43), .B(n44), .Z(DIFF[19]) );
  XOR2_X1 U62 ( .A(B[31]), .B(n19), .Z(DIFF[31]) );
  INV_X1 U63 ( .A(B[12]), .ZN(n57) );
  INV_X1 U64 ( .A(B[14]), .ZN(n59) );
  NOR2_X1 U65 ( .A1(B[1]), .A2(\B[0] ), .ZN(n24) );
  INV_X1 U66 ( .A(B[1]), .ZN(n17) );
  INV_X1 U67 ( .A(B[9]), .ZN(n9) );
  INV_X1 U68 ( .A(B[4]), .ZN(n14) );
  INV_X1 U69 ( .A(B[2]), .ZN(n18) );
  INV_X1 U70 ( .A(B[6]), .ZN(n12) );
  INV_X1 U71 ( .A(B[30]), .ZN(n21) );
  AND3_X1 U72 ( .A1(n69), .A2(n17), .A3(n18), .ZN(n7) );
  INV_X1 U73 ( .A(B[13]), .ZN(n58) );
  INV_X1 U74 ( .A(B[15]), .ZN(n60) );
  INV_X1 U75 ( .A(B[19]), .ZN(n44) );
  INV_X1 U76 ( .A(B[18]), .ZN(n46) );
  INV_X1 U77 ( .A(B[17]), .ZN(n47) );
  INV_X1 U78 ( .A(B[29]), .ZN(n23) );
  INV_X1 U79 ( .A(B[28]), .ZN(n26) );
  INV_X1 U80 ( .A(B[27]), .ZN(n28) );
  INV_X1 U81 ( .A(B[26]), .ZN(n30) );
  INV_X1 U82 ( .A(B[25]), .ZN(n32) );
  INV_X1 U83 ( .A(B[24]), .ZN(n34) );
  INV_X1 U84 ( .A(B[23]), .ZN(n36) );
  INV_X1 U85 ( .A(B[22]), .ZN(n38) );
  INV_X1 U86 ( .A(B[21]), .ZN(n40) );
  INV_X1 U87 ( .A(B[20]), .ZN(n42) );
  INV_X1 U88 ( .A(B[16]), .ZN(n48) );
  INV_X1 U89 ( .A(B[3]), .ZN(n16) );
  INV_X1 U90 ( .A(B[7]), .ZN(n10) );
  INV_X1 U91 ( .A(B[11]), .ZN(n65) );
  INV_X1 U92 ( .A(B[5]), .ZN(n13) );
  INV_X1 U93 ( .A(B[8]), .ZN(n67) );
  INV_X1 U94 ( .A(B[10]), .ZN(n66) );
  INV_X1 U95 ( .A(\B[0] ), .ZN(n69) );
  NAND4_X1 U96 ( .A1(n65), .A2(n66), .A3(n9), .A4(n67), .ZN(n53) );
  NAND4_X1 U97 ( .A1(n17), .A2(n69), .A3(n18), .A4(n16), .ZN(n54) );
  NAND4_X1 U98 ( .A1(n10), .A2(n12), .A3(n13), .A4(n14), .ZN(n52) );
  XNOR2_X1 U99 ( .A(n1), .B(B[16]), .ZN(DIFF[16]) );
  INV_X1 U100 ( .A(n52), .ZN(n51) );
  INV_X1 U101 ( .A(n53), .ZN(n50) );
  XNOR2_X1 U102 ( .A(n62), .B(B[14]), .ZN(DIFF[14]) );
endmodule


module SeqMult_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207;

  AOI21_X1 U2 ( .B1(n103), .B2(n104), .A(n11), .ZN(n10) );
  AND2_X1 U3 ( .A1(n202), .A2(n122), .ZN(SUM[0]) );
  OAI21_X1 U4 ( .B1(n116), .B2(n117), .A(n118), .ZN(n2) );
  INV_X1 U5 ( .A(n169), .ZN(n3) );
  XOR2_X1 U6 ( .A(n164), .B(n4), .Z(SUM[15]) );
  AND2_X1 U7 ( .A1(n144), .A2(n143), .ZN(n4) );
  OAI21_X1 U8 ( .B1(n149), .B2(n169), .A(n151), .ZN(n5) );
  OAI21_X1 U9 ( .B1(n46), .B2(n163), .A(n195), .ZN(n6) );
  XNOR2_X1 U10 ( .A(n10), .B(n7), .ZN(SUM[24]) );
  AND2_X1 U11 ( .A1(n101), .A2(n100), .ZN(n7) );
  INV_X1 U12 ( .A(n102), .ZN(n11) );
  OAI21_X1 U13 ( .B1(n99), .B2(n10), .A(n100), .ZN(n8) );
  INV_X1 U14 ( .A(n83), .ZN(n14) );
  INV_X1 U15 ( .A(n117), .ZN(n9) );
  INV_X1 U16 ( .A(n13), .ZN(n80) );
  INV_X1 U17 ( .A(n125), .ZN(n12) );
  AOI21_X1 U18 ( .B1(n85), .B2(n84), .A(n14), .ZN(n13) );
  XOR2_X1 U19 ( .A(n17), .B(n15), .Z(SUM[22]) );
  NAND2_X1 U20 ( .A1(n108), .A2(n107), .ZN(n15) );
  OR2_X1 U21 ( .A1(B[6]), .A2(A[6]), .ZN(n39) );
  OR2_X1 U22 ( .A1(B[15]), .A2(A[15]), .ZN(n144) );
  OAI21_X1 U23 ( .B1(n46), .B2(n163), .A(n195), .ZN(n27) );
  NAND2_X1 U24 ( .A1(n70), .A2(n68), .ZN(n77) );
  NAND2_X1 U25 ( .A1(n146), .A2(n148), .ZN(n168) );
  NAND2_X1 U26 ( .A1(n178), .A2(n191), .ZN(n192) );
  NAND2_X1 U27 ( .A1(n171), .A2(n151), .ZN(n172) );
  NAND2_X1 U28 ( .A1(n153), .A2(n155), .ZN(n176) );
  NAND2_X1 U29 ( .A1(n139), .A2(n136), .ZN(n140) );
  NAND2_X1 U30 ( .A1(n81), .A2(n79), .ZN(n82) );
  NAND2_X1 U31 ( .A1(n85), .A2(n83), .ZN(n86) );
  NAND2_X1 U32 ( .A1(n33), .A2(n34), .ZN(n32) );
  NAND2_X1 U33 ( .A1(n29), .A2(n30), .ZN(n28) );
  NAND2_X1 U34 ( .A1(n91), .A2(n89), .ZN(n92) );
  NAND2_X1 U35 ( .A1(n97), .A2(n95), .ZN(n98) );
  NAND2_X1 U36 ( .A1(n104), .A2(n102), .ZN(n105) );
  NAND2_X1 U37 ( .A1(n120), .A2(n118), .ZN(n123) );
  NAND2_X1 U38 ( .A1(n128), .A2(n126), .ZN(n129) );
  NAND2_X1 U39 ( .A1(n134), .A2(n132), .ZN(n135) );
  NAND2_X1 U40 ( .A1(n62), .A2(n64), .ZN(n65) );
  INV_X1 U41 ( .A(n144), .ZN(n142) );
  INV_X1 U42 ( .A(n148), .ZN(n147) );
  XNOR2_X1 U43 ( .A(n43), .B(n45), .ZN(SUM[5]) );
  XNOR2_X1 U44 ( .A(n38), .B(n40), .ZN(SUM[6]) );
  NAND2_X1 U45 ( .A1(n39), .A2(n37), .ZN(n40) );
  XNOR2_X1 U46 ( .A(n75), .B(n121), .ZN(SUM[1]) );
  XNOR2_X1 U47 ( .A(n58), .B(n71), .ZN(SUM[2]) );
  NAND2_X1 U48 ( .A1(n72), .A2(n57), .ZN(n71) );
  NAND2_X1 U49 ( .A1(n53), .A2(n54), .ZN(n52) );
  INV_X1 U50 ( .A(n155), .ZN(n154) );
  OAI21_X1 U51 ( .B1(n156), .B2(n157), .A(n158), .ZN(n152) );
  INV_X1 U52 ( .A(n122), .ZN(n75) );
  XOR2_X1 U53 ( .A(n59), .B(n60), .Z(SUM[31]) );
  INV_X1 U54 ( .A(B[31]), .ZN(n60) );
  OR2_X1 U55 ( .A1(B[2]), .A2(A[2]), .ZN(n72) );
  NAND2_X1 U56 ( .A1(B[14]), .A2(A[14]), .ZN(n148) );
  NAND2_X1 U57 ( .A1(B[12]), .A2(A[12]), .ZN(n155) );
  OR2_X2 U58 ( .A1(B[10]), .A2(A[10]), .ZN(n178) );
  NAND2_X1 U59 ( .A1(B[28]), .A2(A[28]), .ZN(n79) );
  NAND2_X1 U60 ( .A1(B[17]), .A2(A[17]), .ZN(n132) );
  NAND2_X1 U61 ( .A1(B[25]), .A2(A[25]), .ZN(n95) );
  NAND2_X1 U62 ( .A1(B[29]), .A2(A[29]), .ZN(n68) );
  NAND2_X1 U63 ( .A1(B[16]), .A2(A[16]), .ZN(n136) );
  OR2_X1 U64 ( .A1(B[20]), .A2(A[20]), .ZN(n114) );
  OR2_X1 U65 ( .A1(B[14]), .A2(A[14]), .ZN(n146) );
  OR2_X1 U66 ( .A1(B[12]), .A2(A[12]), .ZN(n153) );
  OR2_X1 U67 ( .A1(B[7]), .A2(A[7]), .ZN(n33) );
  NAND2_X1 U68 ( .A1(B[30]), .A2(A[30]), .ZN(n64) );
  NAND2_X1 U69 ( .A1(B[26]), .A2(A[26]), .ZN(n89) );
  NAND2_X1 U70 ( .A1(B[19]), .A2(A[19]), .ZN(n118) );
  NAND2_X1 U71 ( .A1(B[24]), .A2(A[24]), .ZN(n100) );
  NAND2_X1 U72 ( .A1(B[23]), .A2(A[23]), .ZN(n102) );
  NAND2_X1 U73 ( .A1(B[27]), .A2(A[27]), .ZN(n83) );
  NAND2_X1 U74 ( .A1(B[15]), .A2(A[15]), .ZN(n143) );
  NAND2_X1 U75 ( .A1(B[22]), .A2(A[22]), .ZN(n107) );
  OR2_X1 U76 ( .A1(B[5]), .A2(A[5]), .ZN(n44) );
  OR2_X1 U77 ( .A1(B[4]), .A2(A[4]), .ZN(n49) );
  OR2_X1 U78 ( .A1(B[29]), .A2(A[29]), .ZN(n70) );
  OR2_X1 U79 ( .A1(B[28]), .A2(A[28]), .ZN(n81) );
  OR2_X1 U80 ( .A1(B[17]), .A2(A[17]), .ZN(n134) );
  OR2_X1 U81 ( .A1(B[25]), .A2(A[25]), .ZN(n97) );
  OR2_X1 U82 ( .A1(B[19]), .A2(A[19]), .ZN(n120) );
  OR2_X1 U83 ( .A1(B[26]), .A2(A[26]), .ZN(n91) );
  OR2_X1 U84 ( .A1(B[24]), .A2(A[24]), .ZN(n101) );
  OR2_X1 U85 ( .A1(B[27]), .A2(A[27]), .ZN(n85) );
  OR2_X1 U86 ( .A1(B[23]), .A2(A[23]), .ZN(n104) );
  OR2_X1 U87 ( .A1(B[22]), .A2(A[22]), .ZN(n108) );
  OR2_X1 U88 ( .A1(B[16]), .A2(A[16]), .ZN(n139) );
  OR2_X1 U89 ( .A1(B[30]), .A2(A[30]), .ZN(n62) );
  OR2_X1 U90 ( .A1(B[3]), .A2(A[3]), .ZN(n53) );
  OR2_X1 U91 ( .A1(B[18]), .A2(A[18]), .ZN(n128) );
  OR2_X1 U92 ( .A1(B[13]), .A2(A[13]), .ZN(n171) );
  INV_X1 U93 ( .A(A[0]), .ZN(n207) );
  OR2_X1 U94 ( .A1(B[11]), .A2(A[11]), .ZN(n179) );
  OR2_X1 U95 ( .A1(B[8]), .A2(A[8]), .ZN(n29) );
  OR2_X1 U96 ( .A1(B[21]), .A2(A[21]), .ZN(n111) );
  NAND2_X1 U97 ( .A1(n206), .A2(n207), .ZN(n202) );
  OAI21_X1 U98 ( .B1(n99), .B2(n10), .A(n100), .ZN(n96) );
  NAND2_X1 U99 ( .A1(n114), .A2(n113), .ZN(n115) );
  INV_X1 U100 ( .A(n113), .ZN(n22) );
  NAND2_X1 U101 ( .A1(B[20]), .A2(A[20]), .ZN(n113) );
  XNOR2_X1 U102 ( .A(n138), .B(n140), .ZN(SUM[16]) );
  OAI21_X1 U103 ( .B1(n141), .B2(n142), .A(n143), .ZN(n138) );
  NAND2_X1 U104 ( .A1(n111), .A2(n109), .ZN(n112) );
  INV_X1 U105 ( .A(n109), .ZN(n18) );
  NAND2_X1 U106 ( .A1(B[21]), .A2(A[21]), .ZN(n109) );
  XNOR2_X1 U107 ( .A(n9), .B(n123), .ZN(SUM[19]) );
  OAI21_X1 U108 ( .B1(n124), .B2(n125), .A(n126), .ZN(n119) );
  XNOR2_X1 U109 ( .A(n187), .B(n188), .ZN(SUM[11]) );
  XNOR2_X1 U110 ( .A(n69), .B(n77), .ZN(SUM[29]) );
  OAI21_X1 U111 ( .B1(n78), .B2(n13), .A(n79), .ZN(n69) );
  OR2_X1 U112 ( .A1(B[9]), .A2(A[9]), .ZN(n25) );
  NAND2_X1 U113 ( .A1(B[2]), .A2(A[2]), .ZN(n57) );
  OR2_X1 U114 ( .A1(B[1]), .A2(A[1]), .ZN(n76) );
  NAND2_X1 U115 ( .A1(B[10]), .A2(A[10]), .ZN(n191) );
  NAND2_X1 U116 ( .A1(B[3]), .A2(A[3]), .ZN(n54) );
  NAND2_X1 U117 ( .A1(B[13]), .A2(A[13]), .ZN(n151) );
  NAND2_X1 U118 ( .A1(B[18]), .A2(A[18]), .ZN(n126) );
  NAND2_X1 U119 ( .A1(B[8]), .A2(A[8]), .ZN(n30) );
  NAND2_X1 U120 ( .A1(B[11]), .A2(A[11]), .ZN(n183) );
  NAND2_X1 U121 ( .A1(n41), .A2(n42), .ZN(n38) );
  OAI21_X1 U122 ( .B1(n46), .B2(n47), .A(n48), .ZN(n43) );
  NAND2_X1 U123 ( .A1(n49), .A2(n48), .ZN(n50) );
  NAND2_X1 U124 ( .A1(B[7]), .A2(A[7]), .ZN(n34) );
  NAND2_X1 U125 ( .A1(B[4]), .A2(A[4]), .ZN(n48) );
  NAND2_X1 U126 ( .A1(B[6]), .A2(A[6]), .ZN(n37) );
  INV_X1 U127 ( .A(n25), .ZN(n16) );
  NAND2_X1 U128 ( .A1(B[9]), .A2(A[9]), .ZN(n26) );
  NAND2_X1 U129 ( .A1(n73), .A2(n74), .ZN(n58) );
  INV_X1 U130 ( .A(B[0]), .ZN(n206) );
  OAI21_X1 U131 ( .B1(n106), .B2(n17), .A(n107), .ZN(n103) );
  AOI21_X1 U132 ( .B1(n111), .B2(n110), .A(n18), .ZN(n17) );
  NAND2_X1 U133 ( .A1(B[0]), .A2(A[0]), .ZN(n122) );
  NOR2_X1 U134 ( .A1(B[1]), .A2(A[1]), .ZN(n19) );
  INV_X1 U135 ( .A(n21), .ZN(n110) );
  OAI21_X1 U136 ( .B1(n173), .B2(n174), .A(n155), .ZN(n170) );
  OAI21_X1 U137 ( .B1(n149), .B2(n169), .A(n151), .ZN(n167) );
  XNOR2_X1 U138 ( .A(n23), .B(n24), .ZN(SUM[9]) );
  NAND2_X1 U139 ( .A1(n30), .A2(n194), .ZN(n23) );
  XNOR2_X1 U140 ( .A(n175), .B(n176), .ZN(SUM[12]) );
  OAI21_X1 U141 ( .B1(n193), .B2(n186), .A(n26), .ZN(n20) );
  OAI21_X1 U142 ( .B1(n193), .B2(n186), .A(n26), .ZN(n190) );
  AOI21_X1 U143 ( .B1(n2), .B2(n114), .A(n22), .ZN(n21) );
  OAI21_X1 U144 ( .B1(n93), .B2(n94), .A(n95), .ZN(n90) );
  OAI21_X1 U145 ( .B1(n130), .B2(n131), .A(n132), .ZN(n127) );
  NAND2_X1 U146 ( .A1(n136), .A2(n137), .ZN(n133) );
  NAND2_X1 U147 ( .A1(n138), .A2(n139), .ZN(n137) );
  AOI21_X1 U148 ( .B1(n184), .B2(n178), .A(n185), .ZN(n182) );
  OAI21_X1 U149 ( .B1(n16), .B2(n30), .A(n26), .ZN(n184) );
  OAI21_X1 U150 ( .B1(n200), .B2(n48), .A(n41), .ZN(n198) );
  AOI21_X1 U151 ( .B1(n198), .B2(n39), .A(n199), .ZN(n197) );
  AOI21_X1 U152 ( .B1(n204), .B2(n72), .A(n205), .ZN(n203) );
  OAI21_X1 U153 ( .B1(n19), .B2(n122), .A(n73), .ZN(n204) );
  OAI21_X1 U154 ( .B1(n66), .B2(n67), .A(n68), .ZN(n61) );
  NAND2_X1 U155 ( .A1(n25), .A2(n26), .ZN(n24) );
  NAND4_X1 U156 ( .A1(n25), .A2(n29), .A3(n178), .A4(n179), .ZN(n157) );
  NAND2_X1 U157 ( .A1(n44), .A2(n41), .ZN(n45) );
  NAND2_X1 U158 ( .A1(n43), .A2(n44), .ZN(n42) );
  NAND4_X1 U159 ( .A1(n44), .A2(n49), .A3(n39), .A4(n33), .ZN(n163) );
  XNOR2_X1 U160 ( .A(n161), .B(n50), .ZN(SUM[4]) );
  NAND2_X1 U161 ( .A1(n158), .A2(n177), .ZN(n175) );
  XNOR2_X1 U162 ( .A(n84), .B(n86), .ZN(SUM[27]) );
  XNOR2_X1 U163 ( .A(n110), .B(n112), .ZN(SUM[21]) );
  XNOR2_X1 U164 ( .A(n133), .B(n135), .ZN(SUM[17]) );
  OAI21_X1 U165 ( .B1(n182), .B2(n181), .A(n183), .ZN(n180) );
  XNOR2_X1 U166 ( .A(n90), .B(n92), .ZN(SUM[26]) );
  OAI21_X1 U167 ( .B1(n87), .B2(n88), .A(n89), .ZN(n84) );
  AOI21_X1 U168 ( .B1(n145), .B2(n146), .A(n147), .ZN(n141) );
  NAND2_X1 U169 ( .A1(B[5]), .A2(A[5]), .ZN(n41) );
  XNOR2_X1 U170 ( .A(n61), .B(n65), .ZN(SUM[30]) );
  AOI21_X1 U171 ( .B1(n61), .B2(n62), .A(n63), .ZN(n59) );
  XNOR2_X1 U172 ( .A(n96), .B(n98), .ZN(SUM[25]) );
  XNOR2_X1 U173 ( .A(n103), .B(n105), .ZN(SUM[23]) );
  XNOR2_X1 U174 ( .A(n2), .B(n115), .ZN(SUM[20]) );
  XNOR2_X1 U175 ( .A(n12), .B(n129), .ZN(SUM[18]) );
  OAI21_X1 U176 ( .B1(n149), .B2(n150), .A(n151), .ZN(n145) );
  XNOR2_X1 U177 ( .A(n80), .B(n82), .ZN(SUM[28]) );
  AOI21_X1 U178 ( .B1(n152), .B2(n153), .A(n154), .ZN(n150) );
  XNOR2_X1 U179 ( .A(n167), .B(n168), .ZN(SUM[14]) );
  XNOR2_X1 U180 ( .A(n3), .B(n172), .ZN(SUM[13]) );
  NAND2_X1 U181 ( .A1(n76), .A2(n73), .ZN(n121) );
  NAND2_X1 U182 ( .A1(n75), .A2(n76), .ZN(n74) );
  OAI21_X1 U183 ( .B1(n197), .B2(n196), .A(n34), .ZN(n162) );
  AOI21_X1 U184 ( .B1(n159), .B2(n161), .A(n162), .ZN(n156) );
  XNOR2_X1 U185 ( .A(n20), .B(n192), .ZN(SUM[10]) );
  XNOR2_X1 U186 ( .A(n27), .B(n28), .ZN(SUM[8]) );
  AOI21_X1 U187 ( .B1(n190), .B2(n178), .A(n185), .ZN(n187) );
  NAND2_X1 U188 ( .A1(n160), .A2(n27), .ZN(n177) );
  NAND2_X1 U189 ( .A1(n29), .A2(n6), .ZN(n194) );
  OAI21_X1 U190 ( .B1(n201), .B2(n203), .A(n54), .ZN(n161) );
  NAND2_X1 U191 ( .A1(B[1]), .A2(A[1]), .ZN(n73) );
  XNOR2_X1 U192 ( .A(n31), .B(n32), .ZN(SUM[7]) );
  OAI21_X1 U193 ( .B1(n35), .B2(n36), .A(n37), .ZN(n31) );
  INV_X1 U194 ( .A(n38), .ZN(n36) );
  INV_X1 U195 ( .A(n39), .ZN(n35) );
  INV_X1 U196 ( .A(n49), .ZN(n47) );
  XNOR2_X1 U197 ( .A(n51), .B(n52), .ZN(SUM[3]) );
  OAI21_X1 U198 ( .B1(n55), .B2(n56), .A(n57), .ZN(n51) );
  INV_X1 U199 ( .A(n58), .ZN(n56) );
  INV_X1 U200 ( .A(n64), .ZN(n63) );
  INV_X1 U201 ( .A(n69), .ZN(n67) );
  INV_X1 U202 ( .A(n70), .ZN(n66) );
  INV_X1 U203 ( .A(n81), .ZN(n78) );
  INV_X1 U204 ( .A(n90), .ZN(n88) );
  INV_X1 U205 ( .A(n91), .ZN(n87) );
  INV_X1 U206 ( .A(n8), .ZN(n94) );
  INV_X1 U207 ( .A(n97), .ZN(n93) );
  INV_X1 U208 ( .A(n101), .ZN(n99) );
  INV_X1 U209 ( .A(n108), .ZN(n106) );
  INV_X1 U210 ( .A(n119), .ZN(n117) );
  INV_X1 U211 ( .A(n120), .ZN(n116) );
  INV_X1 U212 ( .A(n127), .ZN(n125) );
  INV_X1 U213 ( .A(n128), .ZN(n124) );
  INV_X1 U214 ( .A(n133), .ZN(n131) );
  INV_X1 U215 ( .A(n134), .ZN(n130) );
  INV_X1 U216 ( .A(n163), .ZN(n159) );
  OAI21_X1 U217 ( .B1(n165), .B2(n166), .A(n148), .ZN(n164) );
  INV_X1 U218 ( .A(n5), .ZN(n166) );
  INV_X1 U219 ( .A(n146), .ZN(n165) );
  INV_X1 U220 ( .A(n170), .ZN(n169) );
  INV_X1 U221 ( .A(n171), .ZN(n149) );
  INV_X1 U222 ( .A(n175), .ZN(n174) );
  INV_X1 U223 ( .A(n153), .ZN(n173) );
  INV_X1 U224 ( .A(n157), .ZN(n160) );
  INV_X1 U225 ( .A(n180), .ZN(n158) );
  NOR2_X1 U226 ( .A1(n189), .A2(n181), .ZN(n188) );
  INV_X1 U227 ( .A(n179), .ZN(n181) );
  INV_X1 U228 ( .A(n183), .ZN(n189) );
  INV_X1 U229 ( .A(n191), .ZN(n185) );
  INV_X1 U230 ( .A(n25), .ZN(n186) );
  INV_X1 U231 ( .A(n23), .ZN(n193) );
  INV_X1 U232 ( .A(n162), .ZN(n195) );
  INV_X1 U233 ( .A(n37), .ZN(n199) );
  INV_X1 U234 ( .A(n44), .ZN(n200) );
  INV_X1 U235 ( .A(n33), .ZN(n196) );
  INV_X1 U236 ( .A(n161), .ZN(n46) );
  INV_X1 U237 ( .A(n72), .ZN(n55) );
  INV_X1 U238 ( .A(n57), .ZN(n205) );
  INV_X1 U239 ( .A(n53), .ZN(n201) );
endmodule


module SeqMult_DW01_sub_6 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;

  AND4_X1 U3 ( .A1(n28), .A2(n63), .A3(n31), .A4(n44), .ZN(n12) );
  INV_X1 U4 ( .A(n8), .ZN(n19) );
  NAND2_X1 U5 ( .A1(n35), .A2(n34), .ZN(n1) );
  NAND2_X1 U6 ( .A1(n39), .A2(n38), .ZN(n2) );
  NAND2_X1 U7 ( .A1(n37), .A2(n36), .ZN(n3) );
  NAND2_X1 U8 ( .A1(n43), .A2(n42), .ZN(n4) );
  NAND2_X1 U9 ( .A1(n46), .A2(n45), .ZN(n5) );
  NAND2_X1 U10 ( .A1(n54), .A2(n58), .ZN(n6) );
  NAND2_X1 U11 ( .A1(n41), .A2(n40), .ZN(n7) );
  NAND2_X1 U12 ( .A1(n12), .A2(n9), .ZN(n8) );
  AND4_X1 U13 ( .A1(n21), .A2(n23), .A3(n25), .A4(n27), .ZN(n9) );
  AND4_X1 U14 ( .A1(n21), .A2(n23), .A3(n25), .A4(n27), .ZN(n10) );
  AND4_X1 U15 ( .A1(n59), .A2(n60), .A3(n18), .A4(n20), .ZN(n11) );
  XOR2_X1 U16 ( .A(n56), .B(B[15]), .Z(DIFF[15]) );
  XOR2_X1 U17 ( .A(n13), .B(n28), .Z(DIFF[3]) );
  NOR2_X1 U18 ( .A1(B[2]), .A2(n29), .ZN(n13) );
  XOR2_X1 U19 ( .A(B[31]), .B(n14), .Z(DIFF[31]) );
  NAND2_X1 U20 ( .A1(n32), .A2(n33), .ZN(n14) );
  NOR2_X1 U21 ( .A1(n8), .A2(n55), .ZN(n58) );
  NAND4_X1 U22 ( .A1(n59), .A2(n60), .A3(n18), .A4(n20), .ZN(n55) );
  NOR2_X1 U23 ( .A1(B[13]), .A2(n6), .ZN(n57) );
  NOR2_X1 U24 ( .A1(n26), .A2(B[4]), .ZN(n24) );
  NOR2_X1 U25 ( .A1(B[15]), .A2(n50), .ZN(n48) );
  NAND2_X1 U26 ( .A1(n51), .A2(n52), .ZN(n50) );
  NOR2_X1 U27 ( .A1(B[13]), .A2(n53), .ZN(n51) );
  NAND2_X1 U28 ( .A1(n16), .A2(n54), .ZN(n53) );
  NOR2_X1 U29 ( .A1(B[29]), .A2(n1), .ZN(n32) );
  XOR2_X1 U30 ( .A(n17), .B(n18), .Z(DIFF[9]) );
  XOR2_X1 U31 ( .A(n19), .B(n20), .Z(DIFF[8]) );
  XOR2_X1 U32 ( .A(n24), .B(n25), .Z(DIFF[5]) );
  XOR2_X1 U33 ( .A(n12), .B(n27), .Z(DIFF[4]) );
  NOR2_X1 U34 ( .A1(n8), .A2(B[8]), .ZN(n17) );
  NOR2_X1 U35 ( .A1(B[17]), .A2(n47), .ZN(n45) );
  NOR2_X1 U36 ( .A1(B[19]), .A2(n5), .ZN(n42) );
  NOR2_X1 U37 ( .A1(B[21]), .A2(n4), .ZN(n40) );
  NOR2_X1 U38 ( .A1(B[23]), .A2(n7), .ZN(n38) );
  NOR2_X1 U39 ( .A1(B[25]), .A2(n2), .ZN(n36) );
  NOR2_X1 U40 ( .A1(B[27]), .A2(n3), .ZN(n34) );
  XOR2_X1 U41 ( .A(n15), .B(n23), .Z(DIFF[6]) );
  NAND2_X1 U42 ( .A1(n48), .A2(n49), .ZN(n47) );
  AND2_X1 U43 ( .A1(n24), .A2(n25), .ZN(n15) );
  XOR2_X1 U44 ( .A(n4), .B(B[21]), .Z(DIFF[21]) );
  XOR2_X1 U45 ( .A(n5), .B(B[19]), .Z(DIFF[19]) );
  XOR2_X1 U46 ( .A(n45), .B(n46), .Z(DIFF[18]) );
  XOR2_X1 U47 ( .A(n62), .B(n60), .Z(DIFF[10]) );
  XOR2_X1 U48 ( .A(n6), .B(B[13]), .Z(DIFF[13]) );
  XOR2_X1 U49 ( .A(n38), .B(n39), .Z(DIFF[24]) );
  XOR2_X1 U50 ( .A(n58), .B(n54), .Z(DIFF[12]) );
  XOR2_X1 U51 ( .A(n7), .B(B[23]), .Z(DIFF[23]) );
  XOR2_X1 U52 ( .A(n34), .B(n35), .Z(DIFF[28]) );
  XOR2_X1 U53 ( .A(n40), .B(n41), .Z(DIFF[22]) );
  XOR2_X1 U54 ( .A(n42), .B(n43), .Z(DIFF[20]) );
  XOR2_X1 U55 ( .A(n47), .B(B[17]), .Z(DIFF[17]) );
  XOR2_X1 U56 ( .A(n32), .B(n33), .Z(DIFF[30]) );
  XOR2_X1 U57 ( .A(n36), .B(n37), .Z(DIFF[26]) );
  XOR2_X1 U58 ( .A(n1), .B(B[29]), .Z(DIFF[29]) );
  XOR2_X1 U59 ( .A(n2), .B(B[25]), .Z(DIFF[25]) );
  XOR2_X1 U60 ( .A(n3), .B(B[27]), .Z(DIFF[27]) );
  XOR2_X1 U61 ( .A(n48), .B(n49), .Z(DIFF[16]) );
  NAND2_X1 U62 ( .A1(n57), .A2(n52), .ZN(n56) );
  XOR2_X1 U63 ( .A(n30), .B(n31), .Z(DIFF[2]) );
  AND2_X1 U64 ( .A1(n17), .A2(n18), .ZN(n62) );
  NAND2_X1 U65 ( .A1(n15), .A2(n23), .ZN(n22) );
  AND3_X1 U66 ( .A1(n10), .A2(n11), .A3(n12), .ZN(n16) );
  XNOR2_X1 U67 ( .A(n22), .B(n21), .ZN(DIFF[7]) );
  XNOR2_X1 U68 ( .A(n61), .B(n59), .ZN(DIFF[11]) );
  NOR2_X1 U69 ( .A1(B[0]), .A2(B[1]), .ZN(n30) );
  XOR2_X1 U70 ( .A(B[0]), .B(B[1]), .Z(DIFF[1]) );
  INV_X1 U71 ( .A(B[5]), .ZN(n25) );
  INV_X1 U72 ( .A(B[14]), .ZN(n52) );
  INV_X1 U73 ( .A(B[6]), .ZN(n23) );
  INV_X1 U74 ( .A(B[8]), .ZN(n20) );
  INV_X1 U75 ( .A(B[4]), .ZN(n27) );
  INV_X1 U76 ( .A(B[9]), .ZN(n18) );
  INV_X1 U77 ( .A(B[12]), .ZN(n54) );
  INV_X1 U78 ( .A(B[10]), .ZN(n60) );
  INV_X1 U79 ( .A(B[2]), .ZN(n31) );
  INV_X1 U80 ( .A(B[16]), .ZN(n49) );
  INV_X1 U81 ( .A(B[7]), .ZN(n21) );
  INV_X1 U82 ( .A(B[11]), .ZN(n59) );
  INV_X1 U83 ( .A(B[18]), .ZN(n46) );
  INV_X1 U84 ( .A(B[20]), .ZN(n43) );
  INV_X1 U85 ( .A(B[22]), .ZN(n41) );
  INV_X1 U86 ( .A(B[24]), .ZN(n39) );
  INV_X1 U87 ( .A(B[26]), .ZN(n37) );
  INV_X1 U88 ( .A(B[3]), .ZN(n28) );
  INV_X1 U89 ( .A(B[1]), .ZN(n44) );
  INV_X1 U90 ( .A(B[30]), .ZN(n33) );
  INV_X1 U91 ( .A(B[28]), .ZN(n35) );
  NAND2_X1 U92 ( .A1(n62), .A2(n60), .ZN(n61) );
  INV_X1 U93 ( .A(B[0]), .ZN(n63) );
  INV_X1 U94 ( .A(n30), .ZN(n29) );
  XNOR2_X1 U95 ( .A(n57), .B(B[14]), .ZN(DIFF[14]) );
  INV_X1 U96 ( .A(n12), .ZN(n26) );
endmodule


module SeqMult ( clk, internalClk, rst, A, B, P );
  input [31:0] A;
  input [31:0] B;
  output [63:0] P;
  input clk, internalClk, rst;
  wire   N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163,
         N164, N165, N166, N167, N168, N169, N170, N171, N172, N205, N206,
         N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N235, N236, N303, N304, N305,
         N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316,
         N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327,
         N328, N329, N330, N331, N332, N333, N334, N337, N338, N339, N340,
         N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351,
         N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362,
         N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373,
         N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384,
         N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395,
         N396, N397, N398, N399, N400, N465, N466, N467, N468, N469, N470,
         N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503,
         N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514,
         N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525,
         N526, N527, N528, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584,
         N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595,
         N596, N829, N831, N833, N835, N837, N839, N841, N843, N845, N847,
         N849, N851, N853, N855, N857, N859, N861, N863, N865, N867, N869,
         N871, N873, N875, N877, N879, N881, N883, N885, N887, N889, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688,
         N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677,
         N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666,
         \dp_cluster_0/N268 , n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969;
  wire   [31:0] counter;
  wire   [31:0] A_reg;
  wire   [31:0] B_reg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  DFF_X1 \A_reg_reg[31]  ( .D(N40), .CK(clk), .Q(A_reg[31]), .QN(n407) );
  DFF_X1 \A_reg_reg[30]  ( .D(N39), .CK(clk), .Q(A_reg[30]), .QN(n341) );
  DFF_X1 \A_reg_reg[29]  ( .D(N38), .CK(clk), .Q(A_reg[29]), .QN(n343) );
  DFF_X1 \A_reg_reg[28]  ( .D(N37), .CK(clk), .Q(A_reg[28]), .QN(n345) );
  DFF_X1 \A_reg_reg[27]  ( .D(N36), .CK(clk), .Q(A_reg[27]), .QN(n347) );
  DFF_X1 \A_reg_reg[26]  ( .D(N35), .CK(clk), .Q(A_reg[26]), .QN(n349) );
  DFF_X1 \A_reg_reg[25]  ( .D(N34), .CK(clk), .Q(A_reg[25]), .QN(n351) );
  DFF_X1 \A_reg_reg[24]  ( .D(N33), .CK(clk), .Q(A_reg[24]), .QN(n353) );
  DFF_X1 \A_reg_reg[23]  ( .D(N32), .CK(clk), .Q(A_reg[23]), .QN(n355) );
  DFF_X1 \A_reg_reg[22]  ( .D(N31), .CK(clk), .Q(A_reg[22]), .QN(n357) );
  DFF_X1 \A_reg_reg[21]  ( .D(N30), .CK(clk), .Q(A_reg[21]), .QN(n359) );
  DFF_X1 \A_reg_reg[20]  ( .D(N29), .CK(clk), .Q(A_reg[20]), .QN(n361) );
  DFF_X1 \A_reg_reg[19]  ( .D(N28), .CK(clk), .Q(A_reg[19]), .QN(n363) );
  DFF_X1 \A_reg_reg[18]  ( .D(N27), .CK(clk), .Q(A_reg[18]), .QN(n365) );
  DFF_X1 \A_reg_reg[17]  ( .D(N26), .CK(clk), .Q(A_reg[17]), .QN(n367) );
  DFF_X1 \A_reg_reg[16]  ( .D(N25), .CK(clk), .Q(A_reg[16]), .QN(n369) );
  DFF_X1 \A_reg_reg[15]  ( .D(N24), .CK(clk), .Q(A_reg[15]), .QN(n371) );
  DFF_X1 \A_reg_reg[14]  ( .D(N23), .CK(clk), .Q(A_reg[14]), .QN(n373) );
  DFF_X1 \A_reg_reg[13]  ( .D(N22), .CK(clk), .Q(A_reg[13]), .QN(n375) );
  DFF_X1 \A_reg_reg[12]  ( .D(N21), .CK(clk), .Q(A_reg[12]), .QN(n377) );
  DFF_X1 \A_reg_reg[11]  ( .D(N20), .CK(clk), .Q(A_reg[11]), .QN(n379) );
  DFF_X1 \A_reg_reg[10]  ( .D(N19), .CK(clk), .Q(A_reg[10]), .QN(n381) );
  DFF_X1 \A_reg_reg[9]  ( .D(N18), .CK(clk), .Q(A_reg[9]), .QN(n383) );
  DFF_X1 \A_reg_reg[8]  ( .D(N17), .CK(clk), .Q(A_reg[8]), .QN(n385) );
  DFF_X1 \A_reg_reg[7]  ( .D(N16), .CK(clk), .Q(A_reg[7]), .QN(n387) );
  DFF_X1 \A_reg_reg[6]  ( .D(N15), .CK(clk), .Q(A_reg[6]), .QN(n389) );
  DFF_X1 \A_reg_reg[5]  ( .D(N14), .CK(clk), .Q(A_reg[5]), .QN(n391) );
  DFF_X1 \A_reg_reg[4]  ( .D(N13), .CK(clk), .Q(A_reg[4]), .QN(n393) );
  DFF_X1 \A_reg_reg[3]  ( .D(N12), .CK(clk), .Q(A_reg[3]), .QN(n395) );
  DFF_X1 \A_reg_reg[2]  ( .D(N11), .CK(clk), .Q(A_reg[2]), .QN(n397) );
  DFF_X1 \A_reg_reg[1]  ( .D(N10), .CK(clk), .Q(A_reg[1]), .QN(n399) );
  DFF_X1 \A_reg_reg[0]  ( .D(N9), .CK(clk), .Q(A_reg[0]), .QN(n406) );
  DFF_X1 \B_reg_reg[31]  ( .D(N72), .CK(clk), .Q(B_reg[31]), .QN(n338) );
  DFF_X1 \B_reg_reg[30]  ( .D(N71), .CK(clk), .Q(B_reg[30]) );
  DFF_X1 \B_reg_reg[29]  ( .D(N70), .CK(clk), .Q(B_reg[29]) );
  DFF_X1 \B_reg_reg[28]  ( .D(N69), .CK(clk), .Q(B_reg[28]) );
  DFF_X1 \B_reg_reg[27]  ( .D(N68), .CK(clk), .Q(B_reg[27]) );
  DFF_X1 \B_reg_reg[26]  ( .D(N67), .CK(clk), .Q(B_reg[26]) );
  DFF_X1 \B_reg_reg[25]  ( .D(N66), .CK(clk), .Q(B_reg[25]) );
  DFF_X1 \B_reg_reg[24]  ( .D(N65), .CK(clk), .Q(B_reg[24]) );
  DFF_X1 \B_reg_reg[23]  ( .D(N64), .CK(clk), .Q(B_reg[23]) );
  DFF_X1 \B_reg_reg[22]  ( .D(N63), .CK(clk), .Q(B_reg[22]) );
  DFF_X1 \B_reg_reg[21]  ( .D(N62), .CK(clk), .Q(B_reg[21]) );
  DFF_X1 \B_reg_reg[20]  ( .D(N61), .CK(clk), .Q(B_reg[20]) );
  DFF_X1 \B_reg_reg[19]  ( .D(N60), .CK(clk), .Q(B_reg[19]) );
  DFF_X1 \B_reg_reg[18]  ( .D(N59), .CK(clk), .Q(B_reg[18]) );
  DFF_X1 \B_reg_reg[17]  ( .D(N58), .CK(clk), .Q(B_reg[17]) );
  DFF_X1 \B_reg_reg[16]  ( .D(N57), .CK(clk), .Q(B_reg[16]) );
  DFF_X1 \B_reg_reg[15]  ( .D(N56), .CK(clk), .Q(B_reg[15]) );
  DFF_X1 \B_reg_reg[14]  ( .D(N55), .CK(clk), .Q(B_reg[14]) );
  DFF_X1 \B_reg_reg[13]  ( .D(N54), .CK(clk), .Q(B_reg[13]) );
  DFF_X1 \B_reg_reg[12]  ( .D(N53), .CK(clk), .Q(B_reg[12]) );
  DFF_X1 \B_reg_reg[11]  ( .D(N52), .CK(clk), .Q(B_reg[11]) );
  DFF_X1 \B_reg_reg[10]  ( .D(N51), .CK(clk), .Q(B_reg[10]) );
  DFF_X1 \B_reg_reg[9]  ( .D(N50), .CK(clk), .Q(B_reg[9]) );
  DFF_X1 \B_reg_reg[8]  ( .D(N49), .CK(clk), .Q(B_reg[8]) );
  DFF_X1 \B_reg_reg[7]  ( .D(N48), .CK(clk), .Q(B_reg[7]) );
  DFF_X1 \B_reg_reg[6]  ( .D(N47), .CK(clk), .Q(B_reg[6]) );
  DFF_X1 \B_reg_reg[5]  ( .D(N46), .CK(clk), .Q(B_reg[5]) );
  DFF_X1 \B_reg_reg[4]  ( .D(N45), .CK(clk), .Q(B_reg[4]) );
  DFF_X1 \B_reg_reg[3]  ( .D(N44), .CK(clk), .Q(B_reg[3]) );
  DFF_X1 \B_reg_reg[2]  ( .D(N43), .CK(clk), .Q(B_reg[2]) );
  DFF_X1 \B_reg_reg[1]  ( .D(N42), .CK(clk), .Q(B_reg[1]) );
  DFF_X1 \B_reg_reg[0]  ( .D(N41), .CK(clk), .Q(B_reg[0]) );
  DFFR_X1 \counter_reg[0]  ( .D(N497), .CK(internalClk), .RN(n794), .Q(
        counter[0]), .QN(n405) );
  DFFR_X1 \counter_reg[1]  ( .D(N498), .CK(internalClk), .RN(n795), .Q(
        counter[1]), .QN(n404) );
  DFFR_X1 \counter_reg[2]  ( .D(N499), .CK(internalClk), .RN(n796), .Q(
        counter[2]), .QN(n403) );
  DFFR_X1 \counter_reg[3]  ( .D(N500), .CK(internalClk), .RN(n795), .Q(
        counter[3]) );
  DFFR_X1 \counter_reg[4]  ( .D(N501), .CK(internalClk), .RN(n791), .Q(
        counter[4]) );
  DFFR_X1 \counter_reg[5]  ( .D(N502), .CK(internalClk), .RN(n793), .Q(
        counter[5]), .QN(n242) );
  DFFR_X1 \counter_reg[6]  ( .D(N503), .CK(internalClk), .RN(n793), .Q(
        counter[6]), .QN(n712) );
  DFFR_X1 \counter_reg[7]  ( .D(N504), .CK(internalClk), .RN(n791), .Q(
        counter[7]), .QN(n240) );
  DFFR_X1 \counter_reg[8]  ( .D(N505), .CK(internalClk), .RN(n792), .Q(
        counter[8]), .QN(n711) );
  DFFR_X1 \counter_reg[9]  ( .D(N506), .CK(internalClk), .RN(n794), .Q(
        counter[9]), .QN(n710) );
  DFFR_X1 \counter_reg[10]  ( .D(N507), .CK(internalClk), .RN(n791), .Q(
        counter[10]), .QN(n231) );
  DFFR_X1 \counter_reg[11]  ( .D(N508), .CK(internalClk), .RN(n792), .Q(
        counter[11]), .QN(n229) );
  DFFR_X1 \counter_reg[12]  ( .D(N509), .CK(internalClk), .RN(n791), .Q(
        counter[12]), .QN(n230) );
  DFFR_X1 \counter_reg[13]  ( .D(N510), .CK(internalClk), .RN(n791), .Q(
        counter[13]) );
  DFFR_X1 \counter_reg[14]  ( .D(N511), .CK(internalClk), .RN(n795), .Q(
        counter[14]) );
  DFFR_X1 \counter_reg[15]  ( .D(N512), .CK(internalClk), .RN(n792), .Q(
        counter[15]) );
  DFFR_X1 \counter_reg[16]  ( .D(N513), .CK(internalClk), .RN(n793), .Q(
        counter[16]), .QN(n235) );
  DFFR_X1 \counter_reg[17]  ( .D(N514), .CK(internalClk), .RN(n792), .Q(
        counter[17]), .QN(n233) );
  DFFR_X1 \counter_reg[18]  ( .D(N515), .CK(internalClk), .RN(n794), .Q(
        counter[18]), .QN(n234) );
  DFFR_X1 \counter_reg[19]  ( .D(N516), .CK(internalClk), .RN(n795), .Q(
        counter[19]) );
  DFFR_X1 \counter_reg[20]  ( .D(N517), .CK(internalClk), .RN(n792), .Q(
        counter[20]), .QN(n232) );
  DFFR_X1 \counter_reg[21]  ( .D(N518), .CK(internalClk), .RN(n791), .Q(
        counter[21]) );
  DFFR_X1 \counter_reg[22]  ( .D(N519), .CK(internalClk), .RN(n795), .Q(
        counter[22]) );
  DFFR_X1 \counter_reg[23]  ( .D(N520), .CK(internalClk), .RN(n794), .Q(
        counter[23]), .QN(n239) );
  DFFR_X1 \counter_reg[24]  ( .D(N521), .CK(internalClk), .RN(n793), .Q(
        counter[24]), .QN(n237) );
  DFFR_X1 \counter_reg[25]  ( .D(N522), .CK(internalClk), .RN(n795), .Q(
        counter[25]), .QN(n238) );
  DFFR_X1 \counter_reg[26]  ( .D(N523), .CK(internalClk), .RN(n794), .Q(
        counter[26]), .QN(n715) );
  DFFR_X1 \counter_reg[27]  ( .D(N524), .CK(internalClk), .RN(n793), .Q(
        counter[27]), .QN(n236) );
  DFFR_X1 \counter_reg[28]  ( .D(N525), .CK(internalClk), .RN(n792), .Q(
        counter[28]), .QN(n714) );
  DFFR_X1 \counter_reg[29]  ( .D(N526), .CK(internalClk), .RN(n793), .Q(
        counter[29]), .QN(n713) );
  DFFR_X1 \counter_reg[30]  ( .D(N527), .CK(internalClk), .RN(n794), .Q(
        counter[30]), .QN(n243) );
  DFFR_X1 \counter_reg[31]  ( .D(N528), .CK(internalClk), .RN(n796), .Q(
        counter[31]), .QN(n241) );
  DFF_X1 \P_reg[63]  ( .D(N596), .CK(clk), .Q(P[63]) );
  DFF_X1 \P_reg[62]  ( .D(N595), .CK(clk), .Q(P[62]) );
  DFF_X1 \P_reg[61]  ( .D(N594), .CK(clk), .Q(P[61]) );
  DFF_X1 \P_reg[60]  ( .D(N593), .CK(clk), .Q(P[60]) );
  DFF_X1 \P_reg[59]  ( .D(N592), .CK(clk), .Q(P[59]) );
  DFF_X1 \P_reg[58]  ( .D(N591), .CK(clk), .Q(P[58]) );
  DFF_X1 \P_reg[57]  ( .D(N590), .CK(clk), .Q(P[57]) );
  DFF_X1 \P_reg[56]  ( .D(N589), .CK(clk), .Q(P[56]) );
  DFF_X1 \P_reg[55]  ( .D(N588), .CK(clk), .Q(P[55]) );
  DFF_X1 \P_reg[54]  ( .D(N587), .CK(clk), .Q(P[54]) );
  DFF_X1 \P_reg[53]  ( .D(N586), .CK(clk), .Q(P[53]) );
  DFF_X1 \P_reg[52]  ( .D(N585), .CK(clk), .Q(P[52]) );
  DFF_X1 \P_reg[51]  ( .D(N584), .CK(clk), .Q(P[51]) );
  DFF_X1 \P_reg[50]  ( .D(N583), .CK(clk), .Q(P[50]) );
  DFF_X1 \P_reg[49]  ( .D(N582), .CK(clk), .Q(P[49]) );
  DFF_X1 \P_reg[48]  ( .D(N581), .CK(clk), .Q(P[48]) );
  DFF_X1 \P_reg[47]  ( .D(N580), .CK(clk), .Q(P[47]) );
  DFF_X1 \P_reg[46]  ( .D(N579), .CK(clk), .Q(P[46]) );
  DFF_X1 \P_reg[45]  ( .D(N578), .CK(clk), .Q(P[45]) );
  DFF_X1 \P_reg[44]  ( .D(N577), .CK(clk), .Q(P[44]) );
  DFF_X1 \P_reg[43]  ( .D(N576), .CK(clk), .Q(P[43]) );
  DFF_X1 \P_reg[42]  ( .D(N575), .CK(clk), .Q(P[42]) );
  DFF_X1 \P_reg[41]  ( .D(N574), .CK(clk), .Q(P[41]) );
  DFF_X1 \P_reg[40]  ( .D(N573), .CK(clk), .Q(P[40]) );
  DFF_X1 \P_reg[39]  ( .D(N572), .CK(clk), .Q(P[39]) );
  DFF_X1 \P_reg[38]  ( .D(N571), .CK(clk), .Q(P[38]) );
  DFF_X1 \P_reg[37]  ( .D(N570), .CK(clk), .Q(P[37]) );
  DFF_X1 \P_reg[36]  ( .D(N569), .CK(clk), .Q(P[36]) );
  DFF_X1 \P_reg[35]  ( .D(N568), .CK(clk), .Q(P[35]) );
  DFF_X1 \P_reg[34]  ( .D(N567), .CK(clk), .Q(P[34]) );
  DFF_X1 \P_reg[33]  ( .D(N566), .CK(clk), .Q(P[33]) );
  DFF_X1 \P_reg[32]  ( .D(N565), .CK(clk), .Q(P[32]) );
  DFF_X1 \P_reg[31]  ( .D(N564), .CK(clk), .Q(P[31]) );
  DFF_X1 \P_reg[30]  ( .D(N563), .CK(clk), .Q(P[30]) );
  DFF_X1 \P_reg[29]  ( .D(N562), .CK(clk), .Q(P[29]) );
  DFF_X1 \P_reg[28]  ( .D(N561), .CK(clk), .Q(P[28]) );
  DFF_X1 \P_reg[27]  ( .D(N560), .CK(clk), .Q(P[27]) );
  DFF_X1 \P_reg[26]  ( .D(N559), .CK(clk), .Q(P[26]) );
  DFF_X1 \P_reg[25]  ( .D(N558), .CK(clk), .Q(P[25]) );
  DFF_X1 \P_reg[24]  ( .D(N557), .CK(clk), .Q(P[24]) );
  DFF_X1 \P_reg[23]  ( .D(N556), .CK(clk), .Q(P[23]) );
  DFF_X1 \P_reg[22]  ( .D(N555), .CK(clk), .Q(P[22]) );
  DFF_X1 \P_reg[21]  ( .D(N554), .CK(clk), .Q(P[21]) );
  DFF_X1 \P_reg[20]  ( .D(N553), .CK(clk), .Q(P[20]) );
  DFF_X1 \P_reg[19]  ( .D(N552), .CK(clk), .Q(P[19]) );
  DFF_X1 \P_reg[18]  ( .D(N551), .CK(clk), .Q(P[18]) );
  DFF_X1 \P_reg[17]  ( .D(N550), .CK(clk), .Q(P[17]) );
  DFF_X1 \P_reg[16]  ( .D(N549), .CK(clk), .Q(P[16]) );
  DFF_X1 \P_reg[15]  ( .D(N548), .CK(clk), .Q(P[15]) );
  DFF_X1 \P_reg[14]  ( .D(N547), .CK(clk), .Q(P[14]) );
  DFF_X1 \P_reg[13]  ( .D(N546), .CK(clk), .Q(P[13]) );
  DFF_X1 \P_reg[12]  ( .D(N545), .CK(clk), .Q(P[12]) );
  DFF_X1 \P_reg[11]  ( .D(N544), .CK(clk), .Q(P[11]) );
  DFF_X1 \P_reg[10]  ( .D(N543), .CK(clk), .Q(P[10]) );
  DFF_X1 \P_reg[9]  ( .D(N542), .CK(clk), .Q(P[9]) );
  DFF_X1 \P_reg[8]  ( .D(N541), .CK(clk), .Q(P[8]) );
  DFF_X1 \P_reg[7]  ( .D(N540), .CK(clk), .Q(P[7]) );
  DFF_X1 \P_reg[6]  ( .D(N539), .CK(clk), .Q(P[6]) );
  DFF_X1 \P_reg[5]  ( .D(N538), .CK(clk), .Q(P[5]) );
  DFF_X1 \P_reg[4]  ( .D(N537), .CK(clk), .Q(P[4]) );
  DFF_X1 \P_reg[3]  ( .D(N536), .CK(clk), .Q(P[3]) );
  DFF_X1 \P_reg[2]  ( .D(N535), .CK(clk), .Q(P[2]) );
  DFF_X1 \P_reg[1]  ( .D(N534), .CK(clk), .Q(P[1]) );
  DFF_X1 \P_reg[0]  ( .D(N533), .CK(clk), .Q(P[0]) );
  DFF_X1 \multiplier_reg[31]  ( .D(n599), .CK(internalClk), .Q(n634) );
  DFF_X1 \Accumulator_reg[30]  ( .D(n598), .CK(internalClk), .Q(n638), .QN(
        n439) );
  DFF_X1 \Accumulator_reg[29]  ( .D(n597), .CK(internalClk), .Q(n639), .QN(
        n438) );
  DFF_X1 \Accumulator_reg[28]  ( .D(n596), .CK(internalClk), .Q(n640), .QN(
        n437) );
  DFF_X1 \Accumulator_reg[27]  ( .D(n595), .CK(internalClk), .Q(n641), .QN(
        n436) );
  DFF_X1 \Accumulator_reg[26]  ( .D(n594), .CK(internalClk), .Q(n642), .QN(
        n435) );
  DFF_X1 \Accumulator_reg[25]  ( .D(n593), .CK(internalClk), .Q(n643), .QN(
        n434) );
  DFF_X1 \Accumulator_reg[24]  ( .D(n592), .CK(internalClk), .Q(n644), .QN(
        n433) );
  DFF_X1 \Accumulator_reg[23]  ( .D(n591), .CK(internalClk), .Q(n645), .QN(
        n432) );
  DFF_X1 \Accumulator_reg[22]  ( .D(n590), .CK(internalClk), .Q(n646), .QN(
        n431) );
  DFF_X1 \Accumulator_reg[21]  ( .D(n589), .CK(internalClk), .Q(n647), .QN(
        n430) );
  DFF_X1 \Accumulator_reg[20]  ( .D(n588), .CK(internalClk), .Q(n648), .QN(
        n429) );
  DFF_X1 \Accumulator_reg[19]  ( .D(n587), .CK(internalClk), .Q(n649), .QN(
        n428) );
  DFF_X1 \Accumulator_reg[18]  ( .D(n586), .CK(internalClk), .Q(n650), .QN(
        n427) );
  DFF_X1 \Accumulator_reg[17]  ( .D(n585), .CK(internalClk), .Q(n651), .QN(
        n426) );
  DFF_X1 \Accumulator_reg[16]  ( .D(n584), .CK(internalClk), .Q(n652), .QN(
        n425) );
  DFF_X1 \Accumulator_reg[15]  ( .D(n583), .CK(internalClk), .Q(n653), .QN(
        n424) );
  DFF_X1 \Accumulator_reg[14]  ( .D(n582), .CK(internalClk), .Q(n654), .QN(
        n423) );
  DFF_X1 \Accumulator_reg[13]  ( .D(n581), .CK(internalClk), .Q(n655), .QN(
        n422) );
  DFF_X1 \Accumulator_reg[12]  ( .D(n580), .CK(internalClk), .Q(n656), .QN(
        n421) );
  DFF_X1 \Accumulator_reg[11]  ( .D(n579), .CK(internalClk), .Q(n657), .QN(
        n420) );
  DFF_X1 \Accumulator_reg[10]  ( .D(n578), .CK(internalClk), .Q(n658), .QN(
        n419) );
  DFF_X1 \Accumulator_reg[9]  ( .D(n577), .CK(internalClk), .Q(n659), .QN(n418) );
  DFF_X1 \Accumulator_reg[8]  ( .D(n576), .CK(internalClk), .Q(n660), .QN(n417) );
  DFF_X1 \Accumulator_reg[7]  ( .D(n575), .CK(internalClk), .Q(n661), .QN(n416) );
  DFF_X1 \Accumulator_reg[6]  ( .D(n574), .CK(internalClk), .Q(n662), .QN(n415) );
  DFF_X1 \Accumulator_reg[5]  ( .D(n573), .CK(internalClk), .Q(n663), .QN(n414) );
  DFF_X1 \Accumulator_reg[4]  ( .D(n572), .CK(internalClk), .Q(n664), .QN(n413) );
  DFF_X1 \Accumulator_reg[3]  ( .D(n571), .CK(internalClk), .Q(n665), .QN(n412) );
  DFF_X1 \Accumulator_reg[2]  ( .D(n570), .CK(internalClk), .Q(n666), .QN(n411) );
  DFF_X1 \Accumulator_reg[1]  ( .D(n569), .CK(internalClk), .Q(n667), .QN(n410) );
  DFF_X1 \Accumulator_reg[0]  ( .D(n568), .CK(internalClk), .Q(n668), .QN(n409) );
  DFF_X1 \multiplicand_reg[0]  ( .D(n567), .CK(internalClk), .QN(n408) );
  DFF_X1 \multiplicand_reg[1]  ( .D(n566), .CK(internalClk), .QN(n400) );
  DFF_X1 \multiplicand_reg[2]  ( .D(n565), .CK(internalClk), .QN(n398) );
  DFF_X1 \multiplicand_reg[3]  ( .D(n564), .CK(internalClk), .QN(n396) );
  DFF_X1 \multiplicand_reg[4]  ( .D(n563), .CK(internalClk), .QN(n394) );
  DFF_X1 \multiplicand_reg[5]  ( .D(n562), .CK(internalClk), .QN(n392) );
  DFF_X1 \multiplicand_reg[6]  ( .D(n561), .CK(internalClk), .QN(n390) );
  DFF_X1 \multiplicand_reg[7]  ( .D(n560), .CK(internalClk), .QN(n388) );
  DFF_X1 \multiplicand_reg[8]  ( .D(n559), .CK(internalClk), .QN(n386) );
  DFF_X1 \multiplicand_reg[9]  ( .D(n558), .CK(internalClk), .QN(n384) );
  DFF_X1 \multiplicand_reg[10]  ( .D(n557), .CK(internalClk), .QN(n382) );
  DFF_X1 \multiplicand_reg[11]  ( .D(n556), .CK(internalClk), .QN(n380) );
  DFF_X1 \multiplicand_reg[12]  ( .D(n555), .CK(internalClk), .QN(n378) );
  DFF_X1 \multiplicand_reg[13]  ( .D(n554), .CK(internalClk), .QN(n376) );
  DFF_X1 \multiplicand_reg[14]  ( .D(n553), .CK(internalClk), .QN(n374) );
  DFF_X1 \multiplicand_reg[15]  ( .D(n552), .CK(internalClk), .QN(n372) );
  DFF_X1 \multiplicand_reg[16]  ( .D(n551), .CK(internalClk), .QN(n370) );
  DFF_X1 \multiplicand_reg[17]  ( .D(n550), .CK(internalClk), .QN(n368) );
  DFF_X1 \multiplicand_reg[18]  ( .D(n549), .CK(internalClk), .QN(n366) );
  DFF_X1 \multiplicand_reg[19]  ( .D(n548), .CK(internalClk), .QN(n364) );
  DFF_X1 \multiplicand_reg[20]  ( .D(n547), .CK(internalClk), .QN(n362) );
  DFF_X1 \multiplicand_reg[21]  ( .D(n546), .CK(internalClk), .QN(n360) );
  DFF_X1 \multiplicand_reg[22]  ( .D(n545), .CK(internalClk), .QN(n358) );
  DFF_X1 \multiplicand_reg[23]  ( .D(n544), .CK(internalClk), .QN(n356) );
  DFF_X1 \multiplicand_reg[24]  ( .D(n543), .CK(internalClk), .QN(n354) );
  DFF_X1 \multiplicand_reg[25]  ( .D(n542), .CK(internalClk), .QN(n352) );
  DFF_X1 \multiplicand_reg[26]  ( .D(n541), .CK(internalClk), .QN(n350) );
  DFF_X1 \multiplicand_reg[27]  ( .D(n540), .CK(internalClk), .QN(n348) );
  DFF_X1 \multiplicand_reg[28]  ( .D(n539), .CK(internalClk), .QN(n346) );
  DFF_X1 \multiplicand_reg[29]  ( .D(n538), .CK(internalClk), .QN(n344) );
  DFF_X1 \multiplicand_reg[30]  ( .D(n537), .CK(internalClk), .QN(n342) );
  DFF_X1 \multiplicand_reg[31]  ( .D(n536), .CK(internalClk), .QN(n340) );
  DFF_X1 \multiplier_reg[30]  ( .D(n535), .CK(internalClk), .Q(n669), .QN(n339) );
  DFF_X1 \multiplier_reg[29]  ( .D(n534), .CK(internalClk), .Q(n670), .QN(n337) );
  DFF_X1 \multiplier_reg[28]  ( .D(n533), .CK(internalClk), .Q(n671), .QN(n336) );
  DFF_X1 \multiplier_reg[27]  ( .D(n532), .CK(internalClk), .Q(n672), .QN(n335) );
  DFF_X1 \multiplier_reg[26]  ( .D(n531), .CK(internalClk), .Q(n673), .QN(n334) );
  DFF_X1 \multiplier_reg[25]  ( .D(n530), .CK(internalClk), .Q(n674), .QN(n333) );
  DFF_X1 \multiplier_reg[24]  ( .D(n529), .CK(internalClk), .Q(n675), .QN(n332) );
  DFF_X1 \multiplier_reg[23]  ( .D(n528), .CK(internalClk), .Q(n676), .QN(n331) );
  DFF_X1 \multiplier_reg[22]  ( .D(n527), .CK(internalClk), .Q(n677), .QN(n330) );
  DFF_X1 \multiplier_reg[21]  ( .D(n526), .CK(internalClk), .Q(n678), .QN(n329) );
  DFF_X1 \multiplier_reg[20]  ( .D(n525), .CK(internalClk), .Q(n679), .QN(n328) );
  DFF_X1 \multiplier_reg[19]  ( .D(n524), .CK(internalClk), .Q(n680), .QN(n327) );
  DFF_X1 \multiplier_reg[18]  ( .D(n523), .CK(internalClk), .Q(n681), .QN(n326) );
  DFF_X1 \multiplier_reg[17]  ( .D(n522), .CK(internalClk), .Q(n682), .QN(n325) );
  DFF_X1 \multiplier_reg[16]  ( .D(n521), .CK(internalClk), .Q(n683), .QN(n324) );
  DFF_X1 \multiplier_reg[15]  ( .D(n520), .CK(internalClk), .Q(n684), .QN(n323) );
  DFF_X1 \multiplier_reg[14]  ( .D(n519), .CK(internalClk), .Q(n685), .QN(n322) );
  DFF_X1 \multiplier_reg[13]  ( .D(n518), .CK(internalClk), .Q(n686), .QN(n321) );
  DFF_X1 \multiplier_reg[12]  ( .D(n517), .CK(internalClk), .Q(n687), .QN(n320) );
  DFF_X1 \multiplier_reg[11]  ( .D(n516), .CK(internalClk), .Q(n688), .QN(n319) );
  DFF_X1 \multiplier_reg[10]  ( .D(n515), .CK(internalClk), .Q(n689), .QN(n318) );
  DFF_X1 \multiplier_reg[9]  ( .D(n514), .CK(internalClk), .Q(n690), .QN(n317)
         );
  DFF_X1 \multiplier_reg[8]  ( .D(n513), .CK(internalClk), .Q(n691), .QN(n316)
         );
  DFF_X1 \multiplier_reg[7]  ( .D(n512), .CK(internalClk), .Q(n692), .QN(n315)
         );
  DFF_X1 \multiplier_reg[6]  ( .D(n511), .CK(internalClk), .Q(n693), .QN(n314)
         );
  DFF_X1 \multiplier_reg[5]  ( .D(n510), .CK(internalClk), .Q(n694), .QN(n313)
         );
  DFF_X1 \multiplier_reg[4]  ( .D(n509), .CK(internalClk), .Q(n695), .QN(n312)
         );
  DFF_X1 \multiplier_reg[3]  ( .D(n508), .CK(internalClk), .Q(n696), .QN(n311)
         );
  DFF_X1 \multiplier_reg[2]  ( .D(n507), .CK(internalClk), .Q(n697), .QN(n310)
         );
  DFF_X1 \multiplier_reg[1]  ( .D(n506), .CK(internalClk), .Q(n698), .QN(n309)
         );
  DFF_X1 \P_reg_reg[31]  ( .D(n505), .CK(internalClk), .QN(n308) );
  DFF_X1 \P_reg_reg[32]  ( .D(n504), .CK(internalClk), .QN(n307) );
  DFF_X1 \P_reg_reg[33]  ( .D(n503), .CK(internalClk), .QN(n306) );
  DFF_X1 \P_reg_reg[34]  ( .D(n502), .CK(internalClk), .QN(n305) );
  DFF_X1 \P_reg_reg[35]  ( .D(n501), .CK(internalClk), .QN(n304) );
  DFF_X1 \P_reg_reg[36]  ( .D(n500), .CK(internalClk), .QN(n303) );
  DFF_X1 \P_reg_reg[37]  ( .D(n499), .CK(internalClk), .QN(n302) );
  DFF_X1 \P_reg_reg[38]  ( .D(n498), .CK(internalClk), .QN(n301) );
  DFF_X1 \P_reg_reg[39]  ( .D(n497), .CK(internalClk), .QN(n300) );
  DFF_X1 \P_reg_reg[40]  ( .D(n496), .CK(internalClk), .QN(n299) );
  DFF_X1 \P_reg_reg[41]  ( .D(n495), .CK(internalClk), .QN(n298) );
  DFF_X1 \P_reg_reg[42]  ( .D(n494), .CK(internalClk), .QN(n297) );
  DFF_X1 \P_reg_reg[43]  ( .D(n493), .CK(internalClk), .QN(n296) );
  DFF_X1 \P_reg_reg[44]  ( .D(n492), .CK(internalClk), .QN(n295) );
  DFF_X1 \P_reg_reg[45]  ( .D(n491), .CK(internalClk), .QN(n294) );
  DFF_X1 \P_reg_reg[46]  ( .D(n490), .CK(internalClk), .QN(n293) );
  DFF_X1 \P_reg_reg[47]  ( .D(n489), .CK(internalClk), .QN(n292) );
  DFF_X1 \P_reg_reg[48]  ( .D(n488), .CK(internalClk), .QN(n291) );
  DFF_X1 \P_reg_reg[49]  ( .D(n487), .CK(internalClk), .QN(n290) );
  DFF_X1 \P_reg_reg[50]  ( .D(n486), .CK(internalClk), .QN(n289) );
  DFF_X1 \P_reg_reg[51]  ( .D(n485), .CK(internalClk), .QN(n288) );
  DFF_X1 \P_reg_reg[52]  ( .D(n484), .CK(internalClk), .QN(n287) );
  DFF_X1 \P_reg_reg[53]  ( .D(n483), .CK(internalClk), .QN(n286) );
  DFF_X1 \P_reg_reg[54]  ( .D(n482), .CK(internalClk), .QN(n285) );
  DFF_X1 \P_reg_reg[55]  ( .D(n481), .CK(internalClk), .QN(n284) );
  DFF_X1 \P_reg_reg[56]  ( .D(n480), .CK(internalClk), .QN(n283) );
  DFF_X1 \P_reg_reg[57]  ( .D(n479), .CK(internalClk), .QN(n282) );
  DFF_X1 \P_reg_reg[58]  ( .D(n478), .CK(internalClk), .QN(n281) );
  DFF_X1 \P_reg_reg[59]  ( .D(n477), .CK(internalClk), .QN(n280) );
  DFF_X1 \P_reg_reg[60]  ( .D(n476), .CK(internalClk), .QN(n279) );
  DFF_X1 \P_reg_reg[61]  ( .D(n475), .CK(internalClk), .QN(n278) );
  DFF_X1 \P_reg_reg[62]  ( .D(n474), .CK(internalClk), .QN(n277) );
  DFF_X1 \P_reg_reg[63]  ( .D(n473), .CK(internalClk), .Q(n637), .QN(n276) );
  DFF_X1 \multiplier_reg[0]  ( .D(n472), .CK(internalClk), .Q(n699), .QN(n275)
         );
  DFF_X1 \P_reg_reg[0]  ( .D(n471), .CK(internalClk), .QN(n274) );
  DFF_X1 \P_reg_reg[1]  ( .D(n470), .CK(internalClk), .QN(n273) );
  DFF_X1 \P_reg_reg[2]  ( .D(n469), .CK(internalClk), .QN(n272) );
  DFF_X1 \P_reg_reg[3]  ( .D(n468), .CK(internalClk), .QN(n271) );
  DFF_X1 \P_reg_reg[4]  ( .D(n467), .CK(internalClk), .QN(n270) );
  DFF_X1 \P_reg_reg[5]  ( .D(n466), .CK(internalClk), .QN(n269) );
  DFF_X1 \P_reg_reg[6]  ( .D(n465), .CK(internalClk), .QN(n268) );
  DFF_X1 \P_reg_reg[7]  ( .D(n464), .CK(internalClk), .QN(n267) );
  DFF_X1 \P_reg_reg[8]  ( .D(n463), .CK(internalClk), .QN(n266) );
  DFF_X1 \P_reg_reg[9]  ( .D(n462), .CK(internalClk), .QN(n265) );
  DFF_X1 \P_reg_reg[10]  ( .D(n461), .CK(internalClk), .QN(n264) );
  DFF_X1 \P_reg_reg[11]  ( .D(n460), .CK(internalClk), .QN(n263) );
  DFF_X1 \P_reg_reg[12]  ( .D(n459), .CK(internalClk), .QN(n262) );
  DFF_X1 \P_reg_reg[13]  ( .D(n458), .CK(internalClk), .QN(n261) );
  DFF_X1 \P_reg_reg[14]  ( .D(n457), .CK(internalClk), .QN(n260) );
  DFF_X1 \P_reg_reg[15]  ( .D(n456), .CK(internalClk), .QN(n259) );
  DFF_X1 \P_reg_reg[16]  ( .D(n455), .CK(internalClk), .QN(n258) );
  DFF_X1 \P_reg_reg[17]  ( .D(n454), .CK(internalClk), .QN(n257) );
  DFF_X1 \P_reg_reg[18]  ( .D(n453), .CK(internalClk), .QN(n256) );
  DFF_X1 \P_reg_reg[19]  ( .D(n452), .CK(internalClk), .QN(n255) );
  DFF_X1 \P_reg_reg[20]  ( .D(n451), .CK(internalClk), .QN(n254) );
  DFF_X1 \P_reg_reg[21]  ( .D(n450), .CK(internalClk), .QN(n253) );
  DFF_X1 \P_reg_reg[22]  ( .D(n449), .CK(internalClk), .QN(n252) );
  DFF_X1 \P_reg_reg[23]  ( .D(n448), .CK(internalClk), .QN(n251) );
  DFF_X1 \P_reg_reg[24]  ( .D(n447), .CK(internalClk), .QN(n250) );
  DFF_X1 \P_reg_reg[25]  ( .D(n446), .CK(internalClk), .QN(n249) );
  DFF_X1 \P_reg_reg[26]  ( .D(n445), .CK(internalClk), .QN(n248) );
  DFF_X1 \P_reg_reg[27]  ( .D(n444), .CK(internalClk), .QN(n247) );
  DFF_X1 \P_reg_reg[28]  ( .D(n443), .CK(internalClk), .QN(n246) );
  DFF_X1 \P_reg_reg[29]  ( .D(n442), .CK(internalClk), .QN(n245) );
  DFF_X1 \P_reg_reg[30]  ( .D(n441), .CK(internalClk), .QN(n244) );
  SeqMult_DW01_inc_0 add_60 ( .A(counter), .SUM({N496, N495, N494, N493, N492, 
        N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, 
        N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, 
        N467, N466, N465}) );
  SeqMult_DW02_mult_0 mult_add_51_S2_aco ( .A({N205, N206, N207, N208, N209, 
        N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, 
        N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, 
        N234, N235, N236}), .B(\dp_cluster_0/N268 ), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, N697, N696, N695, N694, N693, N692, N691, 
        N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, 
        N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, 
        N666}) );
  SeqMult_DW01_sub_3 sub_59_S2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, N334, 
        N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, 
        N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, 
        N309, N308, N307, N306, N305, N304, N303, n969, n600, n601, n602, n603, 
        n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
        n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
        n628, n629}), .CI(1'b0), .DIFF({N400, N399, N398, N397, N396, N395, 
        N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, 
        N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, 
        N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, 
        N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, 
        N346, N345, N344, N343, N342, N341, N340, N339, N338, N337}) );
  SeqMult_DW01_sub_4 sub_46_S2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B(B_reg), .CI(1'b0), .DIFF({N172, N171, N170, N169, N168, 
        N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, 
        N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, 
        N143, N142, N141}) );
  SeqMult_DW01_add_1 add_51_S2_aco ( .A({1'b0, N829, N831, N833, N835, N837, 
        N839, N841, N843, N845, N847, N849, N851, N853, N855, N857, N859, N861, 
        N863, N865, N867, N869, N871, N873, N875, N877, N879, N881, N883, N885, 
        N887, N889}), .B({N697, N696, N695, N694, N693, N692, N691, N690, N689, 
        N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, 
        N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666}), 
        .CI(1'b0), .SUM({N334, N333, N332, N331, N330, N329, N328, N327, N326, 
        N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, 
        N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303}) );
  SeqMult_DW01_sub_6 sub_43_S2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B(A_reg), .CI(1'b0), .DIFF({N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, 
        SYNOPSYS_UNCONNECTED__1}) );
  AND3_X1 U642 ( .A1(n403), .A2(n404), .A3(n405), .ZN(n633) );
  AND2_X1 U643 ( .A1(n760), .A2(n902), .ZN(n635) );
  AND2_X1 U644 ( .A1(n760), .A2(n901), .ZN(n636) );
  NOR2_X1 U645 ( .A1(n824), .A2(n701), .ZN(n700) );
  NOR2_X1 U646 ( .A1(n824), .A2(n701), .ZN(n897) );
  NAND2_X1 U647 ( .A1(n703), .A2(n633), .ZN(n701) );
  CLKBUF_X1 U648 ( .A(n824), .Z(n702) );
  CLKBUF_X1 U649 ( .A(n742), .Z(n748) );
  NOR2_X1 U650 ( .A1(counter[3]), .A2(counter[4]), .ZN(n703) );
  NOR2_X1 U651 ( .A1(n824), .A2(n704), .ZN(n825) );
  INV_X1 U652 ( .A(n703), .ZN(n704) );
  BUF_X4 U653 ( .A(n744), .Z(n721) );
  OR2_X1 U654 ( .A1(n275), .A2(n742), .ZN(n705) );
  NAND2_X1 U655 ( .A1(n705), .A2(n862), .ZN(\dp_cluster_0/N268 ) );
  NAND2_X1 U656 ( .A1(n722), .A2(A_reg[31]), .ZN(n706) );
  NAND2_X1 U657 ( .A1(n722), .A2(A_reg[31]), .ZN(n707) );
  BUF_X2 U658 ( .A(n745), .Z(n722) );
  BUF_X1 U659 ( .A(n758), .Z(n760) );
  BUF_X1 U660 ( .A(n708), .Z(n736) );
  BUF_X1 U661 ( .A(n758), .Z(n761) );
  BUF_X1 U662 ( .A(n759), .Z(n764) );
  BUF_X1 U663 ( .A(n759), .Z(n763) );
  BUF_X1 U664 ( .A(n758), .Z(n762) );
  BUF_X1 U665 ( .A(n708), .Z(n737) );
  BUF_X1 U666 ( .A(n708), .Z(n738) );
  CLKBUF_X3 U667 ( .A(n742), .Z(n747) );
  INV_X1 U668 ( .A(n797), .ZN(n786) );
  INV_X1 U669 ( .A(n798), .ZN(n787) );
  INV_X1 U670 ( .A(n798), .ZN(n785) );
  INV_X1 U671 ( .A(n797), .ZN(n784) );
  INV_X1 U672 ( .A(n799), .ZN(n788) );
  BUF_X1 U673 ( .A(n766), .Z(n769) );
  BUF_X1 U674 ( .A(n766), .Z(n768) );
  BUF_X1 U675 ( .A(n767), .Z(n772) );
  BUF_X1 U676 ( .A(n767), .Z(n771) );
  BUF_X1 U677 ( .A(n766), .Z(n770) );
  BUF_X1 U678 ( .A(n750), .Z(n752) );
  BUF_X1 U679 ( .A(n750), .Z(n753) );
  BUF_X1 U680 ( .A(n750), .Z(n754) );
  BUF_X1 U681 ( .A(n751), .Z(n755) );
  BUF_X1 U682 ( .A(n751), .Z(n756) );
  AND2_X1 U683 ( .A1(n743), .A2(n799), .ZN(n708) );
  INV_X1 U684 ( .A(n797), .ZN(n782) );
  INV_X1 U685 ( .A(n799), .ZN(n783) );
  INV_X1 U686 ( .A(n798), .ZN(n789) );
  BUF_X1 U687 ( .A(n707), .Z(n720) );
  BUF_X1 U688 ( .A(n860), .Z(n726) );
  BUF_X1 U689 ( .A(n896), .Z(n739) );
  BUF_X1 U690 ( .A(n896), .Z(n740) );
  BUF_X1 U691 ( .A(n896), .Z(n741) );
  BUF_X1 U692 ( .A(n894), .Z(n734) );
  NAND2_X1 U693 ( .A1(n722), .A2(A_reg[31]), .ZN(n899) );
  BUF_X1 U694 ( .A(n893), .Z(n732) );
  BUF_X1 U695 ( .A(n893), .Z(n731) );
  INV_X1 U696 ( .A(n709), .ZN(n749) );
  BUF_X1 U697 ( .A(n893), .Z(n733) );
  BUF_X1 U698 ( .A(n781), .Z(n776) );
  BUF_X1 U699 ( .A(n780), .Z(n777) );
  BUF_X1 U700 ( .A(n780), .Z(n778) );
  BUF_X1 U701 ( .A(n780), .Z(n779) );
  BUF_X1 U702 ( .A(n781), .Z(n774) );
  BUF_X1 U703 ( .A(n781), .Z(n775) );
  NAND2_X1 U704 ( .A1(n407), .A2(n742), .ZN(n894) );
  AND4_X1 U705 ( .A1(n823), .A2(counter[4]), .A3(counter[3]), .A4(n822), .ZN(
        n709) );
  NOR2_X1 U706 ( .A1(n782), .A2(n273), .ZN(N534) );
  NOR2_X1 U707 ( .A1(n782), .A2(n272), .ZN(N535) );
  NOR2_X1 U708 ( .A1(n782), .A2(n271), .ZN(N536) );
  NOR2_X1 U709 ( .A1(n782), .A2(n270), .ZN(N537) );
  NOR2_X1 U710 ( .A1(n782), .A2(n269), .ZN(N538) );
  NOR2_X1 U711 ( .A1(n782), .A2(n268), .ZN(N539) );
  NOR2_X1 U712 ( .A1(n782), .A2(n267), .ZN(N540) );
  NOR2_X1 U713 ( .A1(n782), .A2(n266), .ZN(N541) );
  NOR2_X1 U714 ( .A1(n782), .A2(n265), .ZN(N542) );
  NOR2_X1 U715 ( .A1(n782), .A2(n264), .ZN(N543) );
  NOR2_X1 U716 ( .A1(n782), .A2(n263), .ZN(N544) );
  NOR2_X1 U717 ( .A1(n782), .A2(n262), .ZN(N545) );
  NOR2_X1 U718 ( .A1(n783), .A2(n261), .ZN(N546) );
  NOR2_X1 U719 ( .A1(n783), .A2(n260), .ZN(N547) );
  NOR2_X1 U720 ( .A1(n783), .A2(n259), .ZN(N548) );
  NOR2_X1 U721 ( .A1(n783), .A2(n258), .ZN(N549) );
  NOR2_X1 U722 ( .A1(n783), .A2(n257), .ZN(N550) );
  NOR2_X1 U723 ( .A1(n783), .A2(n256), .ZN(N551) );
  NOR2_X1 U724 ( .A1(n783), .A2(n255), .ZN(N552) );
  NOR2_X1 U725 ( .A1(n783), .A2(n254), .ZN(N553) );
  NOR2_X1 U726 ( .A1(n783), .A2(n253), .ZN(N554) );
  NOR2_X1 U727 ( .A1(n783), .A2(n252), .ZN(N555) );
  NOR2_X1 U728 ( .A1(n783), .A2(n251), .ZN(N556) );
  NOR2_X1 U729 ( .A1(n783), .A2(n250), .ZN(N557) );
  NOR2_X1 U730 ( .A1(n784), .A2(n274), .ZN(N533) );
  NOR2_X1 U731 ( .A1(n784), .A2(n249), .ZN(N558) );
  NOR2_X1 U732 ( .A1(n784), .A2(n248), .ZN(N559) );
  NOR2_X1 U733 ( .A1(n784), .A2(n247), .ZN(N560) );
  NOR2_X1 U734 ( .A1(n784), .A2(n246), .ZN(N561) );
  NOR2_X1 U735 ( .A1(n784), .A2(n245), .ZN(N562) );
  BUF_X1 U736 ( .A(rst), .Z(n781) );
  BUF_X1 U737 ( .A(rst), .Z(n780) );
  CLKBUF_X1 U738 ( .A(n700), .Z(n744) );
  NAND2_X1 U739 ( .A1(n407), .A2(n744), .ZN(n716) );
  NAND2_X1 U740 ( .A1(n407), .A2(n742), .ZN(n719) );
  NAND2_X1 U741 ( .A1(n722), .A2(A_reg[31]), .ZN(n717) );
  INV_X1 U742 ( .A(n829), .ZN(n718) );
  BUF_X1 U743 ( .A(n745), .Z(n723) );
  CLKBUF_X1 U744 ( .A(n894), .Z(n735) );
  BUF_X2 U745 ( .A(n700), .Z(n742) );
  BUF_X1 U746 ( .A(n700), .Z(n745) );
  INV_X1 U747 ( .A(n826), .ZN(n724) );
  CLKBUF_X1 U748 ( .A(n860), .Z(n727) );
  CLKBUF_X1 U749 ( .A(n861), .Z(n730) );
  CLKBUF_X1 U750 ( .A(n861), .Z(n728) );
  CLKBUF_X1 U751 ( .A(n861), .Z(n729) );
  CLKBUF_X1 U752 ( .A(N333), .Z(n725) );
  BUF_X2 U753 ( .A(n748), .Z(n743) );
  BUF_X2 U754 ( .A(n742), .Z(n746) );
  BUF_X1 U755 ( .A(n635), .Z(n750) );
  BUF_X1 U756 ( .A(n635), .Z(n751) );
  BUF_X1 U757 ( .A(n751), .Z(n757) );
  BUF_X1 U758 ( .A(n966), .Z(n758) );
  BUF_X1 U759 ( .A(n966), .Z(n759) );
  BUF_X1 U760 ( .A(n759), .Z(n765) );
  BUF_X1 U761 ( .A(n636), .Z(n766) );
  BUF_X1 U762 ( .A(n636), .Z(n767) );
  BUF_X1 U763 ( .A(n767), .Z(n773) );
  INV_X1 U764 ( .A(n796), .ZN(n790) );
  INV_X1 U765 ( .A(n774), .ZN(n791) );
  INV_X1 U766 ( .A(n774), .ZN(n792) );
  INV_X1 U767 ( .A(n774), .ZN(n793) );
  INV_X1 U768 ( .A(n774), .ZN(n794) );
  INV_X1 U769 ( .A(n775), .ZN(n795) );
  INV_X1 U770 ( .A(n776), .ZN(n796) );
  INV_X1 U771 ( .A(n776), .ZN(n797) );
  INV_X1 U772 ( .A(n776), .ZN(n798) );
  INV_X1 U773 ( .A(n776), .ZN(n799) );
  INV_X1 U774 ( .A(n776), .ZN(n800) );
  INV_X1 U775 ( .A(n777), .ZN(n801) );
  INV_X1 U776 ( .A(n777), .ZN(n802) );
  INV_X1 U777 ( .A(n777), .ZN(n803) );
  INV_X1 U778 ( .A(n777), .ZN(n804) );
  INV_X1 U779 ( .A(n777), .ZN(n805) );
  INV_X1 U780 ( .A(n778), .ZN(n806) );
  INV_X1 U781 ( .A(n778), .ZN(n807) );
  INV_X1 U782 ( .A(n778), .ZN(n808) );
  INV_X1 U783 ( .A(n778), .ZN(n809) );
  INV_X1 U784 ( .A(n778), .ZN(n810) );
  INV_X1 U785 ( .A(n779), .ZN(n811) );
  INV_X1 U786 ( .A(n779), .ZN(n812) );
  AND2_X1 U787 ( .A1(B[0]), .A2(n800), .ZN(N41) );
  INV_X1 U788 ( .A(B[31]), .ZN(n900) );
  NOR2_X1 U789 ( .A1(n788), .A2(n900), .ZN(N72) );
  NAND4_X1 U790 ( .A1(n241), .A2(n713), .A3(n714), .A4(n715), .ZN(n813) );
  NOR4_X1 U791 ( .A1(n813), .A2(counter[19]), .A3(counter[21]), .A4(
        counter[22]), .ZN(n821) );
  NAND3_X1 U792 ( .A1(n710), .A2(n711), .A3(n712), .ZN(n814) );
  NOR4_X1 U793 ( .A1(n814), .A2(counter[13]), .A3(counter[14]), .A4(
        counter[15]), .ZN(n820) );
  NAND3_X1 U794 ( .A1(n236), .A2(n238), .A3(n243), .ZN(n818) );
  NAND4_X1 U795 ( .A1(n232), .A2(n234), .A3(n237), .A4(n239), .ZN(n817) );
  NAND3_X1 U796 ( .A1(n235), .A2(n230), .A3(n233), .ZN(n816) );
  NAND4_X1 U797 ( .A1(n240), .A2(n242), .A3(n229), .A4(n231), .ZN(n815) );
  NOR4_X1 U798 ( .A1(n815), .A2(n817), .A3(n816), .A4(n818), .ZN(n819) );
  NAND3_X1 U799 ( .A1(n819), .A2(n820), .A3(n821), .ZN(n824) );
  INV_X1 U800 ( .A(n702), .ZN(n823) );
  NOR3_X1 U801 ( .A1(n405), .A2(n404), .A3(n403), .ZN(n822) );
  AND2_X1 U802 ( .A1(N470), .A2(n749), .ZN(N502) );
  AND2_X1 U803 ( .A1(N472), .A2(n749), .ZN(N504) );
  AND2_X1 U804 ( .A1(N475), .A2(n749), .ZN(N507) );
  AND2_X1 U805 ( .A1(N476), .A2(n749), .ZN(N508) );
  AND2_X1 U806 ( .A1(N477), .A2(n749), .ZN(N509) );
  AND2_X1 U807 ( .A1(N481), .A2(n749), .ZN(N513) );
  AND2_X1 U808 ( .A1(N482), .A2(n749), .ZN(N514) );
  AND2_X1 U809 ( .A1(N483), .A2(n749), .ZN(N515) );
  AND2_X1 U810 ( .A1(N485), .A2(n749), .ZN(N517) );
  AND2_X1 U811 ( .A1(N488), .A2(n749), .ZN(N520) );
  AND2_X1 U812 ( .A1(N489), .A2(n749), .ZN(N521) );
  AND2_X1 U813 ( .A1(N490), .A2(n749), .ZN(N522) );
  AND2_X1 U814 ( .A1(N492), .A2(n749), .ZN(N524) );
  AND2_X1 U815 ( .A1(N495), .A2(n749), .ZN(N527) );
  AND2_X1 U816 ( .A1(N494), .A2(n749), .ZN(N526) );
  AND2_X1 U817 ( .A1(N493), .A2(n749), .ZN(N525) );
  AND2_X1 U818 ( .A1(N491), .A2(n749), .ZN(N523) );
  AND2_X1 U819 ( .A1(N487), .A2(n749), .ZN(N519) );
  AND2_X1 U820 ( .A1(N486), .A2(n749), .ZN(N518) );
  AND2_X1 U821 ( .A1(N484), .A2(n749), .ZN(N516) );
  AND2_X1 U822 ( .A1(N480), .A2(n749), .ZN(N512) );
  AND2_X1 U823 ( .A1(N479), .A2(n749), .ZN(N511) );
  AND2_X1 U824 ( .A1(N478), .A2(n749), .ZN(N510) );
  AND2_X1 U825 ( .A1(N474), .A2(n749), .ZN(N506) );
  AND2_X1 U826 ( .A1(N473), .A2(n749), .ZN(N505) );
  AND2_X1 U827 ( .A1(N471), .A2(n749), .ZN(N503) );
  AND2_X1 U828 ( .A1(N469), .A2(n749), .ZN(N501) );
  AND2_X1 U829 ( .A1(N468), .A2(n749), .ZN(N500) );
  AND2_X1 U830 ( .A1(N467), .A2(n749), .ZN(N499) );
  AND2_X1 U831 ( .A1(N466), .A2(n749), .ZN(N498) );
  AND2_X1 U832 ( .A1(N496), .A2(n749), .ZN(N528) );
  AND2_X1 U833 ( .A1(N465), .A2(n749), .ZN(N497) );
  AND2_X1 U834 ( .A1(B[30]), .A2(n812), .ZN(N71) );
  AND2_X1 U835 ( .A1(B[29]), .A2(n812), .ZN(N70) );
  AND2_X1 U836 ( .A1(B[28]), .A2(n812), .ZN(N69) );
  AND2_X1 U837 ( .A1(B[27]), .A2(n812), .ZN(N68) );
  AND2_X1 U838 ( .A1(B[26]), .A2(n811), .ZN(N67) );
  AND2_X1 U839 ( .A1(B[25]), .A2(n811), .ZN(N66) );
  AND2_X1 U840 ( .A1(B[24]), .A2(n811), .ZN(N65) );
  AND2_X1 U841 ( .A1(B[23]), .A2(n811), .ZN(N64) );
  AND2_X1 U842 ( .A1(B[22]), .A2(n811), .ZN(N63) );
  AND2_X1 U843 ( .A1(B[21]), .A2(n810), .ZN(N62) );
  AND2_X1 U844 ( .A1(B[20]), .A2(n810), .ZN(N61) );
  AND2_X1 U845 ( .A1(B[19]), .A2(n810), .ZN(N60) );
  AND2_X1 U846 ( .A1(B[18]), .A2(n810), .ZN(N59) );
  AND2_X1 U847 ( .A1(B[17]), .A2(n810), .ZN(N58) );
  AND2_X1 U848 ( .A1(B[16]), .A2(n809), .ZN(N57) );
  AND2_X1 U849 ( .A1(B[15]), .A2(n809), .ZN(N56) );
  AND2_X1 U850 ( .A1(B[14]), .A2(n803), .ZN(N55) );
  AND2_X1 U851 ( .A1(B[13]), .A2(n809), .ZN(N54) );
  AND2_X1 U852 ( .A1(B[12]), .A2(n809), .ZN(N53) );
  AND2_X1 U853 ( .A1(B[11]), .A2(n809), .ZN(N52) );
  AND2_X1 U854 ( .A1(B[10]), .A2(n808), .ZN(N51) );
  AND2_X1 U855 ( .A1(B[9]), .A2(n808), .ZN(N50) );
  AND2_X1 U856 ( .A1(B[8]), .A2(n808), .ZN(N49) );
  AND2_X1 U857 ( .A1(B[7]), .A2(n808), .ZN(N48) );
  AND2_X1 U858 ( .A1(B[6]), .A2(n808), .ZN(N47) );
  AND2_X1 U859 ( .A1(B[5]), .A2(n807), .ZN(N46) );
  AND2_X1 U860 ( .A1(B[4]), .A2(n807), .ZN(N45) );
  AND2_X1 U861 ( .A1(B[3]), .A2(n807), .ZN(N44) );
  AND2_X1 U862 ( .A1(B[2]), .A2(n807), .ZN(N43) );
  AND2_X1 U863 ( .A1(B[1]), .A2(n807), .ZN(N42) );
  MUX2_X1 U864 ( .A(N334), .B(n638), .S(n788), .Z(n598) );
  NAND4_X1 U865 ( .A1(n405), .A2(n404), .A3(n403), .A4(n825), .ZN(n827) );
  NOR2_X1 U866 ( .A1(n439), .A2(n723), .ZN(N829) );
  MUX2_X1 U867 ( .A(n725), .B(n639), .S(n788), .Z(n597) );
  NOR2_X1 U868 ( .A1(n438), .A2(n721), .ZN(N831) );
  MUX2_X1 U869 ( .A(N332), .B(n640), .S(n787), .Z(n596) );
  NOR2_X1 U870 ( .A1(n437), .A2(n721), .ZN(N833) );
  MUX2_X1 U871 ( .A(N331), .B(n641), .S(n788), .Z(n595) );
  NOR2_X1 U872 ( .A1(n436), .A2(n743), .ZN(N835) );
  MUX2_X1 U873 ( .A(N330), .B(n642), .S(n788), .Z(n594) );
  NOR2_X1 U874 ( .A1(n435), .A2(n723), .ZN(N837) );
  MUX2_X1 U875 ( .A(N329), .B(n643), .S(n787), .Z(n593) );
  NOR2_X1 U876 ( .A1(n434), .A2(n721), .ZN(N839) );
  MUX2_X1 U877 ( .A(N328), .B(n644), .S(n786), .Z(n592) );
  NOR2_X1 U878 ( .A1(n433), .A2(n743), .ZN(N841) );
  MUX2_X1 U879 ( .A(N327), .B(n645), .S(n787), .Z(n591) );
  NOR2_X1 U880 ( .A1(n432), .A2(n743), .ZN(N843) );
  MUX2_X1 U881 ( .A(N326), .B(n646), .S(n787), .Z(n590) );
  NOR2_X1 U882 ( .A1(n431), .A2(n747), .ZN(N845) );
  MUX2_X1 U883 ( .A(N325), .B(n647), .S(n787), .Z(n589) );
  NOR2_X1 U884 ( .A1(n430), .A2(n721), .ZN(N847) );
  MUX2_X1 U885 ( .A(N324), .B(n648), .S(n787), .Z(n588) );
  NOR2_X1 U886 ( .A1(n429), .A2(n723), .ZN(N849) );
  MUX2_X1 U887 ( .A(N323), .B(n649), .S(n787), .Z(n587) );
  NOR2_X1 U888 ( .A1(n428), .A2(n723), .ZN(N851) );
  MUX2_X1 U889 ( .A(N322), .B(n650), .S(n787), .Z(n586) );
  NOR2_X1 U890 ( .A1(n427), .A2(n743), .ZN(N853) );
  MUX2_X1 U891 ( .A(N321), .B(n651), .S(n786), .Z(n585) );
  NOR2_X1 U892 ( .A1(n426), .A2(n721), .ZN(N855) );
  MUX2_X1 U893 ( .A(N320), .B(n652), .S(n787), .Z(n584) );
  NOR2_X1 U894 ( .A1(n425), .A2(n721), .ZN(N857) );
  MUX2_X1 U895 ( .A(N319), .B(n653), .S(n786), .Z(n583) );
  NOR2_X1 U896 ( .A1(n424), .A2(n747), .ZN(N859) );
  MUX2_X1 U897 ( .A(N318), .B(n654), .S(n787), .Z(n582) );
  NOR2_X1 U898 ( .A1(n423), .A2(n721), .ZN(N861) );
  MUX2_X1 U899 ( .A(N317), .B(n655), .S(n786), .Z(n581) );
  NOR2_X1 U900 ( .A1(n422), .A2(n747), .ZN(N863) );
  MUX2_X1 U901 ( .A(N316), .B(n656), .S(n787), .Z(n580) );
  NOR2_X1 U902 ( .A1(n421), .A2(n723), .ZN(N865) );
  MUX2_X1 U903 ( .A(N315), .B(n657), .S(n787), .Z(n579) );
  NOR2_X1 U904 ( .A1(n420), .A2(n723), .ZN(N867) );
  MUX2_X1 U905 ( .A(N314), .B(n658), .S(n786), .Z(n578) );
  NOR2_X1 U906 ( .A1(n419), .A2(n743), .ZN(N869) );
  MUX2_X1 U907 ( .A(N313), .B(n659), .S(n787), .Z(n577) );
  NOR2_X1 U908 ( .A1(n418), .A2(n723), .ZN(N871) );
  MUX2_X1 U909 ( .A(N312), .B(n660), .S(n787), .Z(n576) );
  NOR2_X1 U910 ( .A1(n417), .A2(n721), .ZN(N873) );
  MUX2_X1 U911 ( .A(N311), .B(n661), .S(n786), .Z(n575) );
  NOR2_X1 U912 ( .A1(n416), .A2(n743), .ZN(N875) );
  MUX2_X1 U913 ( .A(N310), .B(n662), .S(n787), .Z(n574) );
  NOR2_X1 U914 ( .A1(n415), .A2(n747), .ZN(N877) );
  MUX2_X1 U915 ( .A(N309), .B(n663), .S(n787), .Z(n573) );
  NOR2_X1 U916 ( .A1(n414), .A2(n723), .ZN(N879) );
  MUX2_X1 U917 ( .A(N308), .B(n664), .S(n786), .Z(n572) );
  NOR2_X1 U918 ( .A1(n413), .A2(n721), .ZN(N881) );
  MUX2_X1 U919 ( .A(N307), .B(n665), .S(n786), .Z(n571) );
  NOR2_X1 U920 ( .A1(n412), .A2(n723), .ZN(N883) );
  MUX2_X1 U921 ( .A(N306), .B(n666), .S(n787), .Z(n570) );
  NOR2_X1 U922 ( .A1(n411), .A2(n721), .ZN(N885) );
  MUX2_X1 U923 ( .A(N305), .B(n667), .S(n786), .Z(n569) );
  NOR2_X1 U924 ( .A1(n410), .A2(n743), .ZN(N887) );
  MUX2_X1 U925 ( .A(N304), .B(n668), .S(n786), .Z(n568) );
  NOR2_X1 U926 ( .A1(n409), .A2(n721), .ZN(N889) );
  MUX2_X1 U927 ( .A(N303), .B(n634), .S(n785), .Z(n599) );
  NAND2_X1 U928 ( .A1(n897), .A2(B_reg[31]), .ZN(n826) );
  INV_X1 U929 ( .A(n826), .ZN(n860) );
  AOI22_X1 U930 ( .A1(N172), .A2(n727), .B1(n827), .B2(n634), .ZN(n828) );
  INV_X1 U931 ( .A(n828), .ZN(n969) );
  MUX2_X1 U932 ( .A(n969), .B(n669), .S(n786), .Z(n535) );
  NAND2_X1 U933 ( .A1(n338), .A2(n897), .ZN(n829) );
  INV_X1 U934 ( .A(n829), .ZN(n861) );
  AOI22_X1 U935 ( .A1(B_reg[30]), .A2(n728), .B1(N171), .B2(n727), .ZN(n830)
         );
  OAI21_X1 U936 ( .B1(n339), .B2(n721), .A(n830), .ZN(n600) );
  MUX2_X1 U937 ( .A(n600), .B(n670), .S(n786), .Z(n534) );
  AOI22_X1 U938 ( .A1(B_reg[29]), .A2(n728), .B1(N170), .B2(n726), .ZN(n831)
         );
  OAI21_X1 U939 ( .B1(n337), .B2(n746), .A(n831), .ZN(n601) );
  MUX2_X1 U940 ( .A(n601), .B(n671), .S(n786), .Z(n533) );
  AOI22_X1 U941 ( .A1(B_reg[28]), .A2(n728), .B1(N169), .B2(n726), .ZN(n832)
         );
  OAI21_X1 U942 ( .B1(n336), .B2(n746), .A(n832), .ZN(n602) );
  MUX2_X1 U943 ( .A(n602), .B(n672), .S(n786), .Z(n532) );
  AOI22_X1 U944 ( .A1(B_reg[27]), .A2(n728), .B1(N168), .B2(n726), .ZN(n833)
         );
  OAI21_X1 U945 ( .B1(n335), .B2(n746), .A(n833), .ZN(n603) );
  MUX2_X1 U946 ( .A(n603), .B(n673), .S(n786), .Z(n531) );
  AOI22_X1 U947 ( .A1(B_reg[26]), .A2(n728), .B1(N167), .B2(n726), .ZN(n834)
         );
  OAI21_X1 U948 ( .B1(n334), .B2(n746), .A(n834), .ZN(n604) );
  MUX2_X1 U949 ( .A(n604), .B(n674), .S(n786), .Z(n530) );
  AOI22_X1 U950 ( .A1(B_reg[25]), .A2(n728), .B1(N166), .B2(n727), .ZN(n835)
         );
  OAI21_X1 U951 ( .B1(n333), .B2(n746), .A(n835), .ZN(n605) );
  MUX2_X1 U952 ( .A(n605), .B(n675), .S(n786), .Z(n529) );
  AOI22_X1 U953 ( .A1(B_reg[24]), .A2(n728), .B1(N165), .B2(n726), .ZN(n836)
         );
  OAI21_X1 U954 ( .B1(n332), .B2(n746), .A(n836), .ZN(n606) );
  MUX2_X1 U955 ( .A(n606), .B(n676), .S(n785), .Z(n528) );
  AOI22_X1 U956 ( .A1(B_reg[23]), .A2(n728), .B1(N164), .B2(n726), .ZN(n837)
         );
  OAI21_X1 U957 ( .B1(n331), .B2(n746), .A(n837), .ZN(n607) );
  MUX2_X1 U958 ( .A(n607), .B(n677), .S(n785), .Z(n527) );
  AOI22_X1 U959 ( .A1(B_reg[22]), .A2(n728), .B1(N163), .B2(n726), .ZN(n838)
         );
  OAI21_X1 U960 ( .B1(n330), .B2(n746), .A(n838), .ZN(n608) );
  MUX2_X1 U961 ( .A(n608), .B(n678), .S(n785), .Z(n526) );
  AOI22_X1 U962 ( .A1(B_reg[21]), .A2(n728), .B1(N162), .B2(n727), .ZN(n839)
         );
  OAI21_X1 U963 ( .B1(n329), .B2(n721), .A(n839), .ZN(n609) );
  MUX2_X1 U964 ( .A(n609), .B(n679), .S(n785), .Z(n525) );
  AOI22_X1 U965 ( .A1(B_reg[20]), .A2(n728), .B1(N161), .B2(n726), .ZN(n840)
         );
  OAI21_X1 U966 ( .B1(n328), .B2(n723), .A(n840), .ZN(n610) );
  MUX2_X1 U967 ( .A(n610), .B(n680), .S(n785), .Z(n524) );
  AOI22_X1 U968 ( .A1(B_reg[19]), .A2(n728), .B1(N160), .B2(n726), .ZN(n841)
         );
  OAI21_X1 U969 ( .B1(n327), .B2(n743), .A(n841), .ZN(n611) );
  MUX2_X1 U970 ( .A(n611), .B(n681), .S(n785), .Z(n523) );
  AOI22_X1 U971 ( .A1(B_reg[18]), .A2(n728), .B1(N159), .B2(n727), .ZN(n842)
         );
  OAI21_X1 U972 ( .B1(n326), .B2(n723), .A(n842), .ZN(n612) );
  MUX2_X1 U973 ( .A(n612), .B(n682), .S(n785), .Z(n522) );
  AOI22_X1 U974 ( .A1(B_reg[17]), .A2(n728), .B1(N158), .B2(n726), .ZN(n843)
         );
  OAI21_X1 U975 ( .B1(n325), .B2(n723), .A(n843), .ZN(n613) );
  MUX2_X1 U976 ( .A(n613), .B(n683), .S(n785), .Z(n521) );
  AOI22_X1 U977 ( .A1(B_reg[16]), .A2(n730), .B1(N157), .B2(n726), .ZN(n844)
         );
  OAI21_X1 U978 ( .B1(n324), .B2(n721), .A(n844), .ZN(n614) );
  MUX2_X1 U979 ( .A(n614), .B(n684), .S(n785), .Z(n520) );
  AOI22_X1 U980 ( .A1(B_reg[15]), .A2(n729), .B1(N156), .B2(n726), .ZN(n845)
         );
  OAI21_X1 U981 ( .B1(n323), .B2(n721), .A(n845), .ZN(n615) );
  MUX2_X1 U982 ( .A(n615), .B(n685), .S(n785), .Z(n519) );
  AOI22_X1 U983 ( .A1(B_reg[14]), .A2(n730), .B1(N155), .B2(n727), .ZN(n846)
         );
  OAI21_X1 U984 ( .B1(n322), .B2(n747), .A(n846), .ZN(n616) );
  MUX2_X1 U985 ( .A(n616), .B(n686), .S(n785), .Z(n518) );
  AOI22_X1 U986 ( .A1(B_reg[13]), .A2(n729), .B1(N154), .B2(n726), .ZN(n847)
         );
  OAI21_X1 U987 ( .B1(n321), .B2(n721), .A(n847), .ZN(n617) );
  MUX2_X1 U988 ( .A(n617), .B(n687), .S(n785), .Z(n517) );
  AOI22_X1 U989 ( .A1(B_reg[12]), .A2(n861), .B1(N153), .B2(n860), .ZN(n848)
         );
  OAI21_X1 U990 ( .B1(n320), .B2(n743), .A(n848), .ZN(n618) );
  MUX2_X1 U991 ( .A(n618), .B(n688), .S(n785), .Z(n516) );
  AOI22_X1 U992 ( .A1(B_reg[11]), .A2(n861), .B1(N152), .B2(n860), .ZN(n849)
         );
  OAI21_X1 U993 ( .B1(n319), .B2(n723), .A(n849), .ZN(n619) );
  MUX2_X1 U994 ( .A(n619), .B(n689), .S(n785), .Z(n515) );
  AOI22_X1 U995 ( .A1(B_reg[10]), .A2(n861), .B1(N151), .B2(n860), .ZN(n850)
         );
  OAI21_X1 U996 ( .B1(n318), .B2(n723), .A(n850), .ZN(n620) );
  MUX2_X1 U997 ( .A(n620), .B(n690), .S(n785), .Z(n514) );
  AOI22_X1 U998 ( .A1(B_reg[9]), .A2(n861), .B1(N150), .B2(n860), .ZN(n851) );
  OAI21_X1 U999 ( .B1(n317), .B2(n721), .A(n851), .ZN(n621) );
  MUX2_X1 U1000 ( .A(n621), .B(n691), .S(n785), .Z(n513) );
  AOI22_X1 U1001 ( .A1(B_reg[8]), .A2(n861), .B1(N149), .B2(n860), .ZN(n852)
         );
  OAI21_X1 U1002 ( .B1(n316), .B2(n743), .A(n852), .ZN(n622) );
  MUX2_X1 U1003 ( .A(n622), .B(n692), .S(n784), .Z(n512) );
  AOI22_X1 U1004 ( .A1(B_reg[7]), .A2(n861), .B1(N148), .B2(n860), .ZN(n853)
         );
  OAI21_X1 U1005 ( .B1(n315), .B2(n721), .A(n853), .ZN(n623) );
  MUX2_X1 U1006 ( .A(n623), .B(n693), .S(n784), .Z(n511) );
  AOI22_X1 U1007 ( .A1(B_reg[6]), .A2(n861), .B1(N147), .B2(n860), .ZN(n854)
         );
  OAI21_X1 U1008 ( .B1(n314), .B2(n743), .A(n854), .ZN(n624) );
  MUX2_X1 U1009 ( .A(n624), .B(n694), .S(n784), .Z(n510) );
  AOI22_X1 U1010 ( .A1(B_reg[5]), .A2(n861), .B1(N146), .B2(n860), .ZN(n855)
         );
  OAI21_X1 U1011 ( .B1(n313), .B2(n721), .A(n855), .ZN(n625) );
  MUX2_X1 U1012 ( .A(n625), .B(n695), .S(n784), .Z(n509) );
  AOI22_X1 U1013 ( .A1(B_reg[4]), .A2(n861), .B1(N145), .B2(n860), .ZN(n856)
         );
  OAI21_X1 U1014 ( .B1(n312), .B2(n723), .A(n856), .ZN(n626) );
  MUX2_X1 U1015 ( .A(n626), .B(n696), .S(n784), .Z(n508) );
  AOI22_X1 U1016 ( .A1(B_reg[3]), .A2(n861), .B1(N144), .B2(n860), .ZN(n857)
         );
  OAI21_X1 U1017 ( .B1(n311), .B2(n721), .A(n857), .ZN(n627) );
  MUX2_X1 U1018 ( .A(n627), .B(n697), .S(n784), .Z(n507) );
  AOI22_X1 U1019 ( .A1(B_reg[2]), .A2(n861), .B1(N143), .B2(n860), .ZN(n858)
         );
  OAI21_X1 U1020 ( .B1(n310), .B2(n743), .A(n858), .ZN(n628) );
  MUX2_X1 U1021 ( .A(n628), .B(n698), .S(n784), .Z(n506) );
  AOI22_X1 U1022 ( .A1(B_reg[1]), .A2(n861), .B1(N142), .B2(n860), .ZN(n859)
         );
  OAI21_X1 U1023 ( .B1(n309), .B2(n721), .A(n859), .ZN(n629) );
  MUX2_X1 U1024 ( .A(n629), .B(n699), .S(n784), .Z(n472) );
  AOI22_X1 U1025 ( .A1(B_reg[0]), .A2(n718), .B1(N141), .B2(n724), .ZN(n862)
         );
  INV_X1 U1026 ( .A(A[31]), .ZN(n863) );
  NOR2_X1 U1027 ( .A1(n788), .A2(n863), .ZN(N40) );
  AND2_X1 U1028 ( .A1(A[0]), .A2(n806), .ZN(N9) );
  NAND2_X1 U1029 ( .A1(n736), .A2(A_reg[31]), .ZN(n896) );
  NAND2_X1 U1030 ( .A1(n407), .A2(n736), .ZN(n893) );
  OAI222_X1 U1031 ( .A1(n741), .A2(n406), .B1(n406), .B2(n731), .C1(n408), 
        .C2(n736), .ZN(n567) );
  OAI222_X1 U1032 ( .A1(n899), .A2(n406), .B1(n406), .B2(n716), .C1(n408), 
        .C2(n746), .ZN(N236) );
  AND2_X1 U1033 ( .A1(A[1]), .A2(n806), .ZN(N10) );
  AND2_X1 U1034 ( .A1(A[30]), .A2(n806), .ZN(N39) );
  AND2_X1 U1035 ( .A1(A[29]), .A2(n806), .ZN(N38) );
  AND2_X1 U1036 ( .A1(A[28]), .A2(n806), .ZN(N37) );
  AND2_X1 U1037 ( .A1(A[27]), .A2(n805), .ZN(N36) );
  AND2_X1 U1038 ( .A1(A[26]), .A2(n805), .ZN(N35) );
  AND2_X1 U1039 ( .A1(A[25]), .A2(n805), .ZN(N34) );
  AND2_X1 U1040 ( .A1(A[24]), .A2(n805), .ZN(N33) );
  AND2_X1 U1041 ( .A1(A[23]), .A2(n805), .ZN(N32) );
  AND2_X1 U1042 ( .A1(A[22]), .A2(n804), .ZN(N31) );
  AND2_X1 U1043 ( .A1(A[21]), .A2(n804), .ZN(N30) );
  AND2_X1 U1044 ( .A1(A[20]), .A2(n804), .ZN(N29) );
  AND2_X1 U1045 ( .A1(A[19]), .A2(n804), .ZN(N28) );
  AND2_X1 U1046 ( .A1(A[18]), .A2(n804), .ZN(N27) );
  AND2_X1 U1047 ( .A1(A[17]), .A2(n803), .ZN(N26) );
  AND2_X1 U1048 ( .A1(A[16]), .A2(n803), .ZN(N25) );
  AND2_X1 U1049 ( .A1(A[15]), .A2(n803), .ZN(N24) );
  AND2_X1 U1050 ( .A1(A[14]), .A2(n803), .ZN(N23) );
  AND2_X1 U1051 ( .A1(A[13]), .A2(n802), .ZN(N22) );
  AND2_X1 U1052 ( .A1(A[12]), .A2(n802), .ZN(N21) );
  AND2_X1 U1053 ( .A1(A[11]), .A2(n802), .ZN(N20) );
  AND2_X1 U1054 ( .A1(A[10]), .A2(n802), .ZN(N19) );
  AND2_X1 U1055 ( .A1(A[9]), .A2(n802), .ZN(N18) );
  AND2_X1 U1056 ( .A1(A[8]), .A2(n801), .ZN(N17) );
  AND2_X1 U1057 ( .A1(A[7]), .A2(n801), .ZN(N16) );
  AND2_X1 U1058 ( .A1(A[6]), .A2(n801), .ZN(N15) );
  AND2_X1 U1059 ( .A1(A[5]), .A2(n801), .ZN(N14) );
  AND2_X1 U1060 ( .A1(A[4]), .A2(n801), .ZN(N13) );
  AND2_X1 U1061 ( .A1(A[3]), .A2(n800), .ZN(N12) );
  AND2_X1 U1062 ( .A1(A[2]), .A2(n800), .ZN(N11) );
  INV_X1 U1063 ( .A(N77), .ZN(n864) );
  OAI222_X1 U1064 ( .A1(n741), .A2(n864), .B1(n399), .B2(n731), .C1(n400), 
        .C2(n738), .ZN(n566) );
  OAI222_X1 U1065 ( .A1(n706), .A2(n864), .B1(n399), .B2(n719), .C1(n400), 
        .C2(n746), .ZN(N235) );
  INV_X1 U1066 ( .A(N78), .ZN(n865) );
  OAI222_X1 U1067 ( .A1(n741), .A2(n865), .B1(n397), .B2(n731), .C1(n398), 
        .C2(n738), .ZN(n565) );
  OAI222_X1 U1068 ( .A1(n707), .A2(n865), .B1(n397), .B2(n894), .C1(n398), 
        .C2(n746), .ZN(N234) );
  INV_X1 U1069 ( .A(N79), .ZN(n866) );
  OAI222_X1 U1070 ( .A1(n741), .A2(n866), .B1(n395), .B2(n731), .C1(n396), 
        .C2(n738), .ZN(n564) );
  OAI222_X1 U1071 ( .A1(n899), .A2(n866), .B1(n395), .B2(n719), .C1(n396), 
        .C2(n746), .ZN(N233) );
  INV_X1 U1072 ( .A(N80), .ZN(n867) );
  OAI222_X1 U1073 ( .A1(n741), .A2(n867), .B1(n393), .B2(n731), .C1(n394), 
        .C2(n738), .ZN(n563) );
  OAI222_X1 U1074 ( .A1(n899), .A2(n867), .B1(n393), .B2(n894), .C1(n394), 
        .C2(n748), .ZN(N232) );
  INV_X1 U1075 ( .A(N81), .ZN(n868) );
  OAI222_X1 U1076 ( .A1(n741), .A2(n868), .B1(n391), .B2(n731), .C1(n392), 
        .C2(n738), .ZN(n562) );
  OAI222_X1 U1077 ( .A1(n717), .A2(n868), .B1(n391), .B2(n719), .C1(n392), 
        .C2(n744), .ZN(N231) );
  INV_X1 U1078 ( .A(N82), .ZN(n869) );
  OAI222_X1 U1079 ( .A1(n741), .A2(n869), .B1(n389), .B2(n731), .C1(n390), 
        .C2(n738), .ZN(n561) );
  OAI222_X1 U1080 ( .A1(n706), .A2(n869), .B1(n389), .B2(n894), .C1(n390), 
        .C2(n746), .ZN(N230) );
  INV_X1 U1081 ( .A(N83), .ZN(n870) );
  OAI222_X1 U1082 ( .A1(n741), .A2(n870), .B1(n387), .B2(n731), .C1(n388), 
        .C2(n738), .ZN(n560) );
  OAI222_X1 U1083 ( .A1(n706), .A2(n870), .B1(n387), .B2(n894), .C1(n388), 
        .C2(n747), .ZN(N229) );
  INV_X1 U1084 ( .A(N84), .ZN(n871) );
  OAI222_X1 U1085 ( .A1(n740), .A2(n871), .B1(n385), .B2(n731), .C1(n386), 
        .C2(n738), .ZN(n559) );
  OAI222_X1 U1086 ( .A1(n899), .A2(n871), .B1(n385), .B2(n716), .C1(n386), 
        .C2(n747), .ZN(N228) );
  INV_X1 U1087 ( .A(N85), .ZN(n872) );
  OAI222_X1 U1088 ( .A1(n740), .A2(n872), .B1(n383), .B2(n731), .C1(n384), 
        .C2(n738), .ZN(n558) );
  OAI222_X1 U1089 ( .A1(n706), .A2(n872), .B1(n383), .B2(n716), .C1(n384), 
        .C2(n744), .ZN(N227) );
  INV_X1 U1090 ( .A(N86), .ZN(n873) );
  OAI222_X1 U1091 ( .A1(n740), .A2(n873), .B1(n381), .B2(n731), .C1(n382), 
        .C2(n738), .ZN(n557) );
  OAI222_X1 U1092 ( .A1(n707), .A2(n873), .B1(n381), .B2(n735), .C1(n382), 
        .C2(n748), .ZN(N226) );
  INV_X1 U1093 ( .A(N87), .ZN(n874) );
  OAI222_X1 U1094 ( .A1(n740), .A2(n874), .B1(n379), .B2(n731), .C1(n380), 
        .C2(n737), .ZN(n556) );
  OAI222_X1 U1095 ( .A1(n707), .A2(n874), .B1(n379), .B2(n735), .C1(n380), 
        .C2(n721), .ZN(N225) );
  INV_X1 U1096 ( .A(N88), .ZN(n875) );
  OAI222_X1 U1097 ( .A1(n740), .A2(n875), .B1(n377), .B2(n732), .C1(n378), 
        .C2(n737), .ZN(n555) );
  OAI222_X1 U1098 ( .A1(n720), .A2(n875), .B1(n377), .B2(n894), .C1(n378), 
        .C2(n721), .ZN(N224) );
  INV_X1 U1099 ( .A(N89), .ZN(n876) );
  OAI222_X1 U1100 ( .A1(n740), .A2(n876), .B1(n375), .B2(n732), .C1(n376), 
        .C2(n737), .ZN(n554) );
  OAI222_X1 U1101 ( .A1(n720), .A2(n876), .B1(n375), .B2(n719), .C1(n376), 
        .C2(n721), .ZN(N223) );
  INV_X1 U1102 ( .A(N90), .ZN(n877) );
  OAI222_X1 U1103 ( .A1(n740), .A2(n877), .B1(n373), .B2(n732), .C1(n374), 
        .C2(n737), .ZN(n553) );
  OAI222_X1 U1104 ( .A1(n720), .A2(n877), .B1(n373), .B2(n734), .C1(n374), 
        .C2(n721), .ZN(N222) );
  INV_X1 U1105 ( .A(N91), .ZN(n878) );
  OAI222_X1 U1106 ( .A1(n740), .A2(n878), .B1(n371), .B2(n732), .C1(n372), 
        .C2(n737), .ZN(n552) );
  OAI222_X1 U1107 ( .A1(n720), .A2(n878), .B1(n371), .B2(n734), .C1(n372), 
        .C2(n721), .ZN(N221) );
  INV_X1 U1108 ( .A(N92), .ZN(n879) );
  OAI222_X1 U1109 ( .A1(n740), .A2(n879), .B1(n369), .B2(n732), .C1(n370), 
        .C2(n737), .ZN(n551) );
  OAI222_X1 U1110 ( .A1(n720), .A2(n879), .B1(n369), .B2(n734), .C1(n370), 
        .C2(n721), .ZN(N220) );
  INV_X1 U1111 ( .A(N93), .ZN(n880) );
  OAI222_X1 U1112 ( .A1(n740), .A2(n880), .B1(n367), .B2(n732), .C1(n368), 
        .C2(n737), .ZN(n550) );
  OAI222_X1 U1113 ( .A1(n720), .A2(n880), .B1(n367), .B2(n734), .C1(n368), 
        .C2(n747), .ZN(N219) );
  INV_X1 U1114 ( .A(N94), .ZN(n881) );
  OAI222_X1 U1115 ( .A1(n740), .A2(n881), .B1(n365), .B2(n732), .C1(n366), 
        .C2(n737), .ZN(n549) );
  OAI222_X1 U1116 ( .A1(n720), .A2(n881), .B1(n365), .B2(n734), .C1(n366), 
        .C2(n747), .ZN(N218) );
  INV_X1 U1117 ( .A(N95), .ZN(n882) );
  OAI222_X1 U1118 ( .A1(n740), .A2(n882), .B1(n363), .B2(n732), .C1(n364), 
        .C2(n737), .ZN(n548) );
  OAI222_X1 U1119 ( .A1(n720), .A2(n882), .B1(n363), .B2(n734), .C1(n364), 
        .C2(n747), .ZN(N217) );
  INV_X1 U1120 ( .A(N96), .ZN(n883) );
  OAI222_X1 U1121 ( .A1(n739), .A2(n883), .B1(n361), .B2(n732), .C1(n362), 
        .C2(n737), .ZN(n547) );
  OAI222_X1 U1122 ( .A1(n720), .A2(n883), .B1(n361), .B2(n734), .C1(n362), 
        .C2(n747), .ZN(N216) );
  INV_X1 U1123 ( .A(N97), .ZN(n884) );
  OAI222_X1 U1124 ( .A1(n739), .A2(n884), .B1(n359), .B2(n732), .C1(n360), 
        .C2(n737), .ZN(n546) );
  OAI222_X1 U1125 ( .A1(n720), .A2(n884), .B1(n359), .B2(n734), .C1(n360), 
        .C2(n747), .ZN(N215) );
  INV_X1 U1126 ( .A(N98), .ZN(n885) );
  OAI222_X1 U1127 ( .A1(n739), .A2(n885), .B1(n357), .B2(n732), .C1(n358), 
        .C2(n736), .ZN(n545) );
  OAI222_X1 U1128 ( .A1(n720), .A2(n885), .B1(n357), .B2(n734), .C1(n358), 
        .C2(n747), .ZN(N214) );
  INV_X1 U1129 ( .A(N99), .ZN(n886) );
  OAI222_X1 U1130 ( .A1(n739), .A2(n886), .B1(n355), .B2(n732), .C1(n356), 
        .C2(n737), .ZN(n544) );
  OAI222_X1 U1131 ( .A1(n720), .A2(n886), .B1(n355), .B2(n734), .C1(n356), 
        .C2(n747), .ZN(N213) );
  INV_X1 U1132 ( .A(N100), .ZN(n887) );
  OAI222_X1 U1133 ( .A1(n739), .A2(n887), .B1(n353), .B2(n733), .C1(n354), 
        .C2(n736), .ZN(n543) );
  OAI222_X1 U1134 ( .A1(n720), .A2(n887), .B1(n353), .B2(n734), .C1(n354), 
        .C2(n747), .ZN(N212) );
  INV_X1 U1135 ( .A(N101), .ZN(n888) );
  OAI222_X1 U1136 ( .A1(n739), .A2(n888), .B1(n351), .B2(n733), .C1(n352), 
        .C2(n736), .ZN(n542) );
  OAI222_X1 U1137 ( .A1(n720), .A2(n888), .B1(n351), .B2(n734), .C1(n352), 
        .C2(n747), .ZN(N211) );
  INV_X1 U1138 ( .A(N102), .ZN(n889) );
  OAI222_X1 U1139 ( .A1(n739), .A2(n889), .B1(n349), .B2(n733), .C1(n350), 
        .C2(n736), .ZN(n541) );
  OAI222_X1 U1140 ( .A1(n720), .A2(n889), .B1(n349), .B2(n734), .C1(n350), 
        .C2(n747), .ZN(N210) );
  INV_X1 U1141 ( .A(N103), .ZN(n890) );
  OAI222_X1 U1142 ( .A1(n739), .A2(n890), .B1(n347), .B2(n733), .C1(n348), 
        .C2(n736), .ZN(n540) );
  OAI222_X1 U1143 ( .A1(n720), .A2(n890), .B1(n347), .B2(n734), .C1(n348), 
        .C2(n747), .ZN(N209) );
  INV_X1 U1144 ( .A(N104), .ZN(n891) );
  OAI222_X1 U1145 ( .A1(n739), .A2(n891), .B1(n345), .B2(n733), .C1(n346), 
        .C2(n736), .ZN(n539) );
  OAI222_X1 U1146 ( .A1(n720), .A2(n891), .B1(n345), .B2(n734), .C1(n346), 
        .C2(n747), .ZN(N208) );
  INV_X1 U1147 ( .A(N105), .ZN(n892) );
  OAI222_X1 U1148 ( .A1(n739), .A2(n892), .B1(n343), .B2(n733), .C1(n344), 
        .C2(n736), .ZN(n538) );
  OAI222_X1 U1149 ( .A1(n720), .A2(n892), .B1(n343), .B2(n734), .C1(n344), 
        .C2(n748), .ZN(N207) );
  INV_X1 U1150 ( .A(N106), .ZN(n895) );
  OAI222_X1 U1151 ( .A1(n739), .A2(n895), .B1(n341), .B2(n733), .C1(n342), 
        .C2(n736), .ZN(n537) );
  OAI222_X1 U1152 ( .A1(n720), .A2(n895), .B1(n341), .B2(n734), .C1(n342), 
        .C2(n748), .ZN(N206) );
  INV_X1 U1153 ( .A(N107), .ZN(n898) );
  OAI22_X1 U1154 ( .A1(n898), .A2(n739), .B1(n340), .B2(n736), .ZN(n536) );
  OAI22_X1 U1155 ( .A1(n720), .A2(n898), .B1(n340), .B2(n743), .ZN(N205) );
  NAND2_X1 U1156 ( .A1(n709), .A2(n800), .ZN(n967) );
  INV_X1 U1157 ( .A(n967), .ZN(n966) );
  XOR2_X1 U1158 ( .A(n900), .B(A[31]), .Z(n902) );
  INV_X1 U1159 ( .A(n902), .ZN(n901) );
  AOI22_X1 U1160 ( .A1(N337), .A2(n768), .B1(n757), .B2(n629), .ZN(n903) );
  OAI21_X1 U1161 ( .B1(n274), .B2(n760), .A(n903), .ZN(n471) );
  AOI22_X1 U1162 ( .A1(N338), .A2(n768), .B1(n757), .B2(n628), .ZN(n904) );
  OAI21_X1 U1163 ( .B1(n273), .B2(n760), .A(n904), .ZN(n470) );
  AOI22_X1 U1164 ( .A1(N339), .A2(n768), .B1(n757), .B2(n627), .ZN(n905) );
  OAI21_X1 U1165 ( .B1(n272), .B2(n760), .A(n905), .ZN(n469) );
  AOI22_X1 U1166 ( .A1(N340), .A2(n768), .B1(n756), .B2(n626), .ZN(n906) );
  OAI21_X1 U1167 ( .B1(n271), .B2(n760), .A(n906), .ZN(n468) );
  AOI22_X1 U1168 ( .A1(N341), .A2(n768), .B1(n756), .B2(n625), .ZN(n907) );
  OAI21_X1 U1169 ( .B1(n270), .B2(n760), .A(n907), .ZN(n467) );
  AOI22_X1 U1170 ( .A1(N342), .A2(n768), .B1(n756), .B2(n624), .ZN(n908) );
  OAI21_X1 U1171 ( .B1(n269), .B2(n760), .A(n908), .ZN(n466) );
  AOI22_X1 U1172 ( .A1(N343), .A2(n768), .B1(n756), .B2(n623), .ZN(n909) );
  OAI21_X1 U1173 ( .B1(n268), .B2(n760), .A(n909), .ZN(n465) );
  AOI22_X1 U1174 ( .A1(N344), .A2(n768), .B1(n756), .B2(n622), .ZN(n910) );
  OAI21_X1 U1175 ( .B1(n267), .B2(n760), .A(n910), .ZN(n464) );
  AOI22_X1 U1176 ( .A1(N345), .A2(n768), .B1(n756), .B2(n621), .ZN(n911) );
  OAI21_X1 U1177 ( .B1(n266), .B2(n760), .A(n911), .ZN(n463) );
  AOI22_X1 U1178 ( .A1(N346), .A2(n768), .B1(n756), .B2(n620), .ZN(n912) );
  OAI21_X1 U1179 ( .B1(n265), .B2(n760), .A(n912), .ZN(n462) );
  AOI22_X1 U1180 ( .A1(N347), .A2(n768), .B1(n756), .B2(n619), .ZN(n913) );
  OAI21_X1 U1181 ( .B1(n264), .B2(n761), .A(n913), .ZN(n461) );
  AOI22_X1 U1182 ( .A1(N348), .A2(n768), .B1(n756), .B2(n618), .ZN(n914) );
  OAI21_X1 U1183 ( .B1(n263), .B2(n761), .A(n914), .ZN(n460) );
  AOI22_X1 U1184 ( .A1(N349), .A2(n769), .B1(n756), .B2(n617), .ZN(n915) );
  OAI21_X1 U1185 ( .B1(n262), .B2(n761), .A(n915), .ZN(n459) );
  AOI22_X1 U1186 ( .A1(N350), .A2(n769), .B1(n756), .B2(n616), .ZN(n916) );
  OAI21_X1 U1187 ( .B1(n261), .B2(n761), .A(n916), .ZN(n458) );
  AOI22_X1 U1188 ( .A1(N351), .A2(n769), .B1(n756), .B2(n615), .ZN(n917) );
  OAI21_X1 U1189 ( .B1(n260), .B2(n761), .A(n917), .ZN(n457) );
  AOI22_X1 U1190 ( .A1(N352), .A2(n769), .B1(n755), .B2(n614), .ZN(n918) );
  OAI21_X1 U1191 ( .B1(n259), .B2(n761), .A(n918), .ZN(n456) );
  AOI22_X1 U1192 ( .A1(N353), .A2(n769), .B1(n755), .B2(n613), .ZN(n919) );
  OAI21_X1 U1193 ( .B1(n258), .B2(n761), .A(n919), .ZN(n455) );
  AOI22_X1 U1194 ( .A1(N354), .A2(n769), .B1(n755), .B2(n612), .ZN(n920) );
  OAI21_X1 U1195 ( .B1(n257), .B2(n761), .A(n920), .ZN(n454) );
  AOI22_X1 U1196 ( .A1(N355), .A2(n769), .B1(n755), .B2(n611), .ZN(n921) );
  OAI21_X1 U1197 ( .B1(n256), .B2(n761), .A(n921), .ZN(n453) );
  AOI22_X1 U1198 ( .A1(N356), .A2(n769), .B1(n755), .B2(n610), .ZN(n922) );
  OAI21_X1 U1199 ( .B1(n255), .B2(n761), .A(n922), .ZN(n452) );
  AOI22_X1 U1200 ( .A1(N357), .A2(n769), .B1(n755), .B2(n609), .ZN(n923) );
  OAI21_X1 U1201 ( .B1(n254), .B2(n761), .A(n923), .ZN(n451) );
  AOI22_X1 U1202 ( .A1(N358), .A2(n769), .B1(n755), .B2(n608), .ZN(n924) );
  OAI21_X1 U1203 ( .B1(n253), .B2(n761), .A(n924), .ZN(n450) );
  AOI22_X1 U1204 ( .A1(N359), .A2(n769), .B1(n755), .B2(n607), .ZN(n925) );
  OAI21_X1 U1205 ( .B1(n252), .B2(n762), .A(n925), .ZN(n449) );
  AOI22_X1 U1206 ( .A1(N360), .A2(n769), .B1(n755), .B2(n606), .ZN(n926) );
  OAI21_X1 U1207 ( .B1(n251), .B2(n762), .A(n926), .ZN(n448) );
  AOI22_X1 U1208 ( .A1(N361), .A2(n770), .B1(n755), .B2(n605), .ZN(n927) );
  OAI21_X1 U1209 ( .B1(n250), .B2(n762), .A(n927), .ZN(n447) );
  AOI22_X1 U1210 ( .A1(N362), .A2(n770), .B1(n755), .B2(n604), .ZN(n928) );
  OAI21_X1 U1211 ( .B1(n249), .B2(n762), .A(n928), .ZN(n446) );
  AOI22_X1 U1212 ( .A1(N363), .A2(n770), .B1(n755), .B2(n603), .ZN(n929) );
  OAI21_X1 U1213 ( .B1(n248), .B2(n762), .A(n929), .ZN(n445) );
  AOI22_X1 U1214 ( .A1(N364), .A2(n770), .B1(n754), .B2(n602), .ZN(n930) );
  OAI21_X1 U1215 ( .B1(n247), .B2(n762), .A(n930), .ZN(n444) );
  AOI22_X1 U1216 ( .A1(N365), .A2(n770), .B1(n754), .B2(n601), .ZN(n931) );
  OAI21_X1 U1217 ( .B1(n246), .B2(n762), .A(n931), .ZN(n443) );
  AOI22_X1 U1218 ( .A1(N366), .A2(n770), .B1(n754), .B2(n600), .ZN(n932) );
  OAI21_X1 U1219 ( .B1(n245), .B2(n762), .A(n932), .ZN(n442) );
  AOI22_X1 U1220 ( .A1(N367), .A2(n770), .B1(n754), .B2(n969), .ZN(n933) );
  OAI21_X1 U1221 ( .B1(n244), .B2(n762), .A(n933), .ZN(n441) );
  NOR2_X1 U1222 ( .A1(n244), .A2(n789), .ZN(N563) );
  AOI22_X1 U1223 ( .A1(N368), .A2(n770), .B1(N303), .B2(n754), .ZN(n934) );
  OAI21_X1 U1224 ( .B1(n308), .B2(n762), .A(n934), .ZN(n505) );
  NOR2_X1 U1225 ( .A1(n308), .A2(n788), .ZN(N564) );
  AOI22_X1 U1226 ( .A1(N369), .A2(n770), .B1(N304), .B2(n754), .ZN(n935) );
  OAI21_X1 U1227 ( .B1(n307), .B2(n762), .A(n935), .ZN(n504) );
  NOR2_X1 U1228 ( .A1(n307), .A2(n788), .ZN(N565) );
  AOI22_X1 U1229 ( .A1(N370), .A2(n770), .B1(N305), .B2(n754), .ZN(n936) );
  OAI21_X1 U1230 ( .B1(n306), .B2(n762), .A(n936), .ZN(n503) );
  NOR2_X1 U1231 ( .A1(n306), .A2(n789), .ZN(N566) );
  AOI22_X1 U1232 ( .A1(N371), .A2(n770), .B1(N306), .B2(n754), .ZN(n937) );
  OAI21_X1 U1233 ( .B1(n305), .B2(n763), .A(n937), .ZN(n502) );
  NOR2_X1 U1234 ( .A1(n305), .A2(n788), .ZN(N567) );
  AOI22_X1 U1235 ( .A1(N372), .A2(n770), .B1(N307), .B2(n754), .ZN(n938) );
  OAI21_X1 U1236 ( .B1(n304), .B2(n763), .A(n938), .ZN(n501) );
  NOR2_X1 U1237 ( .A1(n304), .A2(n788), .ZN(N568) );
  AOI22_X1 U1238 ( .A1(N373), .A2(n771), .B1(N308), .B2(n754), .ZN(n939) );
  OAI21_X1 U1239 ( .B1(n303), .B2(n763), .A(n939), .ZN(n500) );
  NOR2_X1 U1240 ( .A1(n303), .A2(n789), .ZN(N569) );
  AOI22_X1 U1241 ( .A1(N374), .A2(n771), .B1(N309), .B2(n754), .ZN(n940) );
  OAI21_X1 U1242 ( .B1(n302), .B2(n763), .A(n940), .ZN(n499) );
  NOR2_X1 U1243 ( .A1(n302), .A2(n789), .ZN(N570) );
  AOI22_X1 U1244 ( .A1(N375), .A2(n771), .B1(N310), .B2(n754), .ZN(n941) );
  OAI21_X1 U1245 ( .B1(n301), .B2(n763), .A(n941), .ZN(n498) );
  NOR2_X1 U1246 ( .A1(n301), .A2(n788), .ZN(N571) );
  AOI22_X1 U1247 ( .A1(N376), .A2(n771), .B1(N311), .B2(n753), .ZN(n942) );
  OAI21_X1 U1248 ( .B1(n300), .B2(n763), .A(n942), .ZN(n497) );
  NOR2_X1 U1249 ( .A1(n300), .A2(n789), .ZN(N572) );
  AOI22_X1 U1250 ( .A1(N377), .A2(n771), .B1(N312), .B2(n753), .ZN(n943) );
  OAI21_X1 U1251 ( .B1(n299), .B2(n763), .A(n943), .ZN(n496) );
  NOR2_X1 U1252 ( .A1(n299), .A2(n788), .ZN(N573) );
  AOI22_X1 U1253 ( .A1(N378), .A2(n771), .B1(N313), .B2(n753), .ZN(n944) );
  OAI21_X1 U1254 ( .B1(n298), .B2(n763), .A(n944), .ZN(n495) );
  NOR2_X1 U1255 ( .A1(n298), .A2(n788), .ZN(N574) );
  AOI22_X1 U1256 ( .A1(N379), .A2(n771), .B1(N314), .B2(n753), .ZN(n945) );
  OAI21_X1 U1257 ( .B1(n297), .B2(n763), .A(n945), .ZN(n494) );
  NOR2_X1 U1258 ( .A1(n297), .A2(n789), .ZN(N575) );
  AOI22_X1 U1259 ( .A1(N380), .A2(n771), .B1(N315), .B2(n753), .ZN(n946) );
  OAI21_X1 U1260 ( .B1(n296), .B2(n763), .A(n946), .ZN(n493) );
  NOR2_X1 U1261 ( .A1(n296), .A2(n788), .ZN(N576) );
  AOI22_X1 U1262 ( .A1(N381), .A2(n771), .B1(N316), .B2(n753), .ZN(n947) );
  OAI21_X1 U1263 ( .B1(n295), .B2(n763), .A(n947), .ZN(n492) );
  NOR2_X1 U1264 ( .A1(n295), .A2(n790), .ZN(N577) );
  AOI22_X1 U1265 ( .A1(N382), .A2(n771), .B1(N317), .B2(n753), .ZN(n948) );
  OAI21_X1 U1266 ( .B1(n294), .B2(n763), .A(n948), .ZN(n491) );
  NOR2_X1 U1267 ( .A1(n294), .A2(n789), .ZN(N578) );
  AOI22_X1 U1268 ( .A1(N383), .A2(n771), .B1(N318), .B2(n753), .ZN(n949) );
  OAI21_X1 U1269 ( .B1(n293), .B2(n764), .A(n949), .ZN(n490) );
  NOR2_X1 U1270 ( .A1(n293), .A2(n788), .ZN(N579) );
  AOI22_X1 U1271 ( .A1(N384), .A2(n771), .B1(N319), .B2(n753), .ZN(n950) );
  OAI21_X1 U1272 ( .B1(n292), .B2(n764), .A(n950), .ZN(n489) );
  NOR2_X1 U1273 ( .A1(n292), .A2(n788), .ZN(N580) );
  AOI22_X1 U1274 ( .A1(N385), .A2(n772), .B1(N320), .B2(n753), .ZN(n951) );
  OAI21_X1 U1275 ( .B1(n291), .B2(n764), .A(n951), .ZN(n488) );
  NOR2_X1 U1276 ( .A1(n291), .A2(n789), .ZN(N581) );
  AOI22_X1 U1277 ( .A1(N386), .A2(n772), .B1(N321), .B2(n753), .ZN(n952) );
  OAI21_X1 U1278 ( .B1(n290), .B2(n764), .A(n952), .ZN(n487) );
  NOR2_X1 U1279 ( .A1(n290), .A2(n788), .ZN(N582) );
  AOI22_X1 U1280 ( .A1(N387), .A2(n772), .B1(N322), .B2(n753), .ZN(n953) );
  OAI21_X1 U1281 ( .B1(n289), .B2(n764), .A(n953), .ZN(n486) );
  NOR2_X1 U1282 ( .A1(n289), .A2(n788), .ZN(N583) );
  AOI22_X1 U1283 ( .A1(N388), .A2(n772), .B1(N323), .B2(n752), .ZN(n954) );
  OAI21_X1 U1284 ( .B1(n288), .B2(n764), .A(n954), .ZN(n485) );
  NOR2_X1 U1285 ( .A1(n288), .A2(n789), .ZN(N584) );
  AOI22_X1 U1286 ( .A1(N389), .A2(n772), .B1(N324), .B2(n752), .ZN(n955) );
  OAI21_X1 U1287 ( .B1(n287), .B2(n764), .A(n955), .ZN(n484) );
  NOR2_X1 U1288 ( .A1(n287), .A2(n789), .ZN(N585) );
  AOI22_X1 U1289 ( .A1(N390), .A2(n772), .B1(N325), .B2(n752), .ZN(n956) );
  OAI21_X1 U1290 ( .B1(n286), .B2(n764), .A(n956), .ZN(n483) );
  NOR2_X1 U1291 ( .A1(n286), .A2(n789), .ZN(N586) );
  AOI22_X1 U1292 ( .A1(N391), .A2(n772), .B1(N326), .B2(n752), .ZN(n957) );
  OAI21_X1 U1293 ( .B1(n285), .B2(n764), .A(n957), .ZN(n482) );
  NOR2_X1 U1294 ( .A1(n285), .A2(n789), .ZN(N587) );
  AOI22_X1 U1295 ( .A1(N392), .A2(n772), .B1(N327), .B2(n752), .ZN(n958) );
  OAI21_X1 U1296 ( .B1(n284), .B2(n764), .A(n958), .ZN(n481) );
  NOR2_X1 U1297 ( .A1(n284), .A2(n789), .ZN(N588) );
  AOI22_X1 U1298 ( .A1(N393), .A2(n772), .B1(N328), .B2(n752), .ZN(n959) );
  OAI21_X1 U1299 ( .B1(n283), .B2(n764), .A(n959), .ZN(n480) );
  NOR2_X1 U1300 ( .A1(n283), .A2(n789), .ZN(N589) );
  AOI22_X1 U1301 ( .A1(N394), .A2(n772), .B1(N329), .B2(n752), .ZN(n960) );
  OAI21_X1 U1302 ( .B1(n282), .B2(n764), .A(n960), .ZN(n479) );
  NOR2_X1 U1303 ( .A1(n282), .A2(n790), .ZN(N590) );
  AOI22_X1 U1304 ( .A1(N395), .A2(n772), .B1(N330), .B2(n752), .ZN(n961) );
  OAI21_X1 U1305 ( .B1(n281), .B2(n765), .A(n961), .ZN(n478) );
  NOR2_X1 U1306 ( .A1(n281), .A2(n789), .ZN(N591) );
  AOI22_X1 U1307 ( .A1(N396), .A2(n772), .B1(N331), .B2(n752), .ZN(n962) );
  OAI21_X1 U1308 ( .B1(n280), .B2(n765), .A(n962), .ZN(n477) );
  NOR2_X1 U1309 ( .A1(n280), .A2(n789), .ZN(N592) );
  AOI22_X1 U1310 ( .A1(N397), .A2(n773), .B1(N332), .B2(n752), .ZN(n963) );
  OAI21_X1 U1311 ( .B1(n279), .B2(n765), .A(n963), .ZN(n476) );
  NOR2_X1 U1312 ( .A1(n279), .A2(n789), .ZN(N593) );
  AOI22_X1 U1313 ( .A1(N398), .A2(n773), .B1(n725), .B2(n752), .ZN(n964) );
  OAI21_X1 U1314 ( .B1(n278), .B2(n765), .A(n964), .ZN(n475) );
  NOR2_X1 U1315 ( .A1(n278), .A2(n789), .ZN(N594) );
  AOI22_X1 U1316 ( .A1(N399), .A2(n773), .B1(N334), .B2(n752), .ZN(n965) );
  OAI21_X1 U1317 ( .B1(n277), .B2(n765), .A(n965), .ZN(n474) );
  NOR2_X1 U1318 ( .A1(n277), .A2(n789), .ZN(N595) );
  AOI22_X1 U1319 ( .A1(n967), .A2(n637), .B1(N400), .B2(n773), .ZN(n968) );
  INV_X1 U1320 ( .A(n968), .ZN(n473) );
  NOR2_X1 U1321 ( .A1(n276), .A2(n790), .ZN(N596) );
endmodule

